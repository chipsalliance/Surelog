module bot ();
endmodule

