/*
:name: resetall-directive
:description: Check for the resetall directive
:should_fail: 0
:tags: 5.6.4
*/

`resetall

module ts();
endmodule
