/*
:name: number_test_60
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = 'h 0;