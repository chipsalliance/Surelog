/*
:name: 22.5.3--undefineall-basic
:description: Test
:should_fail: 0
:tags: 22.5.3
:type: preprocessing
*/
`undefineall
