

package dv_utils_pkg;
 
  `include "dv_macros.vh"
 

endpackage


`define first_half "start of string
module top ();
$display(`first_half end of string");
endmodule
