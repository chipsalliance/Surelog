/*
:name: typedef_test_6
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef struct { int i; bit b; } mystruct;
