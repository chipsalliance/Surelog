
`include "prim_assert.sv"

module top (input logic b, output logic a);
 

`ASSERT(SigintEventCheck_A, sigint_o |-> !event_o)

   assign a = b;

   
`ASSERT(SigintEventCheck_A, 
    sigint_o |-> !event_o)

   assign a = b;


  `define _N(stg) (16 >> stg)

   assign a = b;

     `define _N(stg) (16 >> stg)
  
      // bext / bdep control bit generation   

 assign a = b;



 prim_subreg #(
     .DW      (1)
  ) u_ip0_p7 (
   .clk_i   (clk_i    )
   );



typedef struct packed {
  
 struct packed {
         logic        q;
       } txunderflow;
   } spi_device_reg2hw_intr_enable_reg_t;

   function automatic logic [31:0] prince_shiftrows_32bit(logic [31:0]      state_in,
                                                               logic [15:0][3:0] shifts );
    
   endfunction : prince_shiftrows_32bit

endmodule : toto
