/*
:name: class_member_test_9
:description: Test
:tags: 8.3
*/
class myclass;
extern local static task subtask(arg_type arg);
endclass