/*
:name: integers-token
:description: Testing the integer variable type
:should_fail: 0
:tags: 5.7.1
*/
module top();
  integer a;
endmodule
