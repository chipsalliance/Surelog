/*
:name: string_atoi
:description: string.atoi()  tests
:tags: 6.16.9
*/
module top();
	string a = "1234";
	int b = a.atoi();
endmodule
