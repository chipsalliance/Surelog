/*
:name: typedef_test_14
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef some_package::some_type myalias;