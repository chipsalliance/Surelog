
module dut ();

parameter S = $size(int);

initial begin
  $display();
end

class A;
endclass
   
endmodule
