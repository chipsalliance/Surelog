
`ifndef BP_FE_LCE_VH
`define BP_FE_LCE_VH

`include "bp_common_me_if.vh"

`endif
