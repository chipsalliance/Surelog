package toto1;





class blah1;
endclass












class blah2;
endclass















class blah3;
endclass








endpackage




package toto2;





class blah21;
endclass




class blah22;
endclass




endpackage



module inb ();
endmodule


package toto3;


endpackage

module gap2();
endmodule





























module gap3();
endmodule


package toto4;

class blah31;
endclass












class blah31;
endclass















class blah32;
endclass













class blah31_167;
endclass





endpackage






module gap4_181();












endmodule
