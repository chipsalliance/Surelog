/*
:name: typedef_test_9
:description: Test
:tags: 6.18
*/
parameter j = 3;
parameter k = 2;
typedef bit data_t;

typedef data_t my_array_t [k:0][j:0];
