module dut (a, b);

   function void UVMC_set_config_object (string type_name,
      string contxt,
      string inst_name,
      string field_name,
      bits_t value);
typedef uvmc_default_converter #(uvm_object) converter1;
typedef logic converter2;

uvm_object obj;
uvm_component comp;


   endfunction


 endmodule
 
