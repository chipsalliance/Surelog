module spidpi();
  import "DPI-C" function
    byte tick(input [1:0] d2p_data);
endmodule
