/*
:name: 22.8--default_nettype-redefinition
:description: Test
:tags: 22.8
:type: preprocessing
*/
`default_nettype wire
`default_nettype tri
`default_nettype tri0
`default_nettype tri1
`default_nettype wand
`default_nettype triand
`default_nettype wor
`default_nettype trior
`default_nettype trireg
`default_nettype uwire
`default_nettype none
