/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 3276
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_clkmux_3to1_diff_slvt_tb
// Design view name: config_vlog
// Solver: Spectre

// Library - wphy_gf12lp_ips_lib, Cell - wphy_clkmux_3to1_diff_slvt,
//View - schematic
// LAST TIME SAVED: May 10 06:34:49 2021
// NETLIST TIME: May 18 22:45:57 2021
`timescale 1ps / 1ps

`endif //SYNTHESIS
module wphy_clkmux_3to1_diff_slvt (out_c, out_t,   in01_c,
    in01_t, in10_c, in10_t, in11_c, in11_t, s
`ifdef WLOGIC_NO_PG
`else
 ,vdda
 ,vss
`endif //WLOGIC_NO_PG
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif

output  out_c, out_t;

input  in01_c, in01_t, in10_c, in10_t, in11_c, in11_t;

input [1:0]  s;

// Buses in the design
`ifdef SYNTHESIS
`else

wire  [1:0]  sb;

wire  [1:0]  s_buf;

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV1_1 ( .in(mux_slw_tb), .vss(vss), .out(c1),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV1_0 ( .in(mux_slw_tb), .vss(vss), .out(c1),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV0_1 ( .in(mux_slw_cb), .vss(vss), .out(t1),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV0_0 ( .in(mux_slw_cb), .vss(vss), .out(t1),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_0 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_1 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_2 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_3 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_4 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_5 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_6 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV8_7 ( .in(yb_t), .vss(vss), .out(out_t),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV7 ( .in(s00b), .vss(vss), .out(s00), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV5_1 ( .in(s[1]), .vss(vss), .out(sb[1]),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV5_0 ( .in(s[0]), .vss(vss), .out(sb[0]),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV6_1 ( .in(sb[1]), .vss(vss), .out(s_buf[1]),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV6_0 ( .in(sb[0]), .vss(vss), .out(s_buf[0]),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV4 ( .in(s01b), .vss(vss), .out(s01), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV3 ( .in(s10b), .vss(vss), .out(s10), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV2 ( .in(s11b), .vss(vss), .out(s11), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_0 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_1 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_2 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_3 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_4 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_5 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_6 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT INV9_7 ( .in(yb_c), .vss(vss), .out(out_c),
    .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_PDDUM_D2_GL16_SLVT PDDUM ( .vss(vss), .tielo(vss));

wphy_clkmux_3to1_diff_slvt_NAND2_D1_GL16_SLVT NAND3 ( .y(s00b), .b(sb[0]), .a(sb[1]), .tielo(vss),
    .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_slvt_NAND2_D1_GL16_SLVT NAND2 ( .y(s10b), .b(sb[0]), .a(s_buf[1]),
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_slvt_NAND2_D1_GL16_SLVT NAND1 ( .y(s11b), .b(s_buf[0]), .a(s_buf[1]),
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_slvt_NAND2_D1_GL16_SLVT NAND0 ( .y(s01b), .b(s_buf[0]), .a(sb[1]),
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT3 ( .out(mux_slw_tb), .en(s11), .enb(s11b),
    .vss(vss), .in(in11_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT03 ( .out(mux_slw_cb), .en(s11), .enb(s11b),
    .vss(vss), .in(in11_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT02 ( .out(mux_slw_cb), .en(s10), .enb(s10b),
    .vss(vss), .in(in10_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT4_3 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(t1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT4_2 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(t1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT4_1 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(t1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT4_0 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(t1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT2 ( .out(mux_slw_tb), .en(s10), .enb(s10b),
    .vss(vss), .in(in10_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT1_3 ( .out(yb_c), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT1_2 ( .out(yb_c), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT1_1 ( .out(yb_c), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT1_0 ( .out(yb_c), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT5_3 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(c1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT5_2 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(c1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT5_1 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(c1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT5_0 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]),
    .vss(vss), .in(c1), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT01_3 ( .out(yb_t), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT01_2 ( .out(yb_t), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT01_1 ( .out(yb_t), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT INVT01_0 ( .out(yb_t), .en(s01), .enb(s01b),
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_slvt_PD_D2_GL16_SLVT PD0 ( .vss(vss), .enb(s00), .y(yb_c));

wphy_clkmux_3to1_diff_slvt_PU_D2_GL16_SLVT PU0 ( .vdd(vdda), .en(s00b), .y(yb_t));

wphy_clkmux_3to1_diff_slvt_PUDUM_D2_GL16_SLVT PUDUM ( .vdd(vdda), .tiehi(vdda));

`ifdef WPHY_ANA_TIMING

specify

  if (s==='b01) (in01_t => out_t) = 13;
  if (s==='b10) (in10_t => out_t) = 19;
  if (s==='b11) (in11_t => out_t) = 19;

endspecify

`endif

`endif //SYNTHESIS
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell -
//wphy_clkmux_3to1_diff_slvt_tb, View - schematic
// LAST TIME SAVED: May 18 22:36:33 2021
// NETLIST TIME: May 18 22:45:57 2021
`timescale 1ps / 1ps

 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_gf12lp_dig_lib", "wphy_clkmux_3to1_diff_slvt_PUDUM_D2_GL16_SLVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_PUDUM_D2_GL16_SLVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  input tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_gf12lp_dig_lib", "wphy_clkmux_3to1_diff_slvt_PU_D2_GL16_SLVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_PU_D2_GL16_SLVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;

  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_gf12lp_dig_lib", "wphy_clkmux_3to1_diff_slvt_PD_D2_GL16_SLVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_PD_D2_GL16_SLVT ( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;

  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "INVT_D2_GL16_LVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_INVT_D2_GL16_SLVT( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

assign out = (en) ? ~in:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "NAND2_D1_GL16_LVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_NAND2_D1_GL16_SLVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_gf12lp_dig_lib", "wphy_clkmux_3to1_diff_slvt_PDDUM_D2_GL16_SLVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_PDDUM_D2_GL16_SLVT ( tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "INV_D2_GL16_LVT" "systemVerilog"

module wphy_clkmux_3to1_diff_slvt_INV_D2_GL16_SLVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
`endif //SYNTHESIS
