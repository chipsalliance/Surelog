/*
:name: class_member_test_13
:description: Test
:should_fail: 0
:tags: 8.3
*/
class protected_stuff;
  protected int count;
  protected const int countess = `SSS;
  protected var int counter = 0;
  protected const var int counted = 1;
  protected const myclass::msg_t null_msg = {1'b1, 1'b0};
endclass