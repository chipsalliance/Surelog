//===================================================================
//
// Copyright (C) Wavious 2020 - All Rights Reserved
//
// Unauthorized copying of this file, via any medium is strictly prohibited
//
// Created by sbridges on April/19/2020 at 10:03:15
//
// wav_reg_model_mvp_pll_no_reg_test.svh
//
//===================================================================






