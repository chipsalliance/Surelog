
module top;
    logic [63:0] sxc;

    assign sxc = 'x << 8;
   
endmodule