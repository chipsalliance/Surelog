/*
:name: 22.7--timescale-basic-2
:description: Test
:tags: 22.7
:type: preprocessing
*/
`timescale 10 us / 100 ns
