// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: nettype
:description: user-defined nettype tests
:tags: 6.6.7
*/
module top();
	nettype real real_net;
endmodule
