module top();
function func;
        localparam FUNC_LOCALPARAM = 32 - 1;
        parameter FUNC_PARAMETER = 1 - 0;
endfunction
endmodule
