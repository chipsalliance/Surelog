/*
:name: empty_test_0
:description: Test
:type: preprocessing
:tags: 5.3 5.4
*/
