`define DDR_CMN_PLL_EN_FIELD                                    0:0
`define DDR_CMN_PLL_BIAS_LVL_FIELD                              4:1
`define DDR_CMN_PLL_VCO0_FINE_FIELD                             10:5
`define DDR_CMN_PLL_INT_CTRL_FIELD                              15:11
`define DDR_CMN_PLL_CP_INT_MODE_FIELD                           16:16
`define DDR_CMN_PLL_VCO1_FINE_FIELD                             22:17
`define DDR_CMN_PLL_VCO2_FINE_FIELD                             28:23
`define DDR_CMN_PLL_PROP_CTRL_FIELD                             33:29
`define DDR_CMN_PLL_PROP_R_CTRL_FIELD                           35:34
`define DDR_CMN_PLL_PROP_C_CTRL_FIELD                           37:36
`define DDR_CMN_PLL_VCO1_ENA_FIELD                              38:38
`define DDR_CMN_PLL_VCO1_BAND_FIELD                             44:39
`define DDR_CMN_PLL_VCO1_POST_DIV_FIELD                         46:45
`define DDR_CMN_PLL_VCO1_BYP_CLK_SEL_FIELD                      47:47
`define DDR_CMN_PLL_VCO2_ENA_FIELD                              48:48
`define DDR_CMN_PLL_VCO2_BAND_FIELD                             54:49
`define DDR_CMN_PLL_VCO2_POST_DIV_FIELD                         56:55
`define DDR_CMN_PLL_VCO2_BYP_CLK_SEL_FIELD                      57:57
`define DDR_CMN_PLL_VCO_SEL_FIELD                               59:58
`define DDR_CMN_PLL_PFD_MODE_FIELD                              61:60
`define DDR_CMN_PLL_SEL_REFCLK_ALT_FIELD                        62:62
`define DDR_CMN_PLL_FBDIV_SEL_FIELD                             71:63
`define DDR_CMN_PLL_VCO0_ENA_FIELD                              72:72
`define DDR_CMN_PLL_VCO0_BAND_FIELD                             78:73
`define DDR_CMN_PLL_VCO0_BYP_CLK_SEL_FIELD                      79:79
`define DDR_CMN_PLL_DIV16_EN_FIELD                              80:80
//`define DDR_CMN_PLL_BIAS_SEL_FIELD                              81:81
`define DDR_CMN_PLL_CFG_BUS_WIDTH                               81
`define DDR_CMN_PLL_CFG_BUS_RANGE                               80:0
