/*
:name: shortreal
:description: shortreal type tests
:tags: 6.12
*/
module top();
	shortreal a = 0.5;
endmodule
