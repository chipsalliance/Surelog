/*
:name: memories-basic
:description: Test memories support
:tags: 7.4.4
*/
module top ();

// one-dimensinal array with elements of types
// reg, logic, bit
logic [7:0] mem [0:255];

endmodule
