`define DDR_ANA_DQS_DRVR_LPBK_OVRD_SEL_FIELD       2:0
`define DDR_ANA_DQS_DRVR_LPBK_OVRD_VAL_C_FIELD       3
`define DDR_ANA_DQS_DRVR_LPBK_OVRD_VAL_T_FIELD       4
`define DDR_ANA_DQS_DRVR_LPBK_SW_OVR_FIELD           5
`define DDR_ANA_DQS_DRVR_LPBK_TX_IMPD_FIELD        8:6
`define DDR_ANA_DQS_DRVR_LPBK_RX_IMPD_FIELD       11:9
