/*
:name: string-broken-line
:description: Basic broken line string example
:tags: 5.9
*/
module top();

  initial begin;
    $display("broken \
              line");
  end

endmodule
