module bot ();
sub sub1();
sub sub2();
endmodule

