/*
:name: 22.10--celldefine-basic-2
:description: Test
:should_fail: 0
:tags: 22.10
:type: preprocessing
*/
`celldefine
