module top;
   export "DPI-C" task simutil_memload;
   task simutil_memload;
      input string file;
   endtask
endmodule // top
