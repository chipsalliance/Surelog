/*
Bar.vh
*/

