/*
:name: class_member_test_46
:description: Test
:tags: 8.3
*/
class constructible;
extern function new(string name, int count);
endclass