/*
:name: class_member_test_11
:description: Test
:tags: 8.3
*/
class myclass;
  int buzz_count;
endclass