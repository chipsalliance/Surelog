module DFlipflop8Bit(A1, Q1, A2, Q2);

output reg [7:0] Q1;
input wire [7:0] A1;

output  [7:0] Q2;
input  [7:0] A2;

endmodule


module DFlipflop8Bit2(input [7:0] A3, 
                      input wire [7:0] A4, 
                      output [7:0] Q3, 
                      output reg [7:0] Q4);

endmodule
