/*
:name: info_task
:description: $info test
:should_fail: 0
:tags: 20.10
:type: simulation parsing
*/

module top();

initial begin
	$info("info");
end

endmodule
