/*
:name: class_member_test_49
:description: Test
:tags: 8.3
*/
class myclass;
virtual splinterface grinterface, winterface;
virtual interface foo_if bar_if, baz_if;
endclass