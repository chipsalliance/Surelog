/*
:name: string_itoa
:description: string.itoa()  tests
:tags: 6.16.11
*/
module top();
	string a;
	initial
		a.itoa(12);
endmodule
