module a(
input interconnect b,
input interconnect [2:0] c
	);
interconnect d;
interconnect [1:0] e;
interconnect [4:0] f [5:0];
endmodule


