/*
:name: 22.9--unconnected_drive-invalid-3
:description: Test
:should_fail_because: `nounconnected_drive takes no argument
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull0
`nounconnected_drive pull0
