/*
:name: event
:description: event type tests
:should_fail: 0
:tags: 6.17
*/
module top();
	event a;
endmodule
