
`ifndef BP_COMMON_ME_IF_VH
`define BP_COMMON_ME_IF_VH

typedef enum bit [2:0] 
{
  e_lce_cce_sync_ack         = 3'b000
  ,e_lce_cce_inv_ack         = 3'b001
} bp_lce_cce_resp_type_e;


`endif
