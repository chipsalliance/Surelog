
module prim_pad_wrapper

  #(
  
    parameter int signed AttrDw = 6
  
  ) ();

endmodule // prim_pad_wrapper
