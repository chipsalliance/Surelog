/*
:name: typedef_test_0
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef i_am_a_type_really;