/*
:name: typedef_test_21
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef enum bit[3:0] {
  Global = 4'h2,
  Local = 4'h3
} myenum_fwd;
