`define DDR_CSP_PRECLKDIS_WAIT_FIELD                      3:0
`define DDR_CSP_PRERST_WAIT_FIELD                         7:4
`define DDR_CSP_RST_PULSE_WIDTH_FIELD                     11:8
`define DDR_CSP_PSTRST_WAIT_FIELD                         15:12
`define DDR_CSP_PSTCLKEN_WAIT_FIELD                       19:16
`define DDR_CSP_PSTPIEN_WAIT_FIELD                        23:20
`define DDR_CSP_REQ_COMPLETE_OVR_SEL_FIELD                24:24
`define DDR_CSP_REQ_COMPLETE_OVR_FIELD                    25:25
`define DDR_CSP_REQ_OVR_SEL_FIELD                         26:26
`define DDR_CSP_REQ_OVR_FIELD                             27:27
`define DDR_CSP_CGC_EN_OVR_FIELD                          28:28
`define DDR_CSP_PI_DISABLE_OVR_FIELD                      29:29
`define DDR_CSP_DIV_RST_OVR_FIELD                         30:30
`define DDR_CSP_CLK_DISABLE_OVR_FIELD                     31:31

`define DDR_CSP_CFG_BUS_WIDTH           32
`define DDR_CSP_CFG_BUS_RANGE           31:0
