/*
:name: iface_class_test_1
:description: Test
:should_fail: 0
:tags: 8.3 8.26
*/
interface class base_ic;
endclass : base_ic