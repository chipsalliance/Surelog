/*
:name: empty_test_4
:description: Test
:type: preprocessing
:tags: 5.3 5.4
*/
// comment
