module top();
   import pkg2::*;
   
endmodule
