/*
:name: enum_anon
:description: anonymous enum tests
:should_fail: 0
:tags: 6.19
*/
module top();
	enum {a, b, c} val;
endmodule
