/*
:name: string_atoreal
:description: string.atoreal()  tests
:tags: 6.16.10
*/
module top();
	string a = "4.76";
	real b = a.atoreal();
endmodule
