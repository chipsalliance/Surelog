// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: typedef_test_8
:description: Test
:tags: 6.18
*/
typedef bit some_other_type;
typedef some_other_type myalias;

module test;
endmodule
