/*
:name: class_test_23
:description: Test
:tags: 6.15 8.3
*/
class Foo implements Bar; endclass