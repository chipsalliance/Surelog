module a;assign a = 0'sh0;
endmodule

