module minimal;
reg [7:0] q;
initial begin
q <= '81;
end
endmodule
