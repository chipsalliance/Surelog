/*
:name: class_test_61
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class pp_class;
`ifndef DEBUGGER
`endif
endclass