// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: info_task
:description: $info test
:tags: 20.10
:type: simulation parsing
*/

module top();

initial begin
	$info("info");
end

endmodule
