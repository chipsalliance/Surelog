/*
:name: desc_test_18
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifndef ASIC_OR_FPGA
`else
module module_asic;
endmodule
module module_fpga;
endmodule
`endif
