/*
:name: preproc_test_4
:description: Test
:should_fail: 0
:tags: 5.6.4
:type: preprocessing
*/
`ifdef INSANITY
`define INSANITY // comment
`else
`define SANITY 1
`endif
