/*
:name: non_blocking_assignment
:description: non-blocking assignment test
:tags: 10.4.2
*/
module top();

logic a;

initial begin
	a <= 2;
end

endmodule
