
module dut ();

parameter S = $size(int);

initial begin
  $display();
end

endmodule
