/*
:name: 22.5.2--undef-basic
:description: Test
:tags: 22.5.2
:type: preprocessing
*/
`define FOO "foo"
`undef FOO
