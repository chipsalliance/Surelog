package p;

parameter package_param = 1;
struct { 
  int x; 
} s1;

struct { 
int x; 
} s2;

function
void f();
int x;
endfunction

endpackage


package q;

parameter package_para = 1;
struct { 
  int x; 
} s1;

struct { 
int x; 
} s2;

function
void f();
int x;
endfunction

endpackage



package r;

parameter package_para = 1;
struct { 
  int x; 
} s1;

struct { 
int x; 
} s2;

function
void f();
int x;
endfunction

endpackage



package s;

parameter package_para = 1;
struct { 
  int x; 
} s1;

struct { 
int x; 
} s2;

function
void f();
int x;
endfunction

endpackage




