/*
:name: variable_assignment
:description: Variable assignment tests
:tags: 6.5
*/
module top();
	int v;

	assign v = 12;
endmodule
