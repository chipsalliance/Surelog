module top();
   assign oo = '{8:1};
   assign uu = '{8{1}};
endmodule
