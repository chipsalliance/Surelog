// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.9--unconnected_drive-basic
:description: Test
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull1
`nounconnected_drive
