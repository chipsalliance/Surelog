/*
:name: arrays-key-index
:description: Basic arrays test
:tags: 5.11
*/
module top();
  typedef int triple [1:3];
  triple b = '{1:1, default:0};
endmodule
