/*
:name: typedef_test_6
:description: Test
:tags: 6.18
*/
typedef struct { int i; bit b; } mystruct;
