/*
:name: real
:description: real type tests
:should_fail: 0
:tags: 6.12
*/
module top();
	real a = 0.5;
endmodule
