
nettype real my_real with my_function2;

function automatic real my_function2(input real driver []);
endfunction

