/*
:name: 22.5.2--undef-nonexisting
:description: Test
:should_fail: 0
:tags: 22.5.2
:type: preprocessing
*/
`undef FOO
`undef BAR
