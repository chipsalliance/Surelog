/*
:name: class_member_test_40
:description: Test
:tags: 8.3
*/
class constructible;
function new ();
endfunction
endclass