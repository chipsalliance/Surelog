/*
:name: class_test_5
:description: Test
:tags: 6.15 8.3
*/
virtual class automatic Foo; endclass