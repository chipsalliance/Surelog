/*
:name: desc_test_6
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
module mymod;
endmodule
`endif
