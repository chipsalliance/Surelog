module test(
  output logic [31:0] b
);

  assign b = '1;

endmodule
