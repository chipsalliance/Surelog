/*
:name: finish_task
:description: $finish test
:should_fail: 0
:tags: 20.2
*/
module top();

initial
	$finish;

endmodule
