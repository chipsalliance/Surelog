/*
:name: logic_vector
:description: logic vector tests
:should_fail: 0
:tags: 6.9.1
*/
module top();
	logic [15:0] a;
endmodule
