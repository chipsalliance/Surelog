module top;
   int dynamic [];
   int assoc [int];
   int assoc_string [string];
   int queue [$];
endmodule // top

