module foo;
  parameter int bar = 0;
endmodule

module baz;
endmodule // baz

