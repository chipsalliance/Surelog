/*
:name: iface_class_test_7
:description: Test
:should_fail: 0
:tags: 8.3 8.26
*/
interface class base_ic;
typedef struct { int i; bool b; } mystruct;
typedef enum { RED, GREEN, BLUE } colors;
typedef virtual blah_if harness_if;
typedef some_class#(3, 2, 1) car_type;
endclass