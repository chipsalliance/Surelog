/*
:name: stime_task
:description: $stime test
:tags: 20.3
*/
module top();

initial
	$display($stime);

endmodule
