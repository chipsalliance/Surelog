// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: system-functions
:description: Calling system functions
:tags: 5.6.3
*/
module systemfn();
  /* Note:
   * This does not test all the individual system calls.
   * It just verifies if the concept exists using one of the
   * calls.
   */

  initial $display("hello world");
endmodule
