/*
:name: basic-packed
:description: Test packed arrays support
:should_fail: 0
:tags: 7.4.1 7.4
*/
module top ();

bit [7:0] _bit;
logic [7:0] _logic;
reg [7:0] _reg;

endmodule
