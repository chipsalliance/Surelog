/*
:name: class_member_test_12
:description: Test
:should_fail: 0
:tags: 8.3
*/
class semaphore;
  local chandle p_handle;
endclass