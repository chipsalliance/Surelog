/*
:name: realtime_task
:description: $realtime test
:tags: 20.3
*/
module top();

initial
	$display($realtime);

endmodule
