`ifndef TVIP_AXI_RAL_PREDICTOR_SVH
`define TVIP_AXI_RAL_PREDICTOR_SVH
typedef tue_reg_predictor #(tvip_axi_item) tvip_axi_ral_predictor;
`endif
