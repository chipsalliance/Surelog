`define DDR_ANA_PI_CODE_RANGE                    5:0
`define DDR_ANA_PI_GEAR_RANGE                    9:6
`define DDR_ANA_PI_XCPL_RANGE                    13:10
`define DDR_ANA_PI_EN_RANGE                      14

`define DDR_ANA_PI_THERM_RANGE                   31:16
`define DDR_ANA_PI_QUAD_RANGE                    33:32

`define DDR_ANA_PI_ENC_RANGE                     14:0
`define DDR_ANA_PI_DEC_RANGE                     33:16
