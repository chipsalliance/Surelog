module top(input in,output out);
  SB_DFF dff(out,in,1);
endmodule
