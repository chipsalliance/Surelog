/*
:name: time_task
:description: $time test
:should_fail: 0
:tags: 20.3
*/
module top();

initial
	$display($time);

endmodule
