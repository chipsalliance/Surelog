module aes(clk, reset, load_i, decrypt_i, data_i, key_i, ready_o, data_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  wire _2214_;
  wire _2215_;
  wire _2216_;
  wire _2217_;
  wire _2218_;
  wire _2219_;
  wire _2220_;
  wire _2221_;
  wire _2222_;
  wire _2223_;
  wire _2224_;
  wire _2225_;
  wire _2226_;
  wire _2227_;
  wire _2228_;
  wire _2229_;
  wire _2230_;
  wire _2231_;
  wire _2232_;
  wire _2233_;
  wire _2234_;
  wire _2235_;
  wire _2236_;
  wire _2237_;
  wire _2238_;
  wire _2239_;
  wire _2240_;
  wire _2241_;
  wire _2242_;
  wire _2243_;
  wire _2244_;
  wire _2245_;
  wire _2246_;
  wire _2247_;
  wire _2248_;
  wire _2249_;
  wire _2250_;
  wire _2251_;
  wire _2252_;
  wire _2253_;
  wire _2254_;
  wire _2255_;
  wire _2256_;
  wire _2257_;
  wire _2258_;
  wire _2259_;
  wire _2260_;
  wire _2261_;
  wire _2262_;
  wire _2263_;
  wire _2264_;
  wire _2265_;
  wire _2266_;
  wire _2267_;
  wire _2268_;
  wire _2269_;
  wire _2270_;
  wire _2271_;
  wire _2272_;
  wire _2273_;
  wire _2274_;
  wire _2275_;
  wire _2276_;
  wire _2277_;
  wire _2278_;
  wire _2279_;
  wire _2280_;
  wire _2281_;
  wire _2282_;
  wire _2283_;
  wire _2284_;
  wire _2285_;
  wire _2286_;
  wire _2287_;
  wire _2288_;
  wire _2289_;
  wire _2290_;
  wire _2291_;
  wire _2292_;
  wire _2293_;
  wire _2294_;
  wire _2295_;
  wire _2296_;
  wire _2297_;
  wire _2298_;
  wire _2299_;
  wire _2300_;
  wire _2301_;
  wire _2302_;
  wire _2303_;
  wire _2304_;
  wire _2305_;
  wire _2306_;
  wire _2307_;
  wire _2308_;
  wire _2309_;
  wire _2310_;
  wire _2311_;
  wire _2312_;
  wire _2313_;
  wire _2314_;
  wire _2315_;
  wire _2316_;
  wire _2317_;
  wire _2318_;
  wire _2319_;
  wire _2320_;
  wire _2321_;
  wire _2322_;
  wire _2323_;
  wire _2324_;
  wire _2325_;
  wire _2326_;
  wire _2327_;
  wire _2328_;
  wire _2329_;
  wire _2330_;
  wire _2331_;
  wire _2332_;
  wire _2333_;
  wire _2334_;
  wire _2335_;
  wire _2336_;
  wire _2337_;
  wire _2338_;
  wire _2339_;
  wire _2340_;
  wire _2341_;
  wire _2342_;
  wire _2343_;
  wire _2344_;
  wire _2345_;
  wire _2346_;
  wire _2347_;
  wire _2348_;
  wire _2349_;
  wire _2350_;
  wire _2351_;
  wire _2352_;
  wire _2353_;
  wire _2354_;
  wire _2355_;
  wire _2356_;
  wire _2357_;
  wire _2358_;
  wire _2359_;
  wire _2360_;
  wire _2361_;
  wire _2362_;
  wire _2363_;
  wire _2364_;
  wire _2365_;
  wire _2366_;
  wire _2367_;
  wire _2368_;
  wire _2369_;
  wire _2370_;
  wire _2371_;
  wire _2372_;
  wire _2373_;
  wire _2374_;
  wire _2375_;
  wire _2376_;
  wire _2377_;
  wire _2378_;
  wire _2379_;
  wire _2380_;
  wire _2381_;
  wire _2382_;
  wire _2383_;
  wire _2384_;
  wire _2385_;
  wire _2386_;
  wire _2387_;
  wire _2388_;
  wire _2389_;
  wire _2390_;
  wire _2391_;
  wire _2392_;
  wire _2393_;
  wire _2394_;
  wire _2395_;
  wire _2396_;
  wire _2397_;
  wire _2398_;
  wire _2399_;
  wire _2400_;
  wire _2401_;
  wire _2402_;
  wire _2403_;
  wire _2404_;
  wire _2405_;
  wire _2406_;
  wire _2407_;
  wire _2408_;
  wire _2409_;
  wire _2410_;
  wire _2411_;
  wire _2412_;
  wire _2413_;
  wire _2414_;
  wire _2415_;
  wire _2416_;
  wire _2417_;
  wire _2418_;
  wire _2419_;
  wire _2420_;
  wire _2421_;
  wire _2422_;
  wire _2423_;
  wire _2424_;
  wire _2425_;
  wire _2426_;
  wire _2427_;
  wire _2428_;
  wire _2429_;
  wire _2430_;
  wire _2431_;
  wire _2432_;
  wire _2433_;
  wire _2434_;
  wire _2435_;
  wire _2436_;
  wire _2437_;
  wire _2438_;
  wire _2439_;
  wire _2440_;
  wire _2441_;
  wire _2442_;
  wire _2443_;
  wire _2444_;
  wire _2445_;
  wire _2446_;
  wire _2447_;
  wire _2448_;
  wire _2449_;
  wire _2450_;
  wire _2451_;
  wire _2452_;
  wire _2453_;
  wire _2454_;
  wire _2455_;
  wire _2456_;
  wire _2457_;
  wire _2458_;
  wire _2459_;
  wire _2460_;
  wire _2461_;
  wire _2462_;
  wire _2463_;
  wire _2464_;
  wire _2465_;
  wire _2466_;
  wire _2467_;
  wire _2468_;
  wire _2469_;
  wire _2470_;
  wire _2471_;
  wire _2472_;
  wire _2473_;
  wire _2474_;
  wire _2475_;
  wire _2476_;
  wire _2477_;
  wire _2478_;
  wire _2479_;
  wire _2480_;
  wire _2481_;
  wire _2482_;
  wire _2483_;
  wire _2484_;
  wire _2485_;
  wire _2486_;
  wire _2487_;
  wire _2488_;
  wire _2489_;
  wire _2490_;
  wire _2491_;
  wire _2492_;
  wire _2493_;
  wire _2494_;
  wire _2495_;
  wire _2496_;
  wire _2497_;
  wire _2498_;
  wire _2499_;
  wire _2500_;
  wire _2501_;
  wire _2502_;
  wire _2503_;
  wire _2504_;
  wire _2505_;
  wire _2506_;
  wire _2507_;
  wire _2508_;
  wire _2509_;
  wire _2510_;
  wire _2511_;
  wire _2512_;
  wire _2513_;
  wire _2514_;
  wire _2515_;
  wire _2516_;
  wire _2517_;
  wire _2518_;
  wire _2519_;
  wire _2520_;
  wire _2521_;
  wire _2522_;
  wire _2523_;
  wire _2524_;
  wire _2525_;
  wire _2526_;
  wire _2527_;
  wire _2528_;
  wire _2529_;
  wire _2530_;
  wire _2531_;
  wire _2532_;
  wire _2533_;
  wire _2534_;
  wire _2535_;
  wire _2536_;
  wire _2537_;
  wire _2538_;
  wire _2539_;
  wire _2540_;
  wire _2541_;
  wire _2542_;
  wire _2543_;
  wire _2544_;
  wire _2545_;
  wire _2546_;
  wire _2547_;
  wire _2548_;
  wire _2549_;
  wire _2550_;
  wire _2551_;
  wire _2552_;
  wire _2553_;
  wire _2554_;
  wire _2555_;
  wire _2556_;
  wire _2557_;
  wire _2558_;
  wire _2559_;
  wire _2560_;
  wire _2561_;
  wire _2562_;
  wire _2563_;
  wire _2564_;
  wire _2565_;
  wire _2566_;
  wire _2567_;
  wire _2568_;
  wire _2569_;
  wire _2570_;
  wire _2571_;
  wire _2572_;
  wire _2573_;
  wire _2574_;
  wire _2575_;
  wire _2576_;
  wire _2577_;
  wire _2578_;
  wire _2579_;
  wire _2580_;
  wire _2581_;
  wire _2582_;
  wire _2583_;
  wire _2584_;
  wire _2585_;
  wire _2586_;
  wire _2587_;
  wire _2588_;
  wire _2589_;
  wire _2590_;
  wire _2591_;
  wire _2592_;
  wire _2593_;
  wire _2594_;
  wire _2595_;
  wire _2596_;
  wire _2597_;
  wire _2598_;
  wire _2599_;
  wire _2600_;
  wire _2601_;
  wire _2602_;
  wire _2603_;
  wire _2604_;
  wire _2605_;
  wire _2606_;
  wire _2607_;
  wire _2608_;
  wire _2609_;
  wire _2610_;
  wire _2611_;
  wire _2612_;
  wire _2613_;
  wire _2614_;
  wire _2615_;
  wire _2616_;
  wire _2617_;
  wire _2618_;
  wire _2619_;
  wire _2620_;
  wire _2621_;
  wire _2622_;
  wire _2623_;
  wire _2624_;
  wire _2625_;
  wire _2626_;
  wire _2627_;
  wire _2628_;
  wire _2629_;
  wire _2630_;
  wire _2631_;
  wire _2632_;
  wire _2633_;
  wire _2634_;
  wire _2635_;
  wire _2636_;
  wire _2637_;
  wire _2638_;
  wire _2639_;
  wire _2640_;
  wire _2641_;
  wire _2642_;
  wire _2643_;
  wire _2644_;
  wire _2645_;
  wire _2646_;
  wire _2647_;
  wire _2648_;
  wire _2649_;
  wire _2650_;
  wire _2651_;
  wire _2652_;
  wire _2653_;
  wire _2654_;
  wire _2655_;
  wire _2656_;
  wire _2657_;
  wire _2658_;
  wire _2659_;
  wire _2660_;
  wire _2661_;
  wire _2662_;
  wire _2663_;
  wire _2664_;
  wire _2665_;
  wire _2666_;
  wire _2667_;
  wire _2668_;
  wire _2669_;
  wire _2670_;
  wire _2671_;
  wire _2672_;
  wire _2673_;
  wire _2674_;
  wire _2675_;
  wire _2676_;
  wire _2677_;
  wire _2678_;
  wire _2679_;
  wire _2680_;
  wire _2681_;
  wire _2682_;
  wire _2683_;
  wire _2684_;
  wire _2685_;
  wire _2686_;
  wire _2687_;
  wire _2688_;
  wire _2689_;
  wire _2690_;
  wire _2691_;
  wire _2692_;
  wire _2693_;
  wire _2694_;
  wire _2695_;
  wire _2696_;
  wire _2697_;
  wire _2698_;
  wire _2699_;
  wire _2700_;
  wire _2701_;
  wire _2702_;
  wire _2703_;
  wire _2704_;
  wire _2705_;
  wire _2706_;
  wire _2707_;
  wire _2708_;
  wire _2709_;
  reg [127:0] addroundkey_data_o;
  wire [127:0] addroundkey_data_reg;
  reg addroundkey_ready_o;
  reg [3:0] addroundkey_round;
  reg addroundkey_start_i;
  input clk;
  input [127:0] data_i;
  output [127:0] data_o;
  input decrypt_i;
  reg first_round_reg;
  input [127:0] key_i;
  wire [127:0] keysched_last_key_i;
  wire [127:0] keysched_new_key_o;
  wire keysched_ready_o;
  wire [3:0] keysched_round_i;
  wire keysched_sbox_access_o;
  wire [7:0] keysched_sbox_data_o;
  wire keysched_sbox_decrypt_o;
  wire keysched_start_i;
  input load_i;
  wire [127:0] mixcol_data_i;
  wire [127:0] mixcol_data_o;
  wire mixcol_ready_o;
  wire mixcol_start_i;
  wire [127:0] next_addroundkey_data_reg;
  wire next_addroundkey_ready_o;
  wire [3:0] next_addroundkey_round;
  wire next_addroundkey_start_i;
  wire next_first_round_reg;
  wire next_ready_o;
  wire [3:0] next_round;
  wire next_state;
  output ready_o;
  reg ready_o;
  input reset;
  reg [3:0] round;
  wire [7:0] sbox_data_i;
  wire [7:0] sbox_data_o;
  wire sbox_decrypt_i;
  reg state;
  wire [127:0] subbytes_data_i;
  wire [127:0] subbytes_data_o;
  wire subbytes_ready_o;
  wire [7:0] subbytes_sbox_data_o;
  wire subbytes_sbox_decrypt_o;
  wire subbytes_start_i;
  assign _0000_ = round[1] | round[0];
  assign _0001_ = round[3] | round[2];
  assign _0002_ = _0001_ | _0000_;
  assign _0003_ = ~_0002_;
  assign _0004_ = _0003_ & addroundkey_start_i;
  assign _0005_ = ~addroundkey_round[1];
  assign _0006_ = _0005_ & addroundkey_round[0];
  assign _0007_ = ~addroundkey_round[2];
  assign _0008_ = ~addroundkey_round[3];
  assign _0009_ = _0008_ & _0007_;
  assign _0010_ = _0009_ & _0006_;
  assign _0011_ = ~addroundkey_round[0];
  assign _0012_ = _0005_ & _0011_;
  assign _0013_ = _0012_ & _0009_;
  assign _0014_ = _0013_ | _0010_;
  assign _0015_ = _0014_ ? key_i[0] : keysched_new_key_o[0];
  assign _0016_ = _0002_ & addroundkey_start_i;
  assign _0017_ = ~round[1];
  assign _0018_ = addroundkey_round[1] ^ _0017_;
  assign _0019_ = ~round[0];
  assign _0020_ = addroundkey_round[0] ^ _0019_;
  assign _0021_ = _0020_ & _0018_;
  assign _0022_ = ~round[3];
  assign _0023_ = addroundkey_round[3] ^ _0022_;
  assign _0024_ = ~round[2];
  assign _0025_ = addroundkey_round[2] ^ _0024_;
  assign _0026_ = _0025_ & _0023_;
  assign _0027_ = _0026_ & _0021_;
  assign _0028_ = ~_0027_;
  assign _0029_ = _0028_ & keysched_ready_o;
  assign _0030_ = _0029_ ? keysched_new_key_o[0] : _0015_;
  assign _0031_ = _0016_ ? key_i[0] : _0030_;
  assign keysched_last_key_i[0] = _0004_ ? _0015_ : _0031_;
  assign _0032_ = _0014_ ? key_i[100] : keysched_new_key_o[100];
  assign _0033_ = _0029_ ? keysched_new_key_o[100] : _0032_;
  assign _0034_ = _0016_ ? key_i[100] : _0033_;
  assign keysched_last_key_i[100] = _0004_ ? _0032_ : _0034_;
  assign _0035_ = _0014_ ? key_i[101] : keysched_new_key_o[101];
  assign _0036_ = _0029_ ? keysched_new_key_o[101] : _0035_;
  assign _0037_ = _0016_ ? key_i[101] : _0036_;
  assign keysched_last_key_i[101] = _0004_ ? _0035_ : _0037_;
  assign _0038_ = _0014_ ? key_i[102] : keysched_new_key_o[102];
  assign _0039_ = _0029_ ? keysched_new_key_o[102] : _0038_;
  assign _0040_ = _0016_ ? key_i[102] : _0039_;
  assign keysched_last_key_i[102] = _0004_ ? _0038_ : _0040_;
  assign _0041_ = _0014_ ? key_i[103] : keysched_new_key_o[103];
  assign _0042_ = _0029_ ? keysched_new_key_o[103] : _0041_;
  assign _0043_ = _0016_ ? key_i[103] : _0042_;
  assign keysched_last_key_i[103] = _0004_ ? _0041_ : _0043_;
  assign _0044_ = _0014_ ? key_i[104] : keysched_new_key_o[104];
  assign _0045_ = _0029_ ? keysched_new_key_o[104] : _0044_;
  assign _0046_ = _0016_ ? key_i[104] : _0045_;
  assign keysched_last_key_i[104] = _0004_ ? _0044_ : _0046_;
  assign _0047_ = _0014_ ? key_i[105] : keysched_new_key_o[105];
  assign _0048_ = _0029_ ? keysched_new_key_o[105] : _0047_;
  assign _0049_ = _0016_ ? key_i[105] : _0048_;
  assign keysched_last_key_i[105] = _0004_ ? _0047_ : _0049_;
  assign _0050_ = _0014_ ? key_i[106] : keysched_new_key_o[106];
  assign _0051_ = _0029_ ? keysched_new_key_o[106] : _0050_;
  assign _0052_ = _0016_ ? key_i[106] : _0051_;
  assign keysched_last_key_i[106] = _0004_ ? _0050_ : _0052_;
  assign _0053_ = _0014_ ? key_i[107] : keysched_new_key_o[107];
  assign _0054_ = _0029_ ? keysched_new_key_o[107] : _0053_;
  assign _0055_ = _0016_ ? key_i[107] : _0054_;
  assign keysched_last_key_i[107] = _0004_ ? _0053_ : _0055_;
  assign _0056_ = _0014_ ? key_i[108] : keysched_new_key_o[108];
  assign _0057_ = _0029_ ? keysched_new_key_o[108] : _0056_;
  assign _0058_ = _0016_ ? key_i[108] : _0057_;
  assign keysched_last_key_i[108] = _0004_ ? _0056_ : _0058_;
  assign _0059_ = _0014_ ? key_i[109] : keysched_new_key_o[109];
  assign _0060_ = _0029_ ? keysched_new_key_o[109] : _0059_;
  assign _0061_ = _0016_ ? key_i[109] : _0060_;
  assign keysched_last_key_i[109] = _0004_ ? _0059_ : _0061_;
  assign _0062_ = _0014_ ? key_i[10] : keysched_new_key_o[10];
  assign _0063_ = _0029_ ? keysched_new_key_o[10] : _0062_;
  assign _0064_ = _0016_ ? key_i[10] : _0063_;
  assign keysched_last_key_i[10] = _0004_ ? _0062_ : _0064_;
  assign _0065_ = _0014_ ? key_i[110] : keysched_new_key_o[110];
  assign _0066_ = _0029_ ? keysched_new_key_o[110] : _0065_;
  assign _0067_ = _0016_ ? key_i[110] : _0066_;
  assign keysched_last_key_i[110] = _0004_ ? _0065_ : _0067_;
  assign _0068_ = _0014_ ? key_i[111] : keysched_new_key_o[111];
  assign _0069_ = _0029_ ? keysched_new_key_o[111] : _0068_;
  assign _0070_ = _0016_ ? key_i[111] : _0069_;
  assign keysched_last_key_i[111] = _0004_ ? _0068_ : _0070_;
  assign _0071_ = _0014_ ? key_i[112] : keysched_new_key_o[112];
  assign _0072_ = _0029_ ? keysched_new_key_o[112] : _0071_;
  assign _0073_ = _0016_ ? key_i[112] : _0072_;
  assign keysched_last_key_i[112] = _0004_ ? _0071_ : _0073_;
  assign _0074_ = _0014_ ? key_i[113] : keysched_new_key_o[113];
  assign _0075_ = _0029_ ? keysched_new_key_o[113] : _0074_;
  assign _0076_ = _0016_ ? key_i[113] : _0075_;
  assign keysched_last_key_i[113] = _0004_ ? _0074_ : _0076_;
  assign _0077_ = _0014_ ? key_i[114] : keysched_new_key_o[114];
  assign _0078_ = _0029_ ? keysched_new_key_o[114] : _0077_;
  assign _0079_ = _0016_ ? key_i[114] : _0078_;
  assign keysched_last_key_i[114] = _0004_ ? _0077_ : _0079_;
  assign _0080_ = _0014_ ? key_i[115] : keysched_new_key_o[115];
  assign _0081_ = _0029_ ? keysched_new_key_o[115] : _0080_;
  assign _0082_ = _0016_ ? key_i[115] : _0081_;
  assign keysched_last_key_i[115] = _0004_ ? _0080_ : _0082_;
  assign _0083_ = _0014_ ? key_i[116] : keysched_new_key_o[116];
  assign _0084_ = _0029_ ? keysched_new_key_o[116] : _0083_;
  assign _0085_ = _0016_ ? key_i[116] : _0084_;
  assign keysched_last_key_i[116] = _0004_ ? _0083_ : _0085_;
  assign _0086_ = _0014_ ? key_i[117] : keysched_new_key_o[117];
  assign _0087_ = _0029_ ? keysched_new_key_o[117] : _0086_;
  assign _0088_ = _0016_ ? key_i[117] : _0087_;
  assign keysched_last_key_i[117] = _0004_ ? _0086_ : _0088_;
  assign _0089_ = _0014_ ? key_i[118] : keysched_new_key_o[118];
  assign _0090_ = _0029_ ? keysched_new_key_o[118] : _0089_;
  assign _0091_ = _0016_ ? key_i[118] : _0090_;
  assign keysched_last_key_i[118] = _0004_ ? _0089_ : _0091_;
  assign _0092_ = _0014_ ? key_i[119] : keysched_new_key_o[119];
  assign _0093_ = _0029_ ? keysched_new_key_o[119] : _0092_;
  assign _0094_ = _0016_ ? key_i[119] : _0093_;
  assign keysched_last_key_i[119] = _0004_ ? _0092_ : _0094_;
  assign _0095_ = _0014_ ? key_i[11] : keysched_new_key_o[11];
  assign _0096_ = _0029_ ? keysched_new_key_o[11] : _0095_;
  assign _0097_ = _0016_ ? key_i[11] : _0096_;
  assign keysched_last_key_i[11] = _0004_ ? _0095_ : _0097_;
  assign _0098_ = _0014_ ? key_i[120] : keysched_new_key_o[120];
  assign _0099_ = _0029_ ? keysched_new_key_o[120] : _0098_;
  assign _0100_ = _0016_ ? key_i[120] : _0099_;
  assign keysched_last_key_i[120] = _0004_ ? _0098_ : _0100_;
  assign _0101_ = _0014_ ? key_i[121] : keysched_new_key_o[121];
  assign _0102_ = _0029_ ? keysched_new_key_o[121] : _0101_;
  assign _0103_ = _0016_ ? key_i[121] : _0102_;
  assign keysched_last_key_i[121] = _0004_ ? _0101_ : _0103_;
  assign _0104_ = _0014_ ? key_i[122] : keysched_new_key_o[122];
  assign _0105_ = _0029_ ? keysched_new_key_o[122] : _0104_;
  assign _0106_ = _0016_ ? key_i[122] : _0105_;
  assign keysched_last_key_i[122] = _0004_ ? _0104_ : _0106_;
  assign _0107_ = _0014_ ? key_i[123] : keysched_new_key_o[123];
  assign _0108_ = _0029_ ? keysched_new_key_o[123] : _0107_;
  assign _0109_ = _0016_ ? key_i[123] : _0108_;
  assign keysched_last_key_i[123] = _0004_ ? _0107_ : _0109_;
  assign _0110_ = _0014_ ? key_i[124] : keysched_new_key_o[124];
  assign _0111_ = _0029_ ? keysched_new_key_o[124] : _0110_;
  assign _0112_ = _0016_ ? key_i[124] : _0111_;
  assign keysched_last_key_i[124] = _0004_ ? _0110_ : _0112_;
  assign _0113_ = _0014_ ? key_i[125] : keysched_new_key_o[125];
  assign _0114_ = _0029_ ? keysched_new_key_o[125] : _0113_;
  assign _0115_ = _0016_ ? key_i[125] : _0114_;
  assign keysched_last_key_i[125] = _0004_ ? _0113_ : _0115_;
  assign _0116_ = _0014_ ? key_i[126] : keysched_new_key_o[126];
  assign _0117_ = _0029_ ? keysched_new_key_o[126] : _0116_;
  assign _0118_ = _0016_ ? key_i[126] : _0117_;
  assign keysched_last_key_i[126] = _0004_ ? _0116_ : _0118_;
  assign _0119_ = _0014_ ? key_i[127] : keysched_new_key_o[127];
  assign _0120_ = _0029_ ? keysched_new_key_o[127] : _0119_;
  assign _0121_ = _0016_ ? key_i[127] : _0120_;
  assign keysched_last_key_i[127] = _0004_ ? _0119_ : _0121_;
  assign _0122_ = _0014_ ? key_i[12] : keysched_new_key_o[12];
  assign _0123_ = _0029_ ? keysched_new_key_o[12] : _0122_;
  assign _0124_ = _0016_ ? key_i[12] : _0123_;
  assign keysched_last_key_i[12] = _0004_ ? _0122_ : _0124_;
  assign _0125_ = _0014_ ? key_i[13] : keysched_new_key_o[13];
  assign _0126_ = _0029_ ? keysched_new_key_o[13] : _0125_;
  assign _0127_ = _0016_ ? key_i[13] : _0126_;
  assign keysched_last_key_i[13] = _0004_ ? _0125_ : _0127_;
  assign _0128_ = _0014_ ? key_i[14] : keysched_new_key_o[14];
  assign _0129_ = _0029_ ? keysched_new_key_o[14] : _0128_;
  assign _0130_ = _0016_ ? key_i[14] : _0129_;
  assign keysched_last_key_i[14] = _0004_ ? _0128_ : _0130_;
  assign _0131_ = _0014_ ? key_i[15] : keysched_new_key_o[15];
  assign _0132_ = _0029_ ? keysched_new_key_o[15] : _0131_;
  assign _0133_ = _0016_ ? key_i[15] : _0132_;
  assign keysched_last_key_i[15] = _0004_ ? _0131_ : _0133_;
  assign _0134_ = _0014_ ? key_i[16] : keysched_new_key_o[16];
  assign _0135_ = _0029_ ? keysched_new_key_o[16] : _0134_;
  assign _0136_ = _0016_ ? key_i[16] : _0135_;
  assign keysched_last_key_i[16] = _0004_ ? _0134_ : _0136_;
  assign _0137_ = _0014_ ? key_i[17] : keysched_new_key_o[17];
  assign _0138_ = _0029_ ? keysched_new_key_o[17] : _0137_;
  assign _0139_ = _0016_ ? key_i[17] : _0138_;
  assign keysched_last_key_i[17] = _0004_ ? _0137_ : _0139_;
  assign _0140_ = _0014_ ? key_i[18] : keysched_new_key_o[18];
  assign _0141_ = _0029_ ? keysched_new_key_o[18] : _0140_;
  assign _0142_ = _0016_ ? key_i[18] : _0141_;
  assign keysched_last_key_i[18] = _0004_ ? _0140_ : _0142_;
  assign _0143_ = _0014_ ? key_i[19] : keysched_new_key_o[19];
  assign _0144_ = _0029_ ? keysched_new_key_o[19] : _0143_;
  assign _0145_ = _0016_ ? key_i[19] : _0144_;
  assign keysched_last_key_i[19] = _0004_ ? _0143_ : _0145_;
  assign _0146_ = _0014_ ? key_i[1] : keysched_new_key_o[1];
  assign _0147_ = _0029_ ? keysched_new_key_o[1] : _0146_;
  assign _0148_ = _0016_ ? key_i[1] : _0147_;
  assign keysched_last_key_i[1] = _0004_ ? _0146_ : _0148_;
  assign _0149_ = _0014_ ? key_i[20] : keysched_new_key_o[20];
  assign _0150_ = _0029_ ? keysched_new_key_o[20] : _0149_;
  assign _0151_ = _0016_ ? key_i[20] : _0150_;
  assign keysched_last_key_i[20] = _0004_ ? _0149_ : _0151_;
  assign _0152_ = _0014_ ? key_i[21] : keysched_new_key_o[21];
  assign _0153_ = _0029_ ? keysched_new_key_o[21] : _0152_;
  assign _0154_ = _0016_ ? key_i[21] : _0153_;
  assign keysched_last_key_i[21] = _0004_ ? _0152_ : _0154_;
  assign _0155_ = _0014_ ? key_i[22] : keysched_new_key_o[22];
  assign _0156_ = _0029_ ? keysched_new_key_o[22] : _0155_;
  assign _0157_ = _0016_ ? key_i[22] : _0156_;
  assign keysched_last_key_i[22] = _0004_ ? _0155_ : _0157_;
  assign _0158_ = _0014_ ? key_i[23] : keysched_new_key_o[23];
  assign _0159_ = _0029_ ? keysched_new_key_o[23] : _0158_;
  assign _0160_ = _0016_ ? key_i[23] : _0159_;
  assign keysched_last_key_i[23] = _0004_ ? _0158_ : _0160_;
  assign _0161_ = _0014_ ? key_i[24] : keysched_new_key_o[24];
  assign _0162_ = _0029_ ? keysched_new_key_o[24] : _0161_;
  assign _0163_ = _0016_ ? key_i[24] : _0162_;
  assign keysched_last_key_i[24] = _0004_ ? _0161_ : _0163_;
  assign _0164_ = _0014_ ? key_i[25] : keysched_new_key_o[25];
  assign _0165_ = _0029_ ? keysched_new_key_o[25] : _0164_;
  assign _0166_ = _0016_ ? key_i[25] : _0165_;
  assign keysched_last_key_i[25] = _0004_ ? _0164_ : _0166_;
  assign _0167_ = _0014_ ? key_i[26] : keysched_new_key_o[26];
  assign _0168_ = _0029_ ? keysched_new_key_o[26] : _0167_;
  assign _0169_ = _0016_ ? key_i[26] : _0168_;
  assign keysched_last_key_i[26] = _0004_ ? _0167_ : _0169_;
  assign _0170_ = _0014_ ? key_i[27] : keysched_new_key_o[27];
  assign _0171_ = _0029_ ? keysched_new_key_o[27] : _0170_;
  assign _0172_ = _0016_ ? key_i[27] : _0171_;
  assign keysched_last_key_i[27] = _0004_ ? _0170_ : _0172_;
  assign _0173_ = _0014_ ? key_i[28] : keysched_new_key_o[28];
  assign _0174_ = _0029_ ? keysched_new_key_o[28] : _0173_;
  assign _0175_ = _0016_ ? key_i[28] : _0174_;
  assign keysched_last_key_i[28] = _0004_ ? _0173_ : _0175_;
  assign _0176_ = _0014_ ? key_i[29] : keysched_new_key_o[29];
  assign _0177_ = _0029_ ? keysched_new_key_o[29] : _0176_;
  assign _0178_ = _0016_ ? key_i[29] : _0177_;
  assign keysched_last_key_i[29] = _0004_ ? _0176_ : _0178_;
  assign _0179_ = _0014_ ? key_i[2] : keysched_new_key_o[2];
  assign _0180_ = _0029_ ? keysched_new_key_o[2] : _0179_;
  assign _0181_ = _0016_ ? key_i[2] : _0180_;
  assign keysched_last_key_i[2] = _0004_ ? _0179_ : _0181_;
  assign _0182_ = _0014_ ? key_i[30] : keysched_new_key_o[30];
  assign _0183_ = _0029_ ? keysched_new_key_o[30] : _0182_;
  assign _0184_ = _0016_ ? key_i[30] : _0183_;
  assign keysched_last_key_i[30] = _0004_ ? _0182_ : _0184_;
  assign _0185_ = _0014_ ? key_i[31] : keysched_new_key_o[31];
  assign _0186_ = _0029_ ? keysched_new_key_o[31] : _0185_;
  assign _0187_ = _0016_ ? key_i[31] : _0186_;
  assign keysched_last_key_i[31] = _0004_ ? _0185_ : _0187_;
  assign _0188_ = _0014_ ? key_i[32] : keysched_new_key_o[32];
  assign _0189_ = _0029_ ? keysched_new_key_o[32] : _0188_;
  assign _0190_ = _0016_ ? key_i[32] : _0189_;
  assign keysched_last_key_i[32] = _0004_ ? _0188_ : _0190_;
  assign _0191_ = _0014_ ? key_i[33] : keysched_new_key_o[33];
  assign _0192_ = _0029_ ? keysched_new_key_o[33] : _0191_;
  assign _0193_ = _0016_ ? key_i[33] : _0192_;
  assign keysched_last_key_i[33] = _0004_ ? _0191_ : _0193_;
  assign _0194_ = _0014_ ? key_i[34] : keysched_new_key_o[34];
  assign _0195_ = _0029_ ? keysched_new_key_o[34] : _0194_;
  assign _0196_ = _0016_ ? key_i[34] : _0195_;
  assign keysched_last_key_i[34] = _0004_ ? _0194_ : _0196_;
  assign _0197_ = _0014_ ? key_i[35] : keysched_new_key_o[35];
  assign _0198_ = _0029_ ? keysched_new_key_o[35] : _0197_;
  assign _0199_ = _0016_ ? key_i[35] : _0198_;
  assign keysched_last_key_i[35] = _0004_ ? _0197_ : _0199_;
  assign _0200_ = _0014_ ? key_i[36] : keysched_new_key_o[36];
  assign _0201_ = _0029_ ? keysched_new_key_o[36] : _0200_;
  assign _0202_ = _0016_ ? key_i[36] : _0201_;
  assign keysched_last_key_i[36] = _0004_ ? _0200_ : _0202_;
  assign _0203_ = _0014_ ? key_i[37] : keysched_new_key_o[37];
  assign _0204_ = _0029_ ? keysched_new_key_o[37] : _0203_;
  assign _0205_ = _0016_ ? key_i[37] : _0204_;
  assign keysched_last_key_i[37] = _0004_ ? _0203_ : _0205_;
  assign _0206_ = _0014_ ? key_i[38] : keysched_new_key_o[38];
  assign _0207_ = _0029_ ? keysched_new_key_o[38] : _0206_;
  assign _0208_ = _0016_ ? key_i[38] : _0207_;
  assign keysched_last_key_i[38] = _0004_ ? _0206_ : _0208_;
  assign _0209_ = _0014_ ? key_i[39] : keysched_new_key_o[39];
  assign _0210_ = _0029_ ? keysched_new_key_o[39] : _0209_;
  assign _0211_ = _0016_ ? key_i[39] : _0210_;
  assign keysched_last_key_i[39] = _0004_ ? _0209_ : _0211_;
  assign _0212_ = _0014_ ? key_i[3] : keysched_new_key_o[3];
  assign _0213_ = _0029_ ? keysched_new_key_o[3] : _0212_;
  assign _0214_ = _0016_ ? key_i[3] : _0213_;
  assign keysched_last_key_i[3] = _0004_ ? _0212_ : _0214_;
  assign _0215_ = _0014_ ? key_i[40] : keysched_new_key_o[40];
  assign _0216_ = _0029_ ? keysched_new_key_o[40] : _0215_;
  assign _0217_ = _0016_ ? key_i[40] : _0216_;
  assign keysched_last_key_i[40] = _0004_ ? _0215_ : _0217_;
  assign _0218_ = _0014_ ? key_i[41] : keysched_new_key_o[41];
  assign _0219_ = _0029_ ? keysched_new_key_o[41] : _0218_;
  assign _0220_ = _0016_ ? key_i[41] : _0219_;
  assign keysched_last_key_i[41] = _0004_ ? _0218_ : _0220_;
  assign _0221_ = _0014_ ? key_i[42] : keysched_new_key_o[42];
  assign _0222_ = _0029_ ? keysched_new_key_o[42] : _0221_;
  assign _0223_ = _0016_ ? key_i[42] : _0222_;
  assign keysched_last_key_i[42] = _0004_ ? _0221_ : _0223_;
  assign _0224_ = _0014_ ? key_i[43] : keysched_new_key_o[43];
  assign _0225_ = _0029_ ? keysched_new_key_o[43] : _0224_;
  assign _0226_ = _0016_ ? key_i[43] : _0225_;
  assign keysched_last_key_i[43] = _0004_ ? _0224_ : _0226_;
  assign _0227_ = _0014_ ? key_i[44] : keysched_new_key_o[44];
  assign _0228_ = _0029_ ? keysched_new_key_o[44] : _0227_;
  assign _0229_ = _0016_ ? key_i[44] : _0228_;
  assign keysched_last_key_i[44] = _0004_ ? _0227_ : _0229_;
  assign _0230_ = _0014_ ? key_i[45] : keysched_new_key_o[45];
  assign _0231_ = _0029_ ? keysched_new_key_o[45] : _0230_;
  assign _0232_ = _0016_ ? key_i[45] : _0231_;
  assign keysched_last_key_i[45] = _0004_ ? _0230_ : _0232_;
  assign _0233_ = _0014_ ? key_i[46] : keysched_new_key_o[46];
  assign _0234_ = _0029_ ? keysched_new_key_o[46] : _0233_;
  assign _0235_ = _0016_ ? key_i[46] : _0234_;
  assign keysched_last_key_i[46] = _0004_ ? _0233_ : _0235_;
  assign _0236_ = _0014_ ? key_i[47] : keysched_new_key_o[47];
  assign _0237_ = _0029_ ? keysched_new_key_o[47] : _0236_;
  assign _0238_ = _0016_ ? key_i[47] : _0237_;
  assign keysched_last_key_i[47] = _0004_ ? _0236_ : _0238_;
  assign _0239_ = _0014_ ? key_i[48] : keysched_new_key_o[48];
  assign _0240_ = _0029_ ? keysched_new_key_o[48] : _0239_;
  assign _0241_ = _0016_ ? key_i[48] : _0240_;
  assign keysched_last_key_i[48] = _0004_ ? _0239_ : _0241_;
  assign _0242_ = _0014_ ? key_i[49] : keysched_new_key_o[49];
  assign _0243_ = _0029_ ? keysched_new_key_o[49] : _0242_;
  assign _0244_ = _0016_ ? key_i[49] : _0243_;
  assign keysched_last_key_i[49] = _0004_ ? _0242_ : _0244_;
  assign _0245_ = _0014_ ? key_i[4] : keysched_new_key_o[4];
  assign _0246_ = _0029_ ? keysched_new_key_o[4] : _0245_;
  assign _0247_ = _0016_ ? key_i[4] : _0246_;
  assign keysched_last_key_i[4] = _0004_ ? _0245_ : _0247_;
  assign _0248_ = _0014_ ? key_i[50] : keysched_new_key_o[50];
  assign _0249_ = _0029_ ? keysched_new_key_o[50] : _0248_;
  assign _0250_ = _0016_ ? key_i[50] : _0249_;
  assign keysched_last_key_i[50] = _0004_ ? _0248_ : _0250_;
  assign _0251_ = _0014_ ? key_i[51] : keysched_new_key_o[51];
  assign _0252_ = _0029_ ? keysched_new_key_o[51] : _0251_;
  assign _0253_ = _0016_ ? key_i[51] : _0252_;
  assign keysched_last_key_i[51] = _0004_ ? _0251_ : _0253_;
  assign _0254_ = _0014_ ? key_i[52] : keysched_new_key_o[52];
  assign _0255_ = _0029_ ? keysched_new_key_o[52] : _0254_;
  assign _0256_ = _0016_ ? key_i[52] : _0255_;
  assign keysched_last_key_i[52] = _0004_ ? _0254_ : _0256_;
  assign _0257_ = _0014_ ? key_i[53] : keysched_new_key_o[53];
  assign _0258_ = _0029_ ? keysched_new_key_o[53] : _0257_;
  assign _0259_ = _0016_ ? key_i[53] : _0258_;
  assign keysched_last_key_i[53] = _0004_ ? _0257_ : _0259_;
  assign _0260_ = _0014_ ? key_i[54] : keysched_new_key_o[54];
  assign _0261_ = _0029_ ? keysched_new_key_o[54] : _0260_;
  assign _0262_ = _0016_ ? key_i[54] : _0261_;
  assign keysched_last_key_i[54] = _0004_ ? _0260_ : _0262_;
  assign _0263_ = _0014_ ? key_i[55] : keysched_new_key_o[55];
  assign _0264_ = _0029_ ? keysched_new_key_o[55] : _0263_;
  assign _0265_ = _0016_ ? key_i[55] : _0264_;
  assign keysched_last_key_i[55] = _0004_ ? _0263_ : _0265_;
  assign _0266_ = _0014_ ? key_i[56] : keysched_new_key_o[56];
  assign _0267_ = _0029_ ? keysched_new_key_o[56] : _0266_;
  assign _0268_ = _0016_ ? key_i[56] : _0267_;
  assign keysched_last_key_i[56] = _0004_ ? _0266_ : _0268_;
  assign _0269_ = _0014_ ? key_i[57] : keysched_new_key_o[57];
  assign _0270_ = _0029_ ? keysched_new_key_o[57] : _0269_;
  assign _0271_ = _0016_ ? key_i[57] : _0270_;
  assign keysched_last_key_i[57] = _0004_ ? _0269_ : _0271_;
  assign _0272_ = _0014_ ? key_i[58] : keysched_new_key_o[58];
  assign _0273_ = _0029_ ? keysched_new_key_o[58] : _0272_;
  assign _0274_ = _0016_ ? key_i[58] : _0273_;
  assign keysched_last_key_i[58] = _0004_ ? _0272_ : _0274_;
  assign _0275_ = _0014_ ? key_i[59] : keysched_new_key_o[59];
  assign _0276_ = _0029_ ? keysched_new_key_o[59] : _0275_;
  assign _0277_ = _0016_ ? key_i[59] : _0276_;
  assign keysched_last_key_i[59] = _0004_ ? _0275_ : _0277_;
  assign _0278_ = _0014_ ? key_i[5] : keysched_new_key_o[5];
  assign _0279_ = _0029_ ? keysched_new_key_o[5] : _0278_;
  assign _0280_ = _0016_ ? key_i[5] : _0279_;
  assign keysched_last_key_i[5] = _0004_ ? _0278_ : _0280_;
  assign _0281_ = _0014_ ? key_i[60] : keysched_new_key_o[60];
  assign _0282_ = _0029_ ? keysched_new_key_o[60] : _0281_;
  assign _0283_ = _0016_ ? key_i[60] : _0282_;
  assign keysched_last_key_i[60] = _0004_ ? _0281_ : _0283_;
  assign _0284_ = _0014_ ? key_i[61] : keysched_new_key_o[61];
  assign _0285_ = _0029_ ? keysched_new_key_o[61] : _0284_;
  assign _0286_ = _0016_ ? key_i[61] : _0285_;
  assign keysched_last_key_i[61] = _0004_ ? _0284_ : _0286_;
  assign _0287_ = _0014_ ? key_i[62] : keysched_new_key_o[62];
  assign _0288_ = _0029_ ? keysched_new_key_o[62] : _0287_;
  assign _0289_ = _0016_ ? key_i[62] : _0288_;
  assign keysched_last_key_i[62] = _0004_ ? _0287_ : _0289_;
  assign _0290_ = _0014_ ? key_i[63] : keysched_new_key_o[63];
  assign _0291_ = _0029_ ? keysched_new_key_o[63] : _0290_;
  assign _0292_ = _0016_ ? key_i[63] : _0291_;
  assign keysched_last_key_i[63] = _0004_ ? _0290_ : _0292_;
  assign _0293_ = _0014_ ? key_i[64] : keysched_new_key_o[64];
  assign _0294_ = _0029_ ? keysched_new_key_o[64] : _0293_;
  assign _0295_ = _0016_ ? key_i[64] : _0294_;
  assign keysched_last_key_i[64] = _0004_ ? _0293_ : _0295_;
  assign _0296_ = _0014_ ? key_i[65] : keysched_new_key_o[65];
  assign _0297_ = _0029_ ? keysched_new_key_o[65] : _0296_;
  assign _0298_ = _0016_ ? key_i[65] : _0297_;
  assign keysched_last_key_i[65] = _0004_ ? _0296_ : _0298_;
  assign _0299_ = _0014_ ? key_i[66] : keysched_new_key_o[66];
  assign _0300_ = _0029_ ? keysched_new_key_o[66] : _0299_;
  assign _0301_ = _0016_ ? key_i[66] : _0300_;
  assign keysched_last_key_i[66] = _0004_ ? _0299_ : _0301_;
  assign _0302_ = _0014_ ? key_i[67] : keysched_new_key_o[67];
  assign _0303_ = _0029_ ? keysched_new_key_o[67] : _0302_;
  assign _0304_ = _0016_ ? key_i[67] : _0303_;
  assign keysched_last_key_i[67] = _0004_ ? _0302_ : _0304_;
  assign _0305_ = _0014_ ? key_i[68] : keysched_new_key_o[68];
  assign _0306_ = _0029_ ? keysched_new_key_o[68] : _0305_;
  assign _0307_ = _0016_ ? key_i[68] : _0306_;
  assign keysched_last_key_i[68] = _0004_ ? _0305_ : _0307_;
  assign _0308_ = _0014_ ? key_i[69] : keysched_new_key_o[69];
  assign _0309_ = _0029_ ? keysched_new_key_o[69] : _0308_;
  assign _0310_ = _0016_ ? key_i[69] : _0309_;
  assign keysched_last_key_i[69] = _0004_ ? _0308_ : _0310_;
  assign _0311_ = _0014_ ? key_i[6] : keysched_new_key_o[6];
  assign _0312_ = _0029_ ? keysched_new_key_o[6] : _0311_;
  assign _0313_ = _0016_ ? key_i[6] : _0312_;
  assign keysched_last_key_i[6] = _0004_ ? _0311_ : _0313_;
  assign _0314_ = _0014_ ? key_i[70] : keysched_new_key_o[70];
  assign _0315_ = _0029_ ? keysched_new_key_o[70] : _0314_;
  assign _0316_ = _0016_ ? key_i[70] : _0315_;
  assign keysched_last_key_i[70] = _0004_ ? _0314_ : _0316_;
  assign _0317_ = _0014_ ? key_i[71] : keysched_new_key_o[71];
  assign _0318_ = _0029_ ? keysched_new_key_o[71] : _0317_;
  assign _0319_ = _0016_ ? key_i[71] : _0318_;
  assign keysched_last_key_i[71] = _0004_ ? _0317_ : _0319_;
  assign _0320_ = _0014_ ? key_i[72] : keysched_new_key_o[72];
  assign _0321_ = _0029_ ? keysched_new_key_o[72] : _0320_;
  assign _0322_ = _0016_ ? key_i[72] : _0321_;
  assign keysched_last_key_i[72] = _0004_ ? _0320_ : _0322_;
  assign _0323_ = _0014_ ? key_i[73] : keysched_new_key_o[73];
  assign _0324_ = _0029_ ? keysched_new_key_o[73] : _0323_;
  assign _0325_ = _0016_ ? key_i[73] : _0324_;
  assign keysched_last_key_i[73] = _0004_ ? _0323_ : _0325_;
  assign _0326_ = _0014_ ? key_i[74] : keysched_new_key_o[74];
  assign _0327_ = _0029_ ? keysched_new_key_o[74] : _0326_;
  assign _0328_ = _0016_ ? key_i[74] : _0327_;
  assign keysched_last_key_i[74] = _0004_ ? _0326_ : _0328_;
  assign _0329_ = _0014_ ? key_i[75] : keysched_new_key_o[75];
  assign _0330_ = _0029_ ? keysched_new_key_o[75] : _0329_;
  assign _0331_ = _0016_ ? key_i[75] : _0330_;
  assign keysched_last_key_i[75] = _0004_ ? _0329_ : _0331_;
  assign _0332_ = _0014_ ? key_i[76] : keysched_new_key_o[76];
  assign _0333_ = _0029_ ? keysched_new_key_o[76] : _0332_;
  assign _0334_ = _0016_ ? key_i[76] : _0333_;
  assign keysched_last_key_i[76] = _0004_ ? _0332_ : _0334_;
  assign _0335_ = _0014_ ? key_i[77] : keysched_new_key_o[77];
  assign _0336_ = _0029_ ? keysched_new_key_o[77] : _0335_;
  assign _0337_ = _0016_ ? key_i[77] : _0336_;
  assign keysched_last_key_i[77] = _0004_ ? _0335_ : _0337_;
  assign _0338_ = _0014_ ? key_i[78] : keysched_new_key_o[78];
  assign _0339_ = _0029_ ? keysched_new_key_o[78] : _0338_;
  assign _0340_ = _0016_ ? key_i[78] : _0339_;
  assign keysched_last_key_i[78] = _0004_ ? _0338_ : _0340_;
  assign _0341_ = _0014_ ? key_i[79] : keysched_new_key_o[79];
  assign _0342_ = _0029_ ? keysched_new_key_o[79] : _0341_;
  assign _0343_ = _0016_ ? key_i[79] : _0342_;
  assign keysched_last_key_i[79] = _0004_ ? _0341_ : _0343_;
  assign _0344_ = _0014_ ? key_i[7] : keysched_new_key_o[7];
  assign _0345_ = _0029_ ? keysched_new_key_o[7] : _0344_;
  assign _0346_ = _0016_ ? key_i[7] : _0345_;
  assign keysched_last_key_i[7] = _0004_ ? _0344_ : _0346_;
  assign _0347_ = _0014_ ? key_i[80] : keysched_new_key_o[80];
  assign _0348_ = _0029_ ? keysched_new_key_o[80] : _0347_;
  assign _0349_ = _0016_ ? key_i[80] : _0348_;
  assign keysched_last_key_i[80] = _0004_ ? _0347_ : _0349_;
  assign _0350_ = _0014_ ? key_i[81] : keysched_new_key_o[81];
  assign _0351_ = _0029_ ? keysched_new_key_o[81] : _0350_;
  assign _0352_ = _0016_ ? key_i[81] : _0351_;
  assign keysched_last_key_i[81] = _0004_ ? _0350_ : _0352_;
  assign _0353_ = _0014_ ? key_i[82] : keysched_new_key_o[82];
  assign _0354_ = _0029_ ? keysched_new_key_o[82] : _0353_;
  assign _0355_ = _0016_ ? key_i[82] : _0354_;
  assign keysched_last_key_i[82] = _0004_ ? _0353_ : _0355_;
  assign _0356_ = _0014_ ? key_i[83] : keysched_new_key_o[83];
  assign _0357_ = _0029_ ? keysched_new_key_o[83] : _0356_;
  assign _0358_ = _0016_ ? key_i[83] : _0357_;
  assign keysched_last_key_i[83] = _0004_ ? _0356_ : _0358_;
  assign _0359_ = _0014_ ? key_i[84] : keysched_new_key_o[84];
  assign _0360_ = _0029_ ? keysched_new_key_o[84] : _0359_;
  assign _0361_ = _0016_ ? key_i[84] : _0360_;
  assign keysched_last_key_i[84] = _0004_ ? _0359_ : _0361_;
  assign _0362_ = _0014_ ? key_i[85] : keysched_new_key_o[85];
  assign _0363_ = _0029_ ? keysched_new_key_o[85] : _0362_;
  assign _0364_ = _0016_ ? key_i[85] : _0363_;
  assign keysched_last_key_i[85] = _0004_ ? _0362_ : _0364_;
  assign _0365_ = _0014_ ? key_i[86] : keysched_new_key_o[86];
  assign _0366_ = _0029_ ? keysched_new_key_o[86] : _0365_;
  assign _0367_ = _0016_ ? key_i[86] : _0366_;
  assign keysched_last_key_i[86] = _0004_ ? _0365_ : _0367_;
  assign _0368_ = _0014_ ? key_i[87] : keysched_new_key_o[87];
  assign _0369_ = _0029_ ? keysched_new_key_o[87] : _0368_;
  assign _0370_ = _0016_ ? key_i[87] : _0369_;
  assign keysched_last_key_i[87] = _0004_ ? _0368_ : _0370_;
  assign _0371_ = _0014_ ? key_i[88] : keysched_new_key_o[88];
  assign _0372_ = _0029_ ? keysched_new_key_o[88] : _0371_;
  assign _0373_ = _0016_ ? key_i[88] : _0372_;
  assign keysched_last_key_i[88] = _0004_ ? _0371_ : _0373_;
  assign _0374_ = _0014_ ? key_i[89] : keysched_new_key_o[89];
  assign _0375_ = _0029_ ? keysched_new_key_o[89] : _0374_;
  assign _0376_ = _0016_ ? key_i[89] : _0375_;
  assign keysched_last_key_i[89] = _0004_ ? _0374_ : _0376_;
  assign _0377_ = _0014_ ? key_i[8] : keysched_new_key_o[8];
  assign _0378_ = _0029_ ? keysched_new_key_o[8] : _0377_;
  assign _0379_ = _0016_ ? key_i[8] : _0378_;
  assign keysched_last_key_i[8] = _0004_ ? _0377_ : _0379_;
  assign _0380_ = _0014_ ? key_i[90] : keysched_new_key_o[90];
  assign _0381_ = _0029_ ? keysched_new_key_o[90] : _0380_;
  assign _0382_ = _0016_ ? key_i[90] : _0381_;
  assign keysched_last_key_i[90] = _0004_ ? _0380_ : _0382_;
  assign _0383_ = _0014_ ? key_i[91] : keysched_new_key_o[91];
  assign _0384_ = _0029_ ? keysched_new_key_o[91] : _0383_;
  assign _0385_ = _0016_ ? key_i[91] : _0384_;
  assign keysched_last_key_i[91] = _0004_ ? _0383_ : _0385_;
  assign _0386_ = _0014_ ? key_i[92] : keysched_new_key_o[92];
  assign _0387_ = _0029_ ? keysched_new_key_o[92] : _0386_;
  assign _0388_ = _0016_ ? key_i[92] : _0387_;
  assign keysched_last_key_i[92] = _0004_ ? _0386_ : _0388_;
  assign _0389_ = _0014_ ? key_i[93] : keysched_new_key_o[93];
  assign _0390_ = _0029_ ? keysched_new_key_o[93] : _0389_;
  assign _0391_ = _0016_ ? key_i[93] : _0390_;
  assign keysched_last_key_i[93] = _0004_ ? _0389_ : _0391_;
  assign _0392_ = _0014_ ? key_i[94] : keysched_new_key_o[94];
  assign _0393_ = _0029_ ? keysched_new_key_o[94] : _0392_;
  assign _0394_ = _0016_ ? key_i[94] : _0393_;
  assign keysched_last_key_i[94] = _0004_ ? _0392_ : _0394_;
  assign _0395_ = _0014_ ? key_i[95] : keysched_new_key_o[95];
  assign _0396_ = _0029_ ? keysched_new_key_o[95] : _0395_;
  assign _0397_ = _0016_ ? key_i[95] : _0396_;
  assign keysched_last_key_i[95] = _0004_ ? _0395_ : _0397_;
  assign _0398_ = _0014_ ? key_i[96] : keysched_new_key_o[96];
  assign _0399_ = _0029_ ? keysched_new_key_o[96] : _0398_;
  assign _0400_ = _0016_ ? key_i[96] : _0399_;
  assign keysched_last_key_i[96] = _0004_ ? _0398_ : _0400_;
  assign _0401_ = _0014_ ? key_i[97] : keysched_new_key_o[97];
  assign _0402_ = _0029_ ? keysched_new_key_o[97] : _0401_;
  assign _0403_ = _0016_ ? key_i[97] : _0402_;
  assign keysched_last_key_i[97] = _0004_ ? _0401_ : _0403_;
  assign _0404_ = _0014_ ? key_i[98] : keysched_new_key_o[98];
  assign _0405_ = _0029_ ? keysched_new_key_o[98] : _0404_;
  assign _0406_ = _0016_ ? key_i[98] : _0405_;
  assign keysched_last_key_i[98] = _0004_ ? _0404_ : _0406_;
  assign _0407_ = _0014_ ? key_i[99] : keysched_new_key_o[99];
  assign _0408_ = _0029_ ? keysched_new_key_o[99] : _0407_;
  assign _0409_ = _0016_ ? key_i[99] : _0408_;
  assign keysched_last_key_i[99] = _0004_ ? _0407_ : _0409_;
  assign _0410_ = _0014_ ? key_i[9] : keysched_new_key_o[9];
  assign _0411_ = _0029_ ? keysched_new_key_o[9] : _0410_;
  assign _0412_ = _0016_ ? key_i[9] : _0411_;
  assign keysched_last_key_i[9] = _0004_ ? _0410_ : _0412_;
  assign _0413_ = _0029_ ^ addroundkey_round[0];
  assign _0414_ = _0413_ | _0016_;
  assign keysched_round_i[0] = _0004_ ? addroundkey_round[0] : _0414_;
  assign _0415_ = _0004_ & addroundkey_round[1];
  assign _0416_ = addroundkey_round[1] ^ addroundkey_round[0];
  assign _0417_ = _0029_ ? _0416_ : addroundkey_round[1];
  assign _0418_ = ~_0004_;
  assign _0419_ = ~_0016_;
  assign _0420_ = _0419_ & _0418_;
  assign _0421_ = _0420_ & _0417_;
  assign keysched_round_i[1] = _0421_ | _0415_;
  assign _0422_ = _0004_ & addroundkey_round[2];
  assign _0423_ = addroundkey_round[1] & addroundkey_round[0];
  assign _0424_ = _0423_ ^ addroundkey_round[2];
  assign _0425_ = _0029_ ? _0424_ : addroundkey_round[2];
  assign _0426_ = _0425_ & _0420_;
  assign keysched_round_i[2] = _0426_ | _0422_;
  assign _0427_ = _0004_ & addroundkey_round[3];
  assign _0428_ = _0423_ & addroundkey_round[2];
  assign _0429_ = _0428_ ^ addroundkey_round[3];
  assign _0430_ = _0029_ ? _0429_ : addroundkey_round[3];
  assign _0431_ = _0430_ & _0420_;
  assign keysched_round_i[3] = _0431_ | _0427_;
  assign keysched_start_i = addroundkey_start_i ? _0002_ : _0029_;
  assign _0432_ = _0029_ & _0011_;
  assign _0433_ = ~keysched_ready_o;
  assign _0434_ = _0433_ & addroundkey_round[0];
  assign _0435_ = _0434_ | _0432_;
  assign _0436_ = _0435_ | _0016_;
  assign next_addroundkey_round[0] = _0004_ ? addroundkey_round[0] : _0436_;
  assign _0437_ = _0416_ & _0029_;
  assign _0438_ = _0433_ & addroundkey_round[1];
  assign _0439_ = _0438_ | _0437_;
  assign _0440_ = _0439_ & _0420_;
  assign next_addroundkey_round[1] = _0440_ | _0415_;
  assign _0441_ = _0424_ & _0029_;
  assign _0442_ = _0433_ & addroundkey_round[2];
  assign _0443_ = _0442_ | _0441_;
  assign _0444_ = _0443_ & _0420_;
  assign next_addroundkey_round[2] = _0444_ | _0422_;
  assign _0445_ = _0429_ & _0029_;
  assign _0446_ = _0433_ & addroundkey_round[3];
  assign _0447_ = _0446_ | _0445_;
  assign _0448_ = _0447_ & _0420_;
  assign next_addroundkey_round[3] = _0448_ | _0427_;
  assign _0449_ = ~key_i[0];
  assign _0450_ = ~state;
  assign _0451_ = ~subbytes_data_o[0];
  assign _0452_ = _0017_ | round[0];
  assign _0453_ = _0022_ | round[2];
  assign _0454_ = _0453_ | _0452_;
  assign _0455_ = _0454_ & decrypt_i;
  assign _0456_ = ~mixcol_data_o[0];
  assign _0457_ = ~data_i[0];
  assign _0458_ = ~decrypt_i;
  assign _0459_ = _0002_ & _0458_;
  assign _0460_ = _0459_ ? _0456_ : _0457_;
  assign _0461_ = _0455_ ? _0451_ : _0460_;
  assign _0462_ = decrypt_i ? _0002_ : _0454_;
  assign _0463_ = ~_0462_;
  assign _0464_ = _0002_ | _0458_;
  assign _0465_ = round[1] | _0019_;
  assign _0466_ = _0453_ | decrypt_i;
  assign _0467_ = _0466_ | _0465_;
  assign _0468_ = _0467_ & _0464_;
  assign _0469_ = mixcol_ready_o & _0458_;
  assign _0470_ = subbytes_ready_o & decrypt_i;
  assign _0471_ = _0470_ ? _0451_ : _0461_;
  assign _0472_ = _0469_ ? _0456_ : _0471_;
  assign _0473_ = subbytes_ready_o ? _0451_ : _0472_;
  assign _0474_ = _0468_ ? _0472_ : _0473_;
  assign _0475_ = _0463_ ? _0451_ : _0474_;
  assign _0476_ = _0450_ ? _0461_ : _0475_;
  assign _0477_ = _0476_ ^ _0449_;
  assign _0478_ = _0027_ & keysched_ready_o;
  assign _0479_ = ~_0478_;
  assign _0480_ = ~keysched_new_key_o[0];
  assign _0481_ = _0476_ ^ _0480_;
  assign _0482_ = _0479_ ? addroundkey_data_o[0] : _0481_;
  assign _0483_ = _0016_ ? addroundkey_data_o[0] : _0482_;
  assign next_addroundkey_data_reg[0] = _0004_ ? _0477_ : _0483_;
  assign _0484_ = ~key_i[100];
  assign _0485_ = ~subbytes_data_o[100];
  assign _0486_ = ~mixcol_data_o[100];
  assign _0487_ = ~data_i[100];
  assign _0488_ = _0459_ ? _0486_ : _0487_;
  assign _0489_ = _0455_ ? _0485_ : _0488_;
  assign _0490_ = _0470_ ? _0485_ : _0489_;
  assign _0491_ = _0469_ ? _0486_ : _0490_;
  assign _0492_ = subbytes_ready_o ? _0485_ : _0491_;
  assign _0493_ = _0468_ ? _0491_ : _0492_;
  assign _0494_ = _0463_ ? _0485_ : _0493_;
  assign _0495_ = _0450_ ? _0489_ : _0494_;
  assign _0496_ = _0495_ ^ _0484_;
  assign _0497_ = ~keysched_new_key_o[100];
  assign _0498_ = _0495_ ^ _0497_;
  assign _0499_ = _0479_ ? addroundkey_data_o[100] : _0498_;
  assign _0500_ = _0016_ ? addroundkey_data_o[100] : _0499_;
  assign next_addroundkey_data_reg[100] = _0004_ ? _0496_ : _0500_;
  assign _0501_ = ~key_i[101];
  assign _0502_ = ~subbytes_data_o[101];
  assign _0503_ = ~mixcol_data_o[101];
  assign _0504_ = ~data_i[101];
  assign _0505_ = _0459_ ? _0503_ : _0504_;
  assign _0506_ = _0455_ ? _0502_ : _0505_;
  assign _0507_ = _0470_ ? _0502_ : _0506_;
  assign _0508_ = _0469_ ? _0503_ : _0507_;
  assign _0509_ = subbytes_ready_o ? _0502_ : _0508_;
  assign _0510_ = _0468_ ? _0508_ : _0509_;
  assign _0511_ = _0463_ ? _0502_ : _0510_;
  assign _0512_ = _0450_ ? _0506_ : _0511_;
  assign _0513_ = _0512_ ^ _0501_;
  assign _0514_ = ~keysched_new_key_o[101];
  assign _0515_ = _0512_ ^ _0514_;
  assign _0516_ = _0479_ ? addroundkey_data_o[101] : _0515_;
  assign _0517_ = _0016_ ? addroundkey_data_o[101] : _0516_;
  assign next_addroundkey_data_reg[101] = _0004_ ? _0513_ : _0517_;
  assign _0518_ = ~key_i[102];
  assign _0519_ = ~subbytes_data_o[102];
  assign _0520_ = ~mixcol_data_o[102];
  assign _0521_ = ~data_i[102];
  assign _0522_ = _0459_ ? _0520_ : _0521_;
  assign _0523_ = _0455_ ? _0519_ : _0522_;
  assign _0524_ = _0470_ ? _0519_ : _0523_;
  assign _0525_ = _0469_ ? _0520_ : _0524_;
  assign _0526_ = subbytes_ready_o ? _0519_ : _0525_;
  assign _0527_ = _0468_ ? _0525_ : _0526_;
  assign _0528_ = _0463_ ? _0519_ : _0527_;
  assign _0529_ = _0450_ ? _0523_ : _0528_;
  assign _0530_ = _0529_ ^ _0518_;
  assign _0531_ = ~keysched_new_key_o[102];
  assign _0532_ = _0529_ ^ _0531_;
  assign _0533_ = _0479_ ? addroundkey_data_o[102] : _0532_;
  assign _0534_ = _0016_ ? addroundkey_data_o[102] : _0533_;
  assign next_addroundkey_data_reg[102] = _0004_ ? _0530_ : _0534_;
  assign _0535_ = ~key_i[103];
  assign _0536_ = ~subbytes_data_o[103];
  assign _0537_ = ~mixcol_data_o[103];
  assign _0538_ = ~data_i[103];
  assign _0539_ = _0459_ ? _0537_ : _0538_;
  assign _0540_ = _0455_ ? _0536_ : _0539_;
  assign _0541_ = _0470_ ? _0536_ : _0540_;
  assign _0542_ = _0469_ ? _0537_ : _0541_;
  assign _0543_ = subbytes_ready_o ? _0536_ : _0542_;
  assign _0544_ = _0468_ ? _0542_ : _0543_;
  assign _0545_ = _0463_ ? _0536_ : _0544_;
  assign _0546_ = _0450_ ? _0540_ : _0545_;
  assign _0547_ = _0546_ ^ _0535_;
  assign _0548_ = ~keysched_new_key_o[103];
  assign _0549_ = _0546_ ^ _0548_;
  assign _0550_ = _0479_ ? addroundkey_data_o[103] : _0549_;
  assign _0551_ = _0016_ ? addroundkey_data_o[103] : _0550_;
  assign next_addroundkey_data_reg[103] = _0004_ ? _0547_ : _0551_;
  assign _0552_ = ~key_i[104];
  assign _0553_ = ~subbytes_data_o[104];
  assign _0554_ = ~mixcol_data_o[104];
  assign _0555_ = ~data_i[104];
  assign _0556_ = _0459_ ? _0554_ : _0555_;
  assign _0557_ = _0455_ ? _0553_ : _0556_;
  assign _0558_ = _0470_ ? _0553_ : _0557_;
  assign _0559_ = _0469_ ? _0554_ : _0558_;
  assign _0560_ = subbytes_ready_o ? _0553_ : _0559_;
  assign _0561_ = _0468_ ? _0559_ : _0560_;
  assign _0562_ = _0463_ ? _0553_ : _0561_;
  assign _0563_ = _0450_ ? _0557_ : _0562_;
  assign _0564_ = _0563_ ^ _0552_;
  assign _0565_ = ~keysched_new_key_o[104];
  assign _0566_ = _0563_ ^ _0565_;
  assign _0567_ = _0479_ ? addroundkey_data_o[104] : _0566_;
  assign _0568_ = _0016_ ? addroundkey_data_o[104] : _0567_;
  assign next_addroundkey_data_reg[104] = _0004_ ? _0564_ : _0568_;
  assign _0569_ = ~key_i[105];
  assign _0570_ = ~subbytes_data_o[105];
  assign _0571_ = ~mixcol_data_o[105];
  assign _0572_ = ~data_i[105];
  assign _0573_ = _0459_ ? _0571_ : _0572_;
  assign _0574_ = _0455_ ? _0570_ : _0573_;
  assign _0575_ = _0470_ ? _0570_ : _0574_;
  assign _0576_ = _0469_ ? _0571_ : _0575_;
  assign _0577_ = subbytes_ready_o ? _0570_ : _0576_;
  assign _0578_ = _0468_ ? _0576_ : _0577_;
  assign _0579_ = _0463_ ? _0570_ : _0578_;
  assign _0580_ = _0450_ ? _0574_ : _0579_;
  assign _0581_ = _0580_ ^ _0569_;
  assign _0582_ = ~keysched_new_key_o[105];
  assign _0583_ = _0580_ ^ _0582_;
  assign _0584_ = _0479_ ? addroundkey_data_o[105] : _0583_;
  assign _0585_ = _0016_ ? addroundkey_data_o[105] : _0584_;
  assign next_addroundkey_data_reg[105] = _0004_ ? _0581_ : _0585_;
  assign _0586_ = ~key_i[106];
  assign _0587_ = ~subbytes_data_o[106];
  assign _0588_ = ~mixcol_data_o[106];
  assign _0589_ = ~data_i[106];
  assign _0590_ = _0459_ ? _0588_ : _0589_;
  assign _0591_ = _0455_ ? _0587_ : _0590_;
  assign _0592_ = _0470_ ? _0587_ : _0591_;
  assign _0593_ = _0469_ ? _0588_ : _0592_;
  assign _0594_ = subbytes_ready_o ? _0587_ : _0593_;
  assign _0595_ = _0468_ ? _0593_ : _0594_;
  assign _0596_ = _0463_ ? _0587_ : _0595_;
  assign _0597_ = _0450_ ? _0591_ : _0596_;
  assign _0598_ = _0597_ ^ _0586_;
  assign _0599_ = ~keysched_new_key_o[106];
  assign _0600_ = _0597_ ^ _0599_;
  assign _0601_ = _0479_ ? addroundkey_data_o[106] : _0600_;
  assign _0602_ = _0016_ ? addroundkey_data_o[106] : _0601_;
  assign next_addroundkey_data_reg[106] = _0004_ ? _0598_ : _0602_;
  assign _0603_ = ~key_i[107];
  assign _0604_ = ~subbytes_data_o[107];
  assign _0605_ = ~mixcol_data_o[107];
  assign _0606_ = ~data_i[107];
  assign _0607_ = _0459_ ? _0605_ : _0606_;
  assign _0608_ = _0455_ ? _0604_ : _0607_;
  assign _0609_ = _0470_ ? _0604_ : _0608_;
  assign _0610_ = _0469_ ? _0605_ : _0609_;
  assign _0611_ = subbytes_ready_o ? _0604_ : _0610_;
  assign _0612_ = _0468_ ? _0610_ : _0611_;
  assign _0613_ = _0463_ ? _0604_ : _0612_;
  assign _0614_ = _0450_ ? _0608_ : _0613_;
  assign _0615_ = _0614_ ^ _0603_;
  assign _0616_ = ~keysched_new_key_o[107];
  assign _0617_ = _0614_ ^ _0616_;
  assign _0618_ = _0479_ ? addroundkey_data_o[107] : _0617_;
  assign _0619_ = _0016_ ? addroundkey_data_o[107] : _0618_;
  assign next_addroundkey_data_reg[107] = _0004_ ? _0615_ : _0619_;
  assign _0620_ = ~key_i[108];
  assign _0621_ = ~subbytes_data_o[108];
  assign _0622_ = ~mixcol_data_o[108];
  assign _0623_ = ~data_i[108];
  assign _0624_ = _0459_ ? _0622_ : _0623_;
  assign _0625_ = _0455_ ? _0621_ : _0624_;
  assign _0626_ = _0470_ ? _0621_ : _0625_;
  assign _0627_ = _0469_ ? _0622_ : _0626_;
  assign _0628_ = subbytes_ready_o ? _0621_ : _0627_;
  assign _0629_ = _0468_ ? _0627_ : _0628_;
  assign _0630_ = _0463_ ? _0621_ : _0629_;
  assign _0631_ = _0450_ ? _0625_ : _0630_;
  assign _0632_ = _0631_ ^ _0620_;
  assign _0633_ = ~keysched_new_key_o[108];
  assign _0634_ = _0631_ ^ _0633_;
  assign _0635_ = _0479_ ? addroundkey_data_o[108] : _0634_;
  assign _0636_ = _0016_ ? addroundkey_data_o[108] : _0635_;
  assign next_addroundkey_data_reg[108] = _0004_ ? _0632_ : _0636_;
  assign _0637_ = ~key_i[109];
  assign _0638_ = ~subbytes_data_o[109];
  assign _0639_ = ~mixcol_data_o[109];
  assign _0640_ = ~data_i[109];
  assign _0641_ = _0459_ ? _0639_ : _0640_;
  assign _0642_ = _0455_ ? _0638_ : _0641_;
  assign _0643_ = _0470_ ? _0638_ : _0642_;
  assign _0644_ = _0469_ ? _0639_ : _0643_;
  assign _0645_ = subbytes_ready_o ? _0638_ : _0644_;
  assign _0646_ = _0468_ ? _0644_ : _0645_;
  assign _0647_ = _0463_ ? _0638_ : _0646_;
  assign _0648_ = _0450_ ? _0642_ : _0647_;
  assign _0649_ = _0648_ ^ _0637_;
  assign _0650_ = ~keysched_new_key_o[109];
  assign _0651_ = _0648_ ^ _0650_;
  assign _0652_ = _0479_ ? addroundkey_data_o[109] : _0651_;
  assign _0653_ = _0016_ ? addroundkey_data_o[109] : _0652_;
  assign next_addroundkey_data_reg[109] = _0004_ ? _0649_ : _0653_;
  assign _0654_ = ~key_i[10];
  assign _0655_ = ~subbytes_data_o[10];
  assign _0656_ = ~mixcol_data_o[10];
  assign _0657_ = ~data_i[10];
  assign _0658_ = _0459_ ? _0656_ : _0657_;
  assign _0659_ = _0455_ ? _0655_ : _0658_;
  assign _0660_ = _0470_ ? _0655_ : _0659_;
  assign _0661_ = _0469_ ? _0656_ : _0660_;
  assign _0662_ = subbytes_ready_o ? _0655_ : _0661_;
  assign _0663_ = _0468_ ? _0661_ : _0662_;
  assign _0664_ = _0463_ ? _0655_ : _0663_;
  assign _0665_ = _0450_ ? _0659_ : _0664_;
  assign _0666_ = _0665_ ^ _0654_;
  assign _0667_ = ~keysched_new_key_o[10];
  assign _0668_ = _0665_ ^ _0667_;
  assign _0669_ = _0479_ ? addroundkey_data_o[10] : _0668_;
  assign _0670_ = _0016_ ? addroundkey_data_o[10] : _0669_;
  assign next_addroundkey_data_reg[10] = _0004_ ? _0666_ : _0670_;
  assign _0671_ = ~key_i[110];
  assign _0672_ = ~subbytes_data_o[110];
  assign _0673_ = ~mixcol_data_o[110];
  assign _0674_ = ~data_i[110];
  assign _0675_ = _0459_ ? _0673_ : _0674_;
  assign _0676_ = _0455_ ? _0672_ : _0675_;
  assign _0677_ = _0470_ ? _0672_ : _0676_;
  assign _0678_ = _0469_ ? _0673_ : _0677_;
  assign _0679_ = subbytes_ready_o ? _0672_ : _0678_;
  assign _0680_ = _0468_ ? _0678_ : _0679_;
  assign _0681_ = _0463_ ? _0672_ : _0680_;
  assign _0682_ = _0450_ ? _0676_ : _0681_;
  assign _0683_ = _0682_ ^ _0671_;
  assign _0684_ = ~keysched_new_key_o[110];
  assign _0685_ = _0682_ ^ _0684_;
  assign _0686_ = _0479_ ? addroundkey_data_o[110] : _0685_;
  assign _0687_ = _0016_ ? addroundkey_data_o[110] : _0686_;
  assign next_addroundkey_data_reg[110] = _0004_ ? _0683_ : _0687_;
  assign _0688_ = ~key_i[111];
  assign _0689_ = ~subbytes_data_o[111];
  assign _0690_ = ~mixcol_data_o[111];
  assign _0691_ = ~data_i[111];
  assign _0692_ = _0459_ ? _0690_ : _0691_;
  assign _0693_ = _0455_ ? _0689_ : _0692_;
  assign _0694_ = _0470_ ? _0689_ : _0693_;
  assign _0695_ = _0469_ ? _0690_ : _0694_;
  assign _0696_ = subbytes_ready_o ? _0689_ : _0695_;
  assign _0697_ = _0468_ ? _0695_ : _0696_;
  assign _0698_ = _0463_ ? _0689_ : _0697_;
  assign _0699_ = _0450_ ? _0693_ : _0698_;
  assign _0700_ = _0699_ ^ _0688_;
  assign _0701_ = ~keysched_new_key_o[111];
  assign _0702_ = _0699_ ^ _0701_;
  assign _0703_ = _0479_ ? addroundkey_data_o[111] : _0702_;
  assign _0704_ = _0016_ ? addroundkey_data_o[111] : _0703_;
  assign next_addroundkey_data_reg[111] = _0004_ ? _0700_ : _0704_;
  assign _0705_ = ~key_i[112];
  assign _0706_ = ~subbytes_data_o[112];
  assign _0707_ = ~mixcol_data_o[112];
  assign _0708_ = ~data_i[112];
  assign _0709_ = _0459_ ? _0707_ : _0708_;
  assign _0710_ = _0455_ ? _0706_ : _0709_;
  assign _0711_ = _0470_ ? _0706_ : _0710_;
  assign _0712_ = _0469_ ? _0707_ : _0711_;
  assign _0713_ = subbytes_ready_o ? _0706_ : _0712_;
  assign _0714_ = _0468_ ? _0712_ : _0713_;
  assign _0715_ = _0463_ ? _0706_ : _0714_;
  assign _0716_ = _0450_ ? _0710_ : _0715_;
  assign _0717_ = _0716_ ^ _0705_;
  assign _0718_ = ~keysched_new_key_o[112];
  assign _0719_ = _0716_ ^ _0718_;
  assign _0720_ = _0479_ ? addroundkey_data_o[112] : _0719_;
  assign _0721_ = _0016_ ? addroundkey_data_o[112] : _0720_;
  assign next_addroundkey_data_reg[112] = _0004_ ? _0717_ : _0721_;
  assign _0722_ = ~key_i[113];
  assign _0723_ = ~subbytes_data_o[113];
  assign _0724_ = ~mixcol_data_o[113];
  assign _0725_ = ~data_i[113];
  assign _0726_ = _0459_ ? _0724_ : _0725_;
  assign _0727_ = _0455_ ? _0723_ : _0726_;
  assign _0728_ = _0470_ ? _0723_ : _0727_;
  assign _0729_ = _0469_ ? _0724_ : _0728_;
  assign _0730_ = subbytes_ready_o ? _0723_ : _0729_;
  assign _0731_ = _0468_ ? _0729_ : _0730_;
  assign _0732_ = _0463_ ? _0723_ : _0731_;
  assign _0733_ = _0450_ ? _0727_ : _0732_;
  assign _0734_ = _0733_ ^ _0722_;
  assign _0735_ = ~keysched_new_key_o[113];
  assign _0736_ = _0733_ ^ _0735_;
  assign _0737_ = _0479_ ? addroundkey_data_o[113] : _0736_;
  assign _0738_ = _0016_ ? addroundkey_data_o[113] : _0737_;
  assign next_addroundkey_data_reg[113] = _0004_ ? _0734_ : _0738_;
  assign _0739_ = ~key_i[114];
  assign _0740_ = ~subbytes_data_o[114];
  assign _0741_ = ~mixcol_data_o[114];
  assign _0742_ = ~data_i[114];
  assign _0743_ = _0459_ ? _0741_ : _0742_;
  assign _0744_ = _0455_ ? _0740_ : _0743_;
  assign _0745_ = _0470_ ? _0740_ : _0744_;
  assign _0746_ = _0469_ ? _0741_ : _0745_;
  assign _0747_ = subbytes_ready_o ? _0740_ : _0746_;
  assign _0748_ = _0468_ ? _0746_ : _0747_;
  assign _0749_ = _0463_ ? _0740_ : _0748_;
  assign _0750_ = _0450_ ? _0744_ : _0749_;
  assign _0751_ = _0750_ ^ _0739_;
  assign _0752_ = ~keysched_new_key_o[114];
  assign _0753_ = _0750_ ^ _0752_;
  assign _0754_ = _0479_ ? addroundkey_data_o[114] : _0753_;
  assign _0755_ = _0016_ ? addroundkey_data_o[114] : _0754_;
  assign next_addroundkey_data_reg[114] = _0004_ ? _0751_ : _0755_;
  assign _0756_ = ~key_i[115];
  assign _0757_ = ~subbytes_data_o[115];
  assign _0758_ = ~mixcol_data_o[115];
  assign _0759_ = ~data_i[115];
  assign _0760_ = _0459_ ? _0758_ : _0759_;
  assign _0761_ = _0455_ ? _0757_ : _0760_;
  assign _0762_ = _0470_ ? _0757_ : _0761_;
  assign _0763_ = _0469_ ? _0758_ : _0762_;
  assign _0764_ = subbytes_ready_o ? _0757_ : _0763_;
  assign _0765_ = _0468_ ? _0763_ : _0764_;
  assign _0766_ = _0463_ ? _0757_ : _0765_;
  assign _0767_ = _0450_ ? _0761_ : _0766_;
  assign _0768_ = _0767_ ^ _0756_;
  assign _0769_ = ~keysched_new_key_o[115];
  assign _0770_ = _0767_ ^ _0769_;
  assign _0771_ = _0479_ ? addroundkey_data_o[115] : _0770_;
  assign _0772_ = _0016_ ? addroundkey_data_o[115] : _0771_;
  assign next_addroundkey_data_reg[115] = _0004_ ? _0768_ : _0772_;
  assign _0773_ = ~key_i[116];
  assign _0774_ = ~subbytes_data_o[116];
  assign _0775_ = ~mixcol_data_o[116];
  assign _0776_ = ~data_i[116];
  assign _0777_ = _0459_ ? _0775_ : _0776_;
  assign _0778_ = _0455_ ? _0774_ : _0777_;
  assign _0779_ = _0470_ ? _0774_ : _0778_;
  assign _0780_ = _0469_ ? _0775_ : _0779_;
  assign _0781_ = subbytes_ready_o ? _0774_ : _0780_;
  assign _0782_ = _0468_ ? _0780_ : _0781_;
  assign _0783_ = _0463_ ? _0774_ : _0782_;
  assign _0784_ = _0450_ ? _0778_ : _0783_;
  assign _0785_ = _0784_ ^ _0773_;
  assign _0786_ = ~keysched_new_key_o[116];
  assign _0787_ = _0784_ ^ _0786_;
  assign _0788_ = _0479_ ? addroundkey_data_o[116] : _0787_;
  assign _0789_ = _0016_ ? addroundkey_data_o[116] : _0788_;
  assign next_addroundkey_data_reg[116] = _0004_ ? _0785_ : _0789_;
  assign _0790_ = ~key_i[117];
  assign _0791_ = ~subbytes_data_o[117];
  assign _0792_ = ~mixcol_data_o[117];
  assign _0793_ = ~data_i[117];
  assign _0794_ = _0459_ ? _0792_ : _0793_;
  assign _0795_ = _0455_ ? _0791_ : _0794_;
  assign _0796_ = _0470_ ? _0791_ : _0795_;
  assign _0797_ = _0469_ ? _0792_ : _0796_;
  assign _0798_ = subbytes_ready_o ? _0791_ : _0797_;
  assign _0799_ = _0468_ ? _0797_ : _0798_;
  assign _0800_ = _0463_ ? _0791_ : _0799_;
  assign _0801_ = _0450_ ? _0795_ : _0800_;
  assign _0802_ = _0801_ ^ _0790_;
  assign _0803_ = ~keysched_new_key_o[117];
  assign _0804_ = _0801_ ^ _0803_;
  assign _0805_ = _0479_ ? addroundkey_data_o[117] : _0804_;
  assign _0806_ = _0016_ ? addroundkey_data_o[117] : _0805_;
  assign next_addroundkey_data_reg[117] = _0004_ ? _0802_ : _0806_;
  assign _0807_ = ~key_i[118];
  assign _0808_ = ~subbytes_data_o[118];
  assign _0809_ = ~mixcol_data_o[118];
  assign _0810_ = ~data_i[118];
  assign _0811_ = _0459_ ? _0809_ : _0810_;
  assign _0812_ = _0455_ ? _0808_ : _0811_;
  assign _0813_ = _0470_ ? _0808_ : _0812_;
  assign _0814_ = _0469_ ? _0809_ : _0813_;
  assign _0815_ = subbytes_ready_o ? _0808_ : _0814_;
  assign _0816_ = _0468_ ? _0814_ : _0815_;
  assign _0817_ = _0463_ ? _0808_ : _0816_;
  assign _0818_ = _0450_ ? _0812_ : _0817_;
  assign _0819_ = _0818_ ^ _0807_;
  assign _0820_ = ~keysched_new_key_o[118];
  assign _0821_ = _0818_ ^ _0820_;
  assign _0822_ = _0479_ ? addroundkey_data_o[118] : _0821_;
  assign _0823_ = _0016_ ? addroundkey_data_o[118] : _0822_;
  assign next_addroundkey_data_reg[118] = _0004_ ? _0819_ : _0823_;
  assign _0824_ = ~key_i[119];
  assign _0825_ = ~subbytes_data_o[119];
  assign _0826_ = ~mixcol_data_o[119];
  assign _0827_ = ~data_i[119];
  assign _0828_ = _0459_ ? _0826_ : _0827_;
  assign _0829_ = _0455_ ? _0825_ : _0828_;
  assign _0830_ = _0470_ ? _0825_ : _0829_;
  assign _0831_ = _0469_ ? _0826_ : _0830_;
  assign _0832_ = subbytes_ready_o ? _0825_ : _0831_;
  assign _0833_ = _0468_ ? _0831_ : _0832_;
  assign _0834_ = _0463_ ? _0825_ : _0833_;
  assign _0835_ = _0450_ ? _0829_ : _0834_;
  assign _0836_ = _0835_ ^ _0824_;
  assign _0837_ = ~keysched_new_key_o[119];
  assign _0838_ = _0835_ ^ _0837_;
  assign _0839_ = _0479_ ? addroundkey_data_o[119] : _0838_;
  assign _0840_ = _0016_ ? addroundkey_data_o[119] : _0839_;
  assign next_addroundkey_data_reg[119] = _0004_ ? _0836_ : _0840_;
  assign _0841_ = ~key_i[11];
  assign _0842_ = ~subbytes_data_o[11];
  assign _0843_ = ~mixcol_data_o[11];
  assign _0844_ = ~data_i[11];
  assign _0845_ = _0459_ ? _0843_ : _0844_;
  assign _0846_ = _0455_ ? _0842_ : _0845_;
  assign _0847_ = _0470_ ? _0842_ : _0846_;
  assign _0848_ = _0469_ ? _0843_ : _0847_;
  assign _0849_ = subbytes_ready_o ? _0842_ : _0848_;
  assign _0850_ = _0468_ ? _0848_ : _0849_;
  assign _0851_ = _0463_ ? _0842_ : _0850_;
  assign _0852_ = _0450_ ? _0846_ : _0851_;
  assign _0853_ = _0852_ ^ _0841_;
  assign _0854_ = ~keysched_new_key_o[11];
  assign _0855_ = _0852_ ^ _0854_;
  assign _0856_ = _0479_ ? addroundkey_data_o[11] : _0855_;
  assign _0857_ = _0016_ ? addroundkey_data_o[11] : _0856_;
  assign next_addroundkey_data_reg[11] = _0004_ ? _0853_ : _0857_;
  assign _0858_ = ~key_i[120];
  assign _0859_ = ~subbytes_data_o[120];
  assign _0860_ = ~mixcol_data_o[120];
  assign _0861_ = ~data_i[120];
  assign _0862_ = _0459_ ? _0860_ : _0861_;
  assign _0863_ = _0455_ ? _0859_ : _0862_;
  assign _0864_ = _0470_ ? _0859_ : _0863_;
  assign _0865_ = _0469_ ? _0860_ : _0864_;
  assign _0866_ = subbytes_ready_o ? _0859_ : _0865_;
  assign _0867_ = _0468_ ? _0865_ : _0866_;
  assign _0868_ = _0463_ ? _0859_ : _0867_;
  assign _0869_ = _0450_ ? _0863_ : _0868_;
  assign _0870_ = _0869_ ^ _0858_;
  assign _0871_ = ~keysched_new_key_o[120];
  assign _0872_ = _0869_ ^ _0871_;
  assign _0873_ = _0479_ ? addroundkey_data_o[120] : _0872_;
  assign _0874_ = _0016_ ? addroundkey_data_o[120] : _0873_;
  assign next_addroundkey_data_reg[120] = _0004_ ? _0870_ : _0874_;
  assign _0875_ = ~key_i[121];
  assign _0876_ = ~subbytes_data_o[121];
  assign _0877_ = ~mixcol_data_o[121];
  assign _0878_ = ~data_i[121];
  assign _0879_ = _0459_ ? _0877_ : _0878_;
  assign _0880_ = _0455_ ? _0876_ : _0879_;
  assign _0881_ = _0470_ ? _0876_ : _0880_;
  assign _0882_ = _0469_ ? _0877_ : _0881_;
  assign _0883_ = subbytes_ready_o ? _0876_ : _0882_;
  assign _0884_ = _0468_ ? _0882_ : _0883_;
  assign _0885_ = _0463_ ? _0876_ : _0884_;
  assign _0886_ = _0450_ ? _0880_ : _0885_;
  assign _0887_ = _0886_ ^ _0875_;
  assign _0888_ = ~keysched_new_key_o[121];
  assign _0889_ = _0886_ ^ _0888_;
  assign _0890_ = _0479_ ? addroundkey_data_o[121] : _0889_;
  assign _0891_ = _0016_ ? addroundkey_data_o[121] : _0890_;
  assign next_addroundkey_data_reg[121] = _0004_ ? _0887_ : _0891_;
  assign _0892_ = ~key_i[122];
  assign _0893_ = ~subbytes_data_o[122];
  assign _0894_ = ~mixcol_data_o[122];
  assign _0895_ = ~data_i[122];
  assign _0896_ = _0459_ ? _0894_ : _0895_;
  assign _0897_ = _0455_ ? _0893_ : _0896_;
  assign _0898_ = _0470_ ? _0893_ : _0897_;
  assign _0899_ = _0469_ ? _0894_ : _0898_;
  assign _0900_ = subbytes_ready_o ? _0893_ : _0899_;
  assign _0901_ = _0468_ ? _0899_ : _0900_;
  assign _0902_ = _0463_ ? _0893_ : _0901_;
  assign _0903_ = _0450_ ? _0897_ : _0902_;
  assign _0904_ = _0903_ ^ _0892_;
  assign _0905_ = ~keysched_new_key_o[122];
  assign _0906_ = _0903_ ^ _0905_;
  assign _0907_ = _0479_ ? addroundkey_data_o[122] : _0906_;
  assign _0908_ = _0016_ ? addroundkey_data_o[122] : _0907_;
  assign next_addroundkey_data_reg[122] = _0004_ ? _0904_ : _0908_;
  assign _0909_ = ~key_i[123];
  assign _0910_ = ~subbytes_data_o[123];
  assign _0911_ = ~mixcol_data_o[123];
  assign _0912_ = ~data_i[123];
  assign _0913_ = _0459_ ? _0911_ : _0912_;
  assign _0914_ = _0455_ ? _0910_ : _0913_;
  assign _0915_ = _0470_ ? _0910_ : _0914_;
  assign _0916_ = _0469_ ? _0911_ : _0915_;
  assign _0917_ = subbytes_ready_o ? _0910_ : _0916_;
  assign _0918_ = _0468_ ? _0916_ : _0917_;
  assign _0919_ = _0463_ ? _0910_ : _0918_;
  assign _0920_ = _0450_ ? _0914_ : _0919_;
  assign _0921_ = _0920_ ^ _0909_;
  assign _0922_ = ~keysched_new_key_o[123];
  assign _0923_ = _0920_ ^ _0922_;
  assign _0924_ = _0479_ ? addroundkey_data_o[123] : _0923_;
  assign _0925_ = _0016_ ? addroundkey_data_o[123] : _0924_;
  assign next_addroundkey_data_reg[123] = _0004_ ? _0921_ : _0925_;
  assign _0926_ = ~key_i[124];
  assign _0927_ = ~subbytes_data_o[124];
  assign _0928_ = ~mixcol_data_o[124];
  assign _0929_ = ~data_i[124];
  assign _0930_ = _0459_ ? _0928_ : _0929_;
  assign _0931_ = _0455_ ? _0927_ : _0930_;
  assign _0932_ = _0470_ ? _0927_ : _0931_;
  assign _0933_ = _0469_ ? _0928_ : _0932_;
  assign _0934_ = subbytes_ready_o ? _0927_ : _0933_;
  assign _0935_ = _0468_ ? _0933_ : _0934_;
  assign _0936_ = _0463_ ? _0927_ : _0935_;
  assign _0937_ = _0450_ ? _0931_ : _0936_;
  assign _0938_ = _0937_ ^ _0926_;
  assign _0939_ = ~keysched_new_key_o[124];
  assign _0940_ = _0937_ ^ _0939_;
  assign _0941_ = _0479_ ? addroundkey_data_o[124] : _0940_;
  assign _0942_ = _0016_ ? addroundkey_data_o[124] : _0941_;
  assign next_addroundkey_data_reg[124] = _0004_ ? _0938_ : _0942_;
  assign _0943_ = ~key_i[125];
  assign _0944_ = ~subbytes_data_o[125];
  assign _0945_ = ~mixcol_data_o[125];
  assign _0946_ = ~data_i[125];
  assign _0947_ = _0459_ ? _0945_ : _0946_;
  assign _0948_ = _0455_ ? _0944_ : _0947_;
  assign _0949_ = _0470_ ? _0944_ : _0948_;
  assign _0950_ = _0469_ ? _0945_ : _0949_;
  assign _0951_ = subbytes_ready_o ? _0944_ : _0950_;
  assign _0952_ = _0468_ ? _0950_ : _0951_;
  assign _0953_ = _0463_ ? _0944_ : _0952_;
  assign _0954_ = _0450_ ? _0948_ : _0953_;
  assign _0955_ = _0954_ ^ _0943_;
  assign _0956_ = ~keysched_new_key_o[125];
  assign _0957_ = _0954_ ^ _0956_;
  assign _0958_ = _0479_ ? addroundkey_data_o[125] : _0957_;
  assign _0959_ = _0016_ ? addroundkey_data_o[125] : _0958_;
  assign next_addroundkey_data_reg[125] = _0004_ ? _0955_ : _0959_;
  assign _0960_ = ~key_i[126];
  assign _0961_ = ~subbytes_data_o[126];
  assign _0962_ = ~mixcol_data_o[126];
  assign _0963_ = ~data_i[126];
  assign _0964_ = _0459_ ? _0962_ : _0963_;
  assign _0965_ = _0455_ ? _0961_ : _0964_;
  assign _0966_ = _0470_ ? _0961_ : _0965_;
  assign _0967_ = _0469_ ? _0962_ : _0966_;
  assign _0968_ = subbytes_ready_o ? _0961_ : _0967_;
  assign _0969_ = _0468_ ? _0967_ : _0968_;
  assign _0970_ = _0463_ ? _0961_ : _0969_;
  assign _0971_ = _0450_ ? _0965_ : _0970_;
  assign _0972_ = _0971_ ^ _0960_;
  assign _0973_ = ~keysched_new_key_o[126];
  assign _0974_ = _0971_ ^ _0973_;
  assign _0975_ = _0479_ ? addroundkey_data_o[126] : _0974_;
  assign _0976_ = _0016_ ? addroundkey_data_o[126] : _0975_;
  assign next_addroundkey_data_reg[126] = _0004_ ? _0972_ : _0976_;
  assign _0977_ = ~key_i[127];
  assign _0978_ = ~subbytes_data_o[127];
  assign _0979_ = ~mixcol_data_o[127];
  assign _0980_ = ~data_i[127];
  assign _0981_ = _0459_ ? _0979_ : _0980_;
  assign _0982_ = _0455_ ? _0978_ : _0981_;
  assign _0983_ = _0470_ ? _0978_ : _0982_;
  assign _0984_ = _0469_ ? _0979_ : _0983_;
  assign _0985_ = subbytes_ready_o ? _0978_ : _0984_;
  assign _0986_ = _0468_ ? _0984_ : _0985_;
  assign _0987_ = _0463_ ? _0978_ : _0986_;
  assign _0988_ = _0450_ ? _0982_ : _0987_;
  assign _0989_ = _0988_ ^ _0977_;
  assign _0990_ = ~keysched_new_key_o[127];
  assign _0991_ = _0988_ ^ _0990_;
  assign _0992_ = _0479_ ? addroundkey_data_o[127] : _0991_;
  assign _0993_ = _0016_ ? addroundkey_data_o[127] : _0992_;
  assign next_addroundkey_data_reg[127] = _0004_ ? _0989_ : _0993_;
  assign _0994_ = ~key_i[12];
  assign _0995_ = ~subbytes_data_o[12];
  assign _0996_ = ~mixcol_data_o[12];
  assign _0997_ = ~data_i[12];
  assign _0998_ = _0459_ ? _0996_ : _0997_;
  assign _0999_ = _0455_ ? _0995_ : _0998_;
  assign _1000_ = _0470_ ? _0995_ : _0999_;
  assign _1001_ = _0469_ ? _0996_ : _1000_;
  assign _1002_ = subbytes_ready_o ? _0995_ : _1001_;
  assign _1003_ = _0468_ ? _1001_ : _1002_;
  assign _1004_ = _0463_ ? _0995_ : _1003_;
  assign _1005_ = _0450_ ? _0999_ : _1004_;
  assign _1006_ = _1005_ ^ _0994_;
  assign _1007_ = ~keysched_new_key_o[12];
  assign _1008_ = _1005_ ^ _1007_;
  assign _1009_ = _0479_ ? addroundkey_data_o[12] : _1008_;
  assign _1010_ = _0016_ ? addroundkey_data_o[12] : _1009_;
  assign next_addroundkey_data_reg[12] = _0004_ ? _1006_ : _1010_;
  assign _1011_ = ~key_i[13];
  assign _1012_ = ~subbytes_data_o[13];
  assign _1013_ = ~mixcol_data_o[13];
  assign _1014_ = ~data_i[13];
  assign _1015_ = _0459_ ? _1013_ : _1014_;
  assign _1016_ = _0455_ ? _1012_ : _1015_;
  assign _1017_ = _0470_ ? _1012_ : _1016_;
  assign _1018_ = _0469_ ? _1013_ : _1017_;
  assign _1019_ = subbytes_ready_o ? _1012_ : _1018_;
  assign _1020_ = _0468_ ? _1018_ : _1019_;
  assign _1021_ = _0463_ ? _1012_ : _1020_;
  assign _1022_ = _0450_ ? _1016_ : _1021_;
  assign _1023_ = _1022_ ^ _1011_;
  assign _1024_ = ~keysched_new_key_o[13];
  assign _1025_ = _1022_ ^ _1024_;
  assign _1026_ = _0479_ ? addroundkey_data_o[13] : _1025_;
  assign _1027_ = _0016_ ? addroundkey_data_o[13] : _1026_;
  assign next_addroundkey_data_reg[13] = _0004_ ? _1023_ : _1027_;
  assign _1028_ = ~key_i[14];
  assign _1029_ = ~subbytes_data_o[14];
  assign _1030_ = ~mixcol_data_o[14];
  assign _1031_ = ~data_i[14];
  assign _1032_ = _0459_ ? _1030_ : _1031_;
  assign _1033_ = _0455_ ? _1029_ : _1032_;
  assign _1034_ = _0470_ ? _1029_ : _1033_;
  assign _1035_ = _0469_ ? _1030_ : _1034_;
  assign _1036_ = subbytes_ready_o ? _1029_ : _1035_;
  assign _1037_ = _0468_ ? _1035_ : _1036_;
  assign _1038_ = _0463_ ? _1029_ : _1037_;
  assign _1039_ = _0450_ ? _1033_ : _1038_;
  assign _1040_ = _1039_ ^ _1028_;
  assign _1041_ = ~keysched_new_key_o[14];
  assign _1042_ = _1039_ ^ _1041_;
  assign _1043_ = _0479_ ? addroundkey_data_o[14] : _1042_;
  assign _1044_ = _0016_ ? addroundkey_data_o[14] : _1043_;
  assign next_addroundkey_data_reg[14] = _0004_ ? _1040_ : _1044_;
  assign _1045_ = ~key_i[15];
  assign _1046_ = ~subbytes_data_o[15];
  assign _1047_ = ~mixcol_data_o[15];
  assign _1048_ = ~data_i[15];
  assign _1049_ = _0459_ ? _1047_ : _1048_;
  assign _1050_ = _0455_ ? _1046_ : _1049_;
  assign _1051_ = _0470_ ? _1046_ : _1050_;
  assign _1052_ = _0469_ ? _1047_ : _1051_;
  assign _1053_ = subbytes_ready_o ? _1046_ : _1052_;
  assign _1054_ = _0468_ ? _1052_ : _1053_;
  assign _1055_ = _0463_ ? _1046_ : _1054_;
  assign _1056_ = _0450_ ? _1050_ : _1055_;
  assign _1057_ = _1056_ ^ _1045_;
  assign _1058_ = ~keysched_new_key_o[15];
  assign _1059_ = _1056_ ^ _1058_;
  assign _1060_ = _0479_ ? addroundkey_data_o[15] : _1059_;
  assign _1061_ = _0016_ ? addroundkey_data_o[15] : _1060_;
  assign next_addroundkey_data_reg[15] = _0004_ ? _1057_ : _1061_;
  assign _1062_ = ~key_i[16];
  assign _1063_ = ~subbytes_data_o[16];
  assign _1064_ = ~mixcol_data_o[16];
  assign _1065_ = ~data_i[16];
  assign _1066_ = _0459_ ? _1064_ : _1065_;
  assign _1067_ = _0455_ ? _1063_ : _1066_;
  assign _1068_ = _0470_ ? _1063_ : _1067_;
  assign _1069_ = _0469_ ? _1064_ : _1068_;
  assign _1070_ = subbytes_ready_o ? _1063_ : _1069_;
  assign _1071_ = _0468_ ? _1069_ : _1070_;
  assign _1072_ = _0463_ ? _1063_ : _1071_;
  assign _1073_ = _0450_ ? _1067_ : _1072_;
  assign _1074_ = _1073_ ^ _1062_;
  assign _1075_ = ~keysched_new_key_o[16];
  assign _1076_ = _1073_ ^ _1075_;
  assign _1077_ = _0479_ ? addroundkey_data_o[16] : _1076_;
  assign _1078_ = _0016_ ? addroundkey_data_o[16] : _1077_;
  assign next_addroundkey_data_reg[16] = _0004_ ? _1074_ : _1078_;
  assign _1079_ = ~key_i[17];
  assign _1080_ = ~subbytes_data_o[17];
  assign _1081_ = ~mixcol_data_o[17];
  assign _1082_ = ~data_i[17];
  assign _1083_ = _0459_ ? _1081_ : _1082_;
  assign _1084_ = _0455_ ? _1080_ : _1083_;
  assign _1085_ = _0470_ ? _1080_ : _1084_;
  assign _1086_ = _0469_ ? _1081_ : _1085_;
  assign _1087_ = subbytes_ready_o ? _1080_ : _1086_;
  assign _1088_ = _0468_ ? _1086_ : _1087_;
  assign _1089_ = _0463_ ? _1080_ : _1088_;
  assign _1090_ = _0450_ ? _1084_ : _1089_;
  assign _1091_ = _1090_ ^ _1079_;
  assign _1092_ = ~keysched_new_key_o[17];
  assign _1093_ = _1090_ ^ _1092_;
  assign _1094_ = _0479_ ? addroundkey_data_o[17] : _1093_;
  assign _1095_ = _0016_ ? addroundkey_data_o[17] : _1094_;
  assign next_addroundkey_data_reg[17] = _0004_ ? _1091_ : _1095_;
  assign _1096_ = ~key_i[18];
  assign _1097_ = ~subbytes_data_o[18];
  assign _1098_ = ~mixcol_data_o[18];
  assign _1099_ = ~data_i[18];
  assign _1100_ = _0459_ ? _1098_ : _1099_;
  assign _1101_ = _0455_ ? _1097_ : _1100_;
  assign _1102_ = _0470_ ? _1097_ : _1101_;
  assign _1103_ = _0469_ ? _1098_ : _1102_;
  assign _1104_ = subbytes_ready_o ? _1097_ : _1103_;
  assign _1105_ = _0468_ ? _1103_ : _1104_;
  assign _1106_ = _0463_ ? _1097_ : _1105_;
  assign _1107_ = _0450_ ? _1101_ : _1106_;
  assign _1108_ = _1107_ ^ _1096_;
  assign _1109_ = ~keysched_new_key_o[18];
  assign _1110_ = _1107_ ^ _1109_;
  assign _1111_ = _0479_ ? addroundkey_data_o[18] : _1110_;
  assign _1112_ = _0016_ ? addroundkey_data_o[18] : _1111_;
  assign next_addroundkey_data_reg[18] = _0004_ ? _1108_ : _1112_;
  assign _1113_ = ~key_i[19];
  assign _1114_ = ~subbytes_data_o[19];
  assign _1115_ = ~mixcol_data_o[19];
  assign _1116_ = ~data_i[19];
  assign _1117_ = _0459_ ? _1115_ : _1116_;
  assign _1118_ = _0455_ ? _1114_ : _1117_;
  assign _1119_ = _0470_ ? _1114_ : _1118_;
  assign _1120_ = _0469_ ? _1115_ : _1119_;
  assign _1121_ = subbytes_ready_o ? _1114_ : _1120_;
  assign _1122_ = _0468_ ? _1120_ : _1121_;
  assign _1123_ = _0463_ ? _1114_ : _1122_;
  assign _1124_ = _0450_ ? _1118_ : _1123_;
  assign _1125_ = _1124_ ^ _1113_;
  assign _1126_ = ~keysched_new_key_o[19];
  assign _1127_ = _1124_ ^ _1126_;
  assign _1128_ = _0479_ ? addroundkey_data_o[19] : _1127_;
  assign _1129_ = _0016_ ? addroundkey_data_o[19] : _1128_;
  assign next_addroundkey_data_reg[19] = _0004_ ? _1125_ : _1129_;
  assign _1130_ = ~key_i[1];
  assign _1131_ = ~subbytes_data_o[1];
  assign _1132_ = ~mixcol_data_o[1];
  assign _1133_ = ~data_i[1];
  assign _1134_ = _0459_ ? _1132_ : _1133_;
  assign _1135_ = _0455_ ? _1131_ : _1134_;
  assign _1136_ = _0470_ ? _1131_ : _1135_;
  assign _1137_ = _0469_ ? _1132_ : _1136_;
  assign _1138_ = subbytes_ready_o ? _1131_ : _1137_;
  assign _1139_ = _0468_ ? _1137_ : _1138_;
  assign _1140_ = _0463_ ? _1131_ : _1139_;
  assign _1141_ = _0450_ ? _1135_ : _1140_;
  assign _1142_ = _1141_ ^ _1130_;
  assign _1143_ = ~keysched_new_key_o[1];
  assign _1144_ = _1141_ ^ _1143_;
  assign _1145_ = _0479_ ? addroundkey_data_o[1] : _1144_;
  assign _1146_ = _0016_ ? addroundkey_data_o[1] : _1145_;
  assign next_addroundkey_data_reg[1] = _0004_ ? _1142_ : _1146_;
  assign _1147_ = ~key_i[20];
  assign _1148_ = ~subbytes_data_o[20];
  assign _1149_ = ~mixcol_data_o[20];
  assign _1150_ = ~data_i[20];
  assign _1151_ = _0459_ ? _1149_ : _1150_;
  assign _1152_ = _0455_ ? _1148_ : _1151_;
  assign _1153_ = _0470_ ? _1148_ : _1152_;
  assign _1154_ = _0469_ ? _1149_ : _1153_;
  assign _1155_ = subbytes_ready_o ? _1148_ : _1154_;
  assign _1156_ = _0468_ ? _1154_ : _1155_;
  assign _1157_ = _0463_ ? _1148_ : _1156_;
  assign _1158_ = _0450_ ? _1152_ : _1157_;
  assign _1159_ = _1158_ ^ _1147_;
  assign _1160_ = ~keysched_new_key_o[20];
  assign _1161_ = _1158_ ^ _1160_;
  assign _1162_ = _0479_ ? addroundkey_data_o[20] : _1161_;
  assign _1163_ = _0016_ ? addroundkey_data_o[20] : _1162_;
  assign next_addroundkey_data_reg[20] = _0004_ ? _1159_ : _1163_;
  assign _1164_ = ~key_i[21];
  assign _1165_ = ~subbytes_data_o[21];
  assign _1166_ = ~mixcol_data_o[21];
  assign _1167_ = ~data_i[21];
  assign _1168_ = _0459_ ? _1166_ : _1167_;
  assign _1169_ = _0455_ ? _1165_ : _1168_;
  assign _1170_ = _0470_ ? _1165_ : _1169_;
  assign _1171_ = _0469_ ? _1166_ : _1170_;
  assign _1172_ = subbytes_ready_o ? _1165_ : _1171_;
  assign _1173_ = _0468_ ? _1171_ : _1172_;
  assign _1174_ = _0463_ ? _1165_ : _1173_;
  assign _1175_ = _0450_ ? _1169_ : _1174_;
  assign _1176_ = _1175_ ^ _1164_;
  assign _1177_ = ~keysched_new_key_o[21];
  assign _1178_ = _1175_ ^ _1177_;
  assign _1179_ = _0479_ ? addroundkey_data_o[21] : _1178_;
  assign _1180_ = _0016_ ? addroundkey_data_o[21] : _1179_;
  assign next_addroundkey_data_reg[21] = _0004_ ? _1176_ : _1180_;
  assign _1181_ = ~key_i[22];
  assign _1182_ = ~subbytes_data_o[22];
  assign _1183_ = ~mixcol_data_o[22];
  assign _1184_ = ~data_i[22];
  assign _1185_ = _0459_ ? _1183_ : _1184_;
  assign _1186_ = _0455_ ? _1182_ : _1185_;
  assign _1187_ = _0470_ ? _1182_ : _1186_;
  assign _1188_ = _0469_ ? _1183_ : _1187_;
  assign _1189_ = subbytes_ready_o ? _1182_ : _1188_;
  assign _1190_ = _0468_ ? _1188_ : _1189_;
  assign _1191_ = _0463_ ? _1182_ : _1190_;
  assign _1192_ = _0450_ ? _1186_ : _1191_;
  assign _1193_ = _1192_ ^ _1181_;
  assign _1194_ = ~keysched_new_key_o[22];
  assign _1195_ = _1192_ ^ _1194_;
  assign _1196_ = _0479_ ? addroundkey_data_o[22] : _1195_;
  assign _1197_ = _0016_ ? addroundkey_data_o[22] : _1196_;
  assign next_addroundkey_data_reg[22] = _0004_ ? _1193_ : _1197_;
  assign _1198_ = ~key_i[23];
  assign _1199_ = ~subbytes_data_o[23];
  assign _1200_ = ~mixcol_data_o[23];
  assign _1201_ = ~data_i[23];
  assign _1202_ = _0459_ ? _1200_ : _1201_;
  assign _1203_ = _0455_ ? _1199_ : _1202_;
  assign _1204_ = _0470_ ? _1199_ : _1203_;
  assign _1205_ = _0469_ ? _1200_ : _1204_;
  assign _1206_ = subbytes_ready_o ? _1199_ : _1205_;
  assign _1207_ = _0468_ ? _1205_ : _1206_;
  assign _1208_ = _0463_ ? _1199_ : _1207_;
  assign _1209_ = _0450_ ? _1203_ : _1208_;
  assign _1210_ = _1209_ ^ _1198_;
  assign _1211_ = ~keysched_new_key_o[23];
  assign _1212_ = _1209_ ^ _1211_;
  assign _1213_ = _0479_ ? addroundkey_data_o[23] : _1212_;
  assign _1214_ = _0016_ ? addroundkey_data_o[23] : _1213_;
  assign next_addroundkey_data_reg[23] = _0004_ ? _1210_ : _1214_;
  assign _1215_ = ~key_i[24];
  assign _1216_ = ~subbytes_data_o[24];
  assign _1217_ = ~mixcol_data_o[24];
  assign _1218_ = ~data_i[24];
  assign _1219_ = _0459_ ? _1217_ : _1218_;
  assign _1220_ = _0455_ ? _1216_ : _1219_;
  assign _1221_ = _0470_ ? _1216_ : _1220_;
  assign _1222_ = _0469_ ? _1217_ : _1221_;
  assign _1223_ = subbytes_ready_o ? _1216_ : _1222_;
  assign _1224_ = _0468_ ? _1222_ : _1223_;
  assign _1225_ = _0463_ ? _1216_ : _1224_;
  assign _1226_ = _0450_ ? _1220_ : _1225_;
  assign _1227_ = _1226_ ^ _1215_;
  assign _1228_ = ~keysched_new_key_o[24];
  assign _1229_ = _1226_ ^ _1228_;
  assign _1230_ = _0479_ ? addroundkey_data_o[24] : _1229_;
  assign _1231_ = _0016_ ? addroundkey_data_o[24] : _1230_;
  assign next_addroundkey_data_reg[24] = _0004_ ? _1227_ : _1231_;
  assign _1232_ = ~key_i[25];
  assign _1233_ = ~subbytes_data_o[25];
  assign _1234_ = ~mixcol_data_o[25];
  assign _1235_ = ~data_i[25];
  assign _1236_ = _0459_ ? _1234_ : _1235_;
  assign _1237_ = _0455_ ? _1233_ : _1236_;
  assign _1238_ = _0470_ ? _1233_ : _1237_;
  assign _1239_ = _0469_ ? _1234_ : _1238_;
  assign _1240_ = subbytes_ready_o ? _1233_ : _1239_;
  assign _1241_ = _0468_ ? _1239_ : _1240_;
  assign _1242_ = _0463_ ? _1233_ : _1241_;
  assign _1243_ = _0450_ ? _1237_ : _1242_;
  assign _1244_ = _1243_ ^ _1232_;
  assign _1245_ = ~keysched_new_key_o[25];
  assign _1246_ = _1243_ ^ _1245_;
  assign _1247_ = _0479_ ? addroundkey_data_o[25] : _1246_;
  assign _1248_ = _0016_ ? addroundkey_data_o[25] : _1247_;
  assign next_addroundkey_data_reg[25] = _0004_ ? _1244_ : _1248_;
  assign _1249_ = ~key_i[26];
  assign _1250_ = ~subbytes_data_o[26];
  assign _1251_ = ~mixcol_data_o[26];
  assign _1252_ = ~data_i[26];
  assign _1253_ = _0459_ ? _1251_ : _1252_;
  assign _1254_ = _0455_ ? _1250_ : _1253_;
  assign _1255_ = _0470_ ? _1250_ : _1254_;
  assign _1256_ = _0469_ ? _1251_ : _1255_;
  assign _1257_ = subbytes_ready_o ? _1250_ : _1256_;
  assign _1258_ = _0468_ ? _1256_ : _1257_;
  assign _1259_ = _0463_ ? _1250_ : _1258_;
  assign _1260_ = _0450_ ? _1254_ : _1259_;
  assign _1261_ = _1260_ ^ _1249_;
  assign _1262_ = ~keysched_new_key_o[26];
  assign _1263_ = _1260_ ^ _1262_;
  assign _1264_ = _0479_ ? addroundkey_data_o[26] : _1263_;
  assign _1265_ = _0016_ ? addroundkey_data_o[26] : _1264_;
  assign next_addroundkey_data_reg[26] = _0004_ ? _1261_ : _1265_;
  assign _1266_ = ~key_i[27];
  assign _1267_ = ~subbytes_data_o[27];
  assign _1268_ = ~mixcol_data_o[27];
  assign _1269_ = ~data_i[27];
  assign _1270_ = _0459_ ? _1268_ : _1269_;
  assign _1271_ = _0455_ ? _1267_ : _1270_;
  assign _1272_ = _0470_ ? _1267_ : _1271_;
  assign _1273_ = _0469_ ? _1268_ : _1272_;
  assign _1274_ = subbytes_ready_o ? _1267_ : _1273_;
  assign _1275_ = _0468_ ? _1273_ : _1274_;
  assign _1276_ = _0463_ ? _1267_ : _1275_;
  assign _1277_ = _0450_ ? _1271_ : _1276_;
  assign _1278_ = _1277_ ^ _1266_;
  assign _1279_ = ~keysched_new_key_o[27];
  assign _1280_ = _1277_ ^ _1279_;
  assign _1281_ = _0479_ ? addroundkey_data_o[27] : _1280_;
  assign _1282_ = _0016_ ? addroundkey_data_o[27] : _1281_;
  assign next_addroundkey_data_reg[27] = _0004_ ? _1278_ : _1282_;
  assign _1283_ = ~key_i[28];
  assign _1284_ = ~subbytes_data_o[28];
  assign _1285_ = ~mixcol_data_o[28];
  assign _1286_ = ~data_i[28];
  assign _1287_ = _0459_ ? _1285_ : _1286_;
  assign _1288_ = _0455_ ? _1284_ : _1287_;
  assign _1289_ = _0470_ ? _1284_ : _1288_;
  assign _1290_ = _0469_ ? _1285_ : _1289_;
  assign _1291_ = subbytes_ready_o ? _1284_ : _1290_;
  assign _1292_ = _0468_ ? _1290_ : _1291_;
  assign _1293_ = _0463_ ? _1284_ : _1292_;
  assign _1294_ = _0450_ ? _1288_ : _1293_;
  assign _1295_ = _1294_ ^ _1283_;
  assign _1296_ = ~keysched_new_key_o[28];
  assign _1297_ = _1294_ ^ _1296_;
  assign _1298_ = _0479_ ? addroundkey_data_o[28] : _1297_;
  assign _1299_ = _0016_ ? addroundkey_data_o[28] : _1298_;
  assign next_addroundkey_data_reg[28] = _0004_ ? _1295_ : _1299_;
  assign _1300_ = ~key_i[29];
  assign _1301_ = ~subbytes_data_o[29];
  assign _1302_ = ~mixcol_data_o[29];
  assign _1303_ = ~data_i[29];
  assign _1304_ = _0459_ ? _1302_ : _1303_;
  assign _1305_ = _0455_ ? _1301_ : _1304_;
  assign _1306_ = _0470_ ? _1301_ : _1305_;
  assign _1307_ = _0469_ ? _1302_ : _1306_;
  assign _1308_ = subbytes_ready_o ? _1301_ : _1307_;
  assign _1309_ = _0468_ ? _1307_ : _1308_;
  assign _1310_ = _0463_ ? _1301_ : _1309_;
  assign _1311_ = _0450_ ? _1305_ : _1310_;
  assign _1312_ = _1311_ ^ _1300_;
  assign _1313_ = ~keysched_new_key_o[29];
  assign _1314_ = _1311_ ^ _1313_;
  assign _1315_ = _0479_ ? addroundkey_data_o[29] : _1314_;
  assign _1316_ = _0016_ ? addroundkey_data_o[29] : _1315_;
  assign next_addroundkey_data_reg[29] = _0004_ ? _1312_ : _1316_;
  assign _1317_ = ~key_i[2];
  assign _1318_ = ~subbytes_data_o[2];
  assign _1319_ = ~mixcol_data_o[2];
  assign _1320_ = ~data_i[2];
  assign _1321_ = _0459_ ? _1319_ : _1320_;
  assign _1322_ = _0455_ ? _1318_ : _1321_;
  assign _1323_ = _0470_ ? _1318_ : _1322_;
  assign _1324_ = _0469_ ? _1319_ : _1323_;
  assign _1325_ = subbytes_ready_o ? _1318_ : _1324_;
  assign _1326_ = _0468_ ? _1324_ : _1325_;
  assign _1327_ = _0463_ ? _1318_ : _1326_;
  assign _1328_ = _0450_ ? _1322_ : _1327_;
  assign _1329_ = _1328_ ^ _1317_;
  assign _1330_ = ~keysched_new_key_o[2];
  assign _1331_ = _1328_ ^ _1330_;
  assign _1332_ = _0479_ ? addroundkey_data_o[2] : _1331_;
  assign _1333_ = _0016_ ? addroundkey_data_o[2] : _1332_;
  assign next_addroundkey_data_reg[2] = _0004_ ? _1329_ : _1333_;
  assign _1334_ = ~key_i[30];
  assign _1335_ = ~subbytes_data_o[30];
  assign _1336_ = ~mixcol_data_o[30];
  assign _1337_ = ~data_i[30];
  assign _1338_ = _0459_ ? _1336_ : _1337_;
  assign _1339_ = _0455_ ? _1335_ : _1338_;
  assign _1340_ = _0470_ ? _1335_ : _1339_;
  assign _1341_ = _0469_ ? _1336_ : _1340_;
  assign _1342_ = subbytes_ready_o ? _1335_ : _1341_;
  assign _1343_ = _0468_ ? _1341_ : _1342_;
  assign _1344_ = _0463_ ? _1335_ : _1343_;
  assign _1345_ = _0450_ ? _1339_ : _1344_;
  assign _1346_ = _1345_ ^ _1334_;
  assign _1347_ = ~keysched_new_key_o[30];
  assign _1348_ = _1345_ ^ _1347_;
  assign _1349_ = _0479_ ? addroundkey_data_o[30] : _1348_;
  assign _1350_ = _0016_ ? addroundkey_data_o[30] : _1349_;
  assign next_addroundkey_data_reg[30] = _0004_ ? _1346_ : _1350_;
  assign _1351_ = ~key_i[31];
  assign _1352_ = ~subbytes_data_o[31];
  assign _1353_ = ~mixcol_data_o[31];
  assign _1354_ = ~data_i[31];
  assign _1355_ = _0459_ ? _1353_ : _1354_;
  assign _1356_ = _0455_ ? _1352_ : _1355_;
  assign _1357_ = _0470_ ? _1352_ : _1356_;
  assign _1358_ = _0469_ ? _1353_ : _1357_;
  assign _1359_ = subbytes_ready_o ? _1352_ : _1358_;
  assign _1360_ = _0468_ ? _1358_ : _1359_;
  assign _1361_ = _0463_ ? _1352_ : _1360_;
  assign _1362_ = _0450_ ? _1356_ : _1361_;
  assign _1363_ = _1362_ ^ _1351_;
  assign _1364_ = ~keysched_new_key_o[31];
  assign _1365_ = _1362_ ^ _1364_;
  assign _1366_ = _0479_ ? addroundkey_data_o[31] : _1365_;
  assign _1367_ = _0016_ ? addroundkey_data_o[31] : _1366_;
  assign next_addroundkey_data_reg[31] = _0004_ ? _1363_ : _1367_;
  assign _1368_ = ~key_i[32];
  assign _1369_ = ~subbytes_data_o[32];
  assign _1370_ = ~mixcol_data_o[32];
  assign _1371_ = ~data_i[32];
  assign _1372_ = _0459_ ? _1370_ : _1371_;
  assign _1373_ = _0455_ ? _1369_ : _1372_;
  assign _1374_ = _0470_ ? _1369_ : _1373_;
  assign _1375_ = _0469_ ? _1370_ : _1374_;
  assign _1376_ = subbytes_ready_o ? _1369_ : _1375_;
  assign _1377_ = _0468_ ? _1375_ : _1376_;
  assign _1378_ = _0463_ ? _1369_ : _1377_;
  assign _1379_ = _0450_ ? _1373_ : _1378_;
  assign _1380_ = _1379_ ^ _1368_;
  assign _1381_ = ~keysched_new_key_o[32];
  assign _1382_ = _1379_ ^ _1381_;
  assign _1383_ = _0479_ ? addroundkey_data_o[32] : _1382_;
  assign _1384_ = _0016_ ? addroundkey_data_o[32] : _1383_;
  assign next_addroundkey_data_reg[32] = _0004_ ? _1380_ : _1384_;
  assign _1385_ = ~key_i[33];
  assign _1386_ = ~subbytes_data_o[33];
  assign _1387_ = ~mixcol_data_o[33];
  assign _1388_ = ~data_i[33];
  assign _1389_ = _0459_ ? _1387_ : _1388_;
  assign _1390_ = _0455_ ? _1386_ : _1389_;
  assign _1391_ = _0470_ ? _1386_ : _1390_;
  assign _1392_ = _0469_ ? _1387_ : _1391_;
  assign _1393_ = subbytes_ready_o ? _1386_ : _1392_;
  assign _1394_ = _0468_ ? _1392_ : _1393_;
  assign _1395_ = _0463_ ? _1386_ : _1394_;
  assign _1396_ = _0450_ ? _1390_ : _1395_;
  assign _1397_ = _1396_ ^ _1385_;
  assign _1398_ = ~keysched_new_key_o[33];
  assign _1399_ = _1396_ ^ _1398_;
  assign _1400_ = _0479_ ? addroundkey_data_o[33] : _1399_;
  assign _1401_ = _0016_ ? addroundkey_data_o[33] : _1400_;
  assign next_addroundkey_data_reg[33] = _0004_ ? _1397_ : _1401_;
  assign _1402_ = ~key_i[34];
  assign _1403_ = ~subbytes_data_o[34];
  assign _1404_ = ~mixcol_data_o[34];
  assign _1405_ = ~data_i[34];
  assign _1406_ = _0459_ ? _1404_ : _1405_;
  assign _1407_ = _0455_ ? _1403_ : _1406_;
  assign _1408_ = _0470_ ? _1403_ : _1407_;
  assign _1409_ = _0469_ ? _1404_ : _1408_;
  assign _1410_ = subbytes_ready_o ? _1403_ : _1409_;
  assign _1411_ = _0468_ ? _1409_ : _1410_;
  assign _1412_ = _0463_ ? _1403_ : _1411_;
  assign _1413_ = _0450_ ? _1407_ : _1412_;
  assign _1414_ = _1413_ ^ _1402_;
  assign _1415_ = ~keysched_new_key_o[34];
  assign _1416_ = _1413_ ^ _1415_;
  assign _1417_ = _0479_ ? addroundkey_data_o[34] : _1416_;
  assign _1418_ = _0016_ ? addroundkey_data_o[34] : _1417_;
  assign next_addroundkey_data_reg[34] = _0004_ ? _1414_ : _1418_;
  assign _1419_ = ~key_i[35];
  assign _1420_ = ~subbytes_data_o[35];
  assign _1421_ = ~mixcol_data_o[35];
  assign _1422_ = ~data_i[35];
  assign _1423_ = _0459_ ? _1421_ : _1422_;
  assign _1424_ = _0455_ ? _1420_ : _1423_;
  assign _1425_ = _0470_ ? _1420_ : _1424_;
  assign _1426_ = _0469_ ? _1421_ : _1425_;
  assign _1427_ = subbytes_ready_o ? _1420_ : _1426_;
  assign _1428_ = _0468_ ? _1426_ : _1427_;
  assign _1429_ = _0463_ ? _1420_ : _1428_;
  assign _1430_ = _0450_ ? _1424_ : _1429_;
  assign _1431_ = _1430_ ^ _1419_;
  assign _1432_ = ~keysched_new_key_o[35];
  assign _1433_ = _1430_ ^ _1432_;
  assign _1434_ = _0479_ ? addroundkey_data_o[35] : _1433_;
  assign _1435_ = _0016_ ? addroundkey_data_o[35] : _1434_;
  assign next_addroundkey_data_reg[35] = _0004_ ? _1431_ : _1435_;
  assign _1436_ = ~key_i[36];
  assign _1437_ = ~subbytes_data_o[36];
  assign _1438_ = ~mixcol_data_o[36];
  assign _1439_ = ~data_i[36];
  assign _1440_ = _0459_ ? _1438_ : _1439_;
  assign _1441_ = _0455_ ? _1437_ : _1440_;
  assign _1442_ = _0470_ ? _1437_ : _1441_;
  assign _1443_ = _0469_ ? _1438_ : _1442_;
  assign _1444_ = subbytes_ready_o ? _1437_ : _1443_;
  assign _1445_ = _0468_ ? _1443_ : _1444_;
  assign _1446_ = _0463_ ? _1437_ : _1445_;
  assign _1447_ = _0450_ ? _1441_ : _1446_;
  assign _1448_ = _1447_ ^ _1436_;
  assign _1449_ = ~keysched_new_key_o[36];
  assign _1450_ = _1447_ ^ _1449_;
  assign _1451_ = _0479_ ? addroundkey_data_o[36] : _1450_;
  assign _1452_ = _0016_ ? addroundkey_data_o[36] : _1451_;
  assign next_addroundkey_data_reg[36] = _0004_ ? _1448_ : _1452_;
  assign _1453_ = ~key_i[37];
  assign _1454_ = ~subbytes_data_o[37];
  assign _1455_ = ~mixcol_data_o[37];
  assign _1456_ = ~data_i[37];
  assign _1457_ = _0459_ ? _1455_ : _1456_;
  assign _1458_ = _0455_ ? _1454_ : _1457_;
  assign _1459_ = _0470_ ? _1454_ : _1458_;
  assign _1460_ = _0469_ ? _1455_ : _1459_;
  assign _1461_ = subbytes_ready_o ? _1454_ : _1460_;
  assign _1462_ = _0468_ ? _1460_ : _1461_;
  assign _1463_ = _0463_ ? _1454_ : _1462_;
  assign _1464_ = _0450_ ? _1458_ : _1463_;
  assign _1465_ = _1464_ ^ _1453_;
  assign _1466_ = ~keysched_new_key_o[37];
  assign _1467_ = _1464_ ^ _1466_;
  assign _1468_ = _0479_ ? addroundkey_data_o[37] : _1467_;
  assign _1469_ = _0016_ ? addroundkey_data_o[37] : _1468_;
  assign next_addroundkey_data_reg[37] = _0004_ ? _1465_ : _1469_;
  assign _1470_ = ~key_i[38];
  assign _1471_ = ~subbytes_data_o[38];
  assign _1472_ = ~mixcol_data_o[38];
  assign _1473_ = ~data_i[38];
  assign _1474_ = _0459_ ? _1472_ : _1473_;
  assign _1475_ = _0455_ ? _1471_ : _1474_;
  assign _1476_ = _0470_ ? _1471_ : _1475_;
  assign _1477_ = _0469_ ? _1472_ : _1476_;
  assign _1478_ = subbytes_ready_o ? _1471_ : _1477_;
  assign _1479_ = _0468_ ? _1477_ : _1478_;
  assign _1480_ = _0463_ ? _1471_ : _1479_;
  assign _1481_ = _0450_ ? _1475_ : _1480_;
  assign _1482_ = _1481_ ^ _1470_;
  assign _1483_ = ~keysched_new_key_o[38];
  assign _1484_ = _1481_ ^ _1483_;
  assign _1485_ = _0479_ ? addroundkey_data_o[38] : _1484_;
  assign _1486_ = _0016_ ? addroundkey_data_o[38] : _1485_;
  assign next_addroundkey_data_reg[38] = _0004_ ? _1482_ : _1486_;
  assign _1487_ = ~key_i[39];
  assign _1488_ = ~subbytes_data_o[39];
  assign _1489_ = ~mixcol_data_o[39];
  assign _1490_ = ~data_i[39];
  assign _1491_ = _0459_ ? _1489_ : _1490_;
  assign _1492_ = _0455_ ? _1488_ : _1491_;
  assign _1493_ = _0470_ ? _1488_ : _1492_;
  assign _1494_ = _0469_ ? _1489_ : _1493_;
  assign _1495_ = subbytes_ready_o ? _1488_ : _1494_;
  assign _1496_ = _0468_ ? _1494_ : _1495_;
  assign _1497_ = _0463_ ? _1488_ : _1496_;
  assign _1498_ = _0450_ ? _1492_ : _1497_;
  assign _1499_ = _1498_ ^ _1487_;
  assign _1500_ = ~keysched_new_key_o[39];
  assign _1501_ = _1498_ ^ _1500_;
  assign _1502_ = _0479_ ? addroundkey_data_o[39] : _1501_;
  assign _1503_ = _0016_ ? addroundkey_data_o[39] : _1502_;
  assign next_addroundkey_data_reg[39] = _0004_ ? _1499_ : _1503_;
  assign _1504_ = ~key_i[3];
  assign _1505_ = ~subbytes_data_o[3];
  assign _1506_ = ~mixcol_data_o[3];
  assign _1507_ = ~data_i[3];
  assign _1508_ = _0459_ ? _1506_ : _1507_;
  assign _1509_ = _0455_ ? _1505_ : _1508_;
  assign _1510_ = _0470_ ? _1505_ : _1509_;
  assign _1511_ = _0469_ ? _1506_ : _1510_;
  assign _1512_ = subbytes_ready_o ? _1505_ : _1511_;
  assign _1513_ = _0468_ ? _1511_ : _1512_;
  assign _1514_ = _0463_ ? _1505_ : _1513_;
  assign _1515_ = _0450_ ? _1509_ : _1514_;
  assign _1516_ = _1515_ ^ _1504_;
  assign _1517_ = ~keysched_new_key_o[3];
  assign _1518_ = _1515_ ^ _1517_;
  assign _1519_ = _0479_ ? addroundkey_data_o[3] : _1518_;
  assign _1520_ = _0016_ ? addroundkey_data_o[3] : _1519_;
  assign next_addroundkey_data_reg[3] = _0004_ ? _1516_ : _1520_;
  assign _1521_ = ~key_i[40];
  assign _1522_ = ~subbytes_data_o[40];
  assign _1523_ = ~mixcol_data_o[40];
  assign _1524_ = ~data_i[40];
  assign _1525_ = _0459_ ? _1523_ : _1524_;
  assign _1526_ = _0455_ ? _1522_ : _1525_;
  assign _1527_ = _0470_ ? _1522_ : _1526_;
  assign _1528_ = _0469_ ? _1523_ : _1527_;
  assign _1529_ = subbytes_ready_o ? _1522_ : _1528_;
  assign _1530_ = _0468_ ? _1528_ : _1529_;
  assign _1531_ = _0463_ ? _1522_ : _1530_;
  assign _1532_ = _0450_ ? _1526_ : _1531_;
  assign _1533_ = _1532_ ^ _1521_;
  assign _1534_ = ~keysched_new_key_o[40];
  assign _1535_ = _1532_ ^ _1534_;
  assign _1536_ = _0479_ ? addroundkey_data_o[40] : _1535_;
  assign _1537_ = _0016_ ? addroundkey_data_o[40] : _1536_;
  assign next_addroundkey_data_reg[40] = _0004_ ? _1533_ : _1537_;
  assign _1538_ = ~key_i[41];
  assign _1539_ = ~subbytes_data_o[41];
  assign _1540_ = ~mixcol_data_o[41];
  assign _1541_ = ~data_i[41];
  assign _1542_ = _0459_ ? _1540_ : _1541_;
  assign _1543_ = _0455_ ? _1539_ : _1542_;
  assign _1544_ = _0470_ ? _1539_ : _1543_;
  assign _1545_ = _0469_ ? _1540_ : _1544_;
  assign _1546_ = subbytes_ready_o ? _1539_ : _1545_;
  assign _1547_ = _0468_ ? _1545_ : _1546_;
  assign _1548_ = _0463_ ? _1539_ : _1547_;
  assign _1549_ = _0450_ ? _1543_ : _1548_;
  assign _1550_ = _1549_ ^ _1538_;
  assign _1551_ = ~keysched_new_key_o[41];
  assign _1552_ = _1549_ ^ _1551_;
  assign _1553_ = _0479_ ? addroundkey_data_o[41] : _1552_;
  assign _1554_ = _0016_ ? addroundkey_data_o[41] : _1553_;
  assign next_addroundkey_data_reg[41] = _0004_ ? _1550_ : _1554_;
  assign _1555_ = ~key_i[42];
  assign _1556_ = ~subbytes_data_o[42];
  assign _1557_ = ~mixcol_data_o[42];
  assign _1558_ = ~data_i[42];
  assign _1559_ = _0459_ ? _1557_ : _1558_;
  assign _1560_ = _0455_ ? _1556_ : _1559_;
  assign _1561_ = _0470_ ? _1556_ : _1560_;
  assign _1562_ = _0469_ ? _1557_ : _1561_;
  assign _1563_ = subbytes_ready_o ? _1556_ : _1562_;
  assign _1564_ = _0468_ ? _1562_ : _1563_;
  assign _1565_ = _0463_ ? _1556_ : _1564_;
  assign _1566_ = _0450_ ? _1560_ : _1565_;
  assign _1567_ = _1566_ ^ _1555_;
  assign _1568_ = ~keysched_new_key_o[42];
  assign _1569_ = _1566_ ^ _1568_;
  assign _1570_ = _0479_ ? addroundkey_data_o[42] : _1569_;
  assign _1571_ = _0016_ ? addroundkey_data_o[42] : _1570_;
  assign next_addroundkey_data_reg[42] = _0004_ ? _1567_ : _1571_;
  assign _1572_ = ~key_i[43];
  assign _1573_ = ~subbytes_data_o[43];
  assign _1574_ = ~mixcol_data_o[43];
  assign _1575_ = ~data_i[43];
  assign _1576_ = _0459_ ? _1574_ : _1575_;
  assign _1577_ = _0455_ ? _1573_ : _1576_;
  assign _1578_ = _0470_ ? _1573_ : _1577_;
  assign _1579_ = _0469_ ? _1574_ : _1578_;
  assign _1580_ = subbytes_ready_o ? _1573_ : _1579_;
  assign _1581_ = _0468_ ? _1579_ : _1580_;
  assign _1582_ = _0463_ ? _1573_ : _1581_;
  assign _1583_ = _0450_ ? _1577_ : _1582_;
  assign _1584_ = _1583_ ^ _1572_;
  assign _1585_ = ~keysched_new_key_o[43];
  assign _1586_ = _1583_ ^ _1585_;
  assign _1587_ = _0479_ ? addroundkey_data_o[43] : _1586_;
  assign _1588_ = _0016_ ? addroundkey_data_o[43] : _1587_;
  assign next_addroundkey_data_reg[43] = _0004_ ? _1584_ : _1588_;
  assign _1589_ = ~key_i[44];
  assign _1590_ = ~subbytes_data_o[44];
  assign _1591_ = ~mixcol_data_o[44];
  assign _1592_ = ~data_i[44];
  assign _1593_ = _0459_ ? _1591_ : _1592_;
  assign _1594_ = _0455_ ? _1590_ : _1593_;
  assign _1595_ = _0470_ ? _1590_ : _1594_;
  assign _1596_ = _0469_ ? _1591_ : _1595_;
  assign _1597_ = subbytes_ready_o ? _1590_ : _1596_;
  assign _1598_ = _0468_ ? _1596_ : _1597_;
  assign _1599_ = _0463_ ? _1590_ : _1598_;
  assign _1600_ = _0450_ ? _1594_ : _1599_;
  assign _1601_ = _1600_ ^ _1589_;
  assign _1602_ = ~keysched_new_key_o[44];
  assign _1603_ = _1600_ ^ _1602_;
  assign _1604_ = _0479_ ? addroundkey_data_o[44] : _1603_;
  assign _1605_ = _0016_ ? addroundkey_data_o[44] : _1604_;
  assign next_addroundkey_data_reg[44] = _0004_ ? _1601_ : _1605_;
  assign _1606_ = ~key_i[45];
  assign _1607_ = ~subbytes_data_o[45];
  assign _1608_ = ~mixcol_data_o[45];
  assign _1609_ = ~data_i[45];
  assign _1610_ = _0459_ ? _1608_ : _1609_;
  assign _1611_ = _0455_ ? _1607_ : _1610_;
  assign _1612_ = _0470_ ? _1607_ : _1611_;
  assign _1613_ = _0469_ ? _1608_ : _1612_;
  assign _1614_ = subbytes_ready_o ? _1607_ : _1613_;
  assign _1615_ = _0468_ ? _1613_ : _1614_;
  assign _1616_ = _0463_ ? _1607_ : _1615_;
  assign _1617_ = _0450_ ? _1611_ : _1616_;
  assign _1618_ = _1617_ ^ _1606_;
  assign _1619_ = ~keysched_new_key_o[45];
  assign _1620_ = _1617_ ^ _1619_;
  assign _1621_ = _0479_ ? addroundkey_data_o[45] : _1620_;
  assign _1622_ = _0016_ ? addroundkey_data_o[45] : _1621_;
  assign next_addroundkey_data_reg[45] = _0004_ ? _1618_ : _1622_;
  assign _1623_ = ~key_i[46];
  assign _1624_ = ~subbytes_data_o[46];
  assign _1625_ = ~mixcol_data_o[46];
  assign _1626_ = ~data_i[46];
  assign _1627_ = _0459_ ? _1625_ : _1626_;
  assign _1628_ = _0455_ ? _1624_ : _1627_;
  assign _1629_ = _0470_ ? _1624_ : _1628_;
  assign _1630_ = _0469_ ? _1625_ : _1629_;
  assign _1631_ = subbytes_ready_o ? _1624_ : _1630_;
  assign _1632_ = _0468_ ? _1630_ : _1631_;
  assign _1633_ = _0463_ ? _1624_ : _1632_;
  assign _1634_ = _0450_ ? _1628_ : _1633_;
  assign _1635_ = _1634_ ^ _1623_;
  assign _1636_ = ~keysched_new_key_o[46];
  assign _1637_ = _1634_ ^ _1636_;
  assign _1638_ = _0479_ ? addroundkey_data_o[46] : _1637_;
  assign _1639_ = _0016_ ? addroundkey_data_o[46] : _1638_;
  assign next_addroundkey_data_reg[46] = _0004_ ? _1635_ : _1639_;
  assign _1640_ = ~key_i[47];
  assign _1641_ = ~subbytes_data_o[47];
  assign _1642_ = ~mixcol_data_o[47];
  assign _1643_ = ~data_i[47];
  assign _1644_ = _0459_ ? _1642_ : _1643_;
  assign _1645_ = _0455_ ? _1641_ : _1644_;
  assign _1646_ = _0470_ ? _1641_ : _1645_;
  assign _1647_ = _0469_ ? _1642_ : _1646_;
  assign _1648_ = subbytes_ready_o ? _1641_ : _1647_;
  assign _1649_ = _0468_ ? _1647_ : _1648_;
  assign _1650_ = _0463_ ? _1641_ : _1649_;
  assign _1651_ = _0450_ ? _1645_ : _1650_;
  assign _1652_ = _1651_ ^ _1640_;
  assign _1653_ = ~keysched_new_key_o[47];
  assign _1654_ = _1651_ ^ _1653_;
  assign _1655_ = _0479_ ? addroundkey_data_o[47] : _1654_;
  assign _1656_ = _0016_ ? addroundkey_data_o[47] : _1655_;
  assign next_addroundkey_data_reg[47] = _0004_ ? _1652_ : _1656_;
  assign _1657_ = ~key_i[48];
  assign _1658_ = ~subbytes_data_o[48];
  assign _1659_ = ~mixcol_data_o[48];
  assign _1660_ = ~data_i[48];
  assign _1661_ = _0459_ ? _1659_ : _1660_;
  assign _1662_ = _0455_ ? _1658_ : _1661_;
  assign _1663_ = _0470_ ? _1658_ : _1662_;
  assign _1664_ = _0469_ ? _1659_ : _1663_;
  assign _1665_ = subbytes_ready_o ? _1658_ : _1664_;
  assign _1666_ = _0468_ ? _1664_ : _1665_;
  assign _1667_ = _0463_ ? _1658_ : _1666_;
  assign _1668_ = _0450_ ? _1662_ : _1667_;
  assign _1669_ = _1668_ ^ _1657_;
  assign _1670_ = ~keysched_new_key_o[48];
  assign _1671_ = _1668_ ^ _1670_;
  assign _1672_ = _0479_ ? addroundkey_data_o[48] : _1671_;
  assign _1673_ = _0016_ ? addroundkey_data_o[48] : _1672_;
  assign next_addroundkey_data_reg[48] = _0004_ ? _1669_ : _1673_;
  assign _1674_ = ~key_i[49];
  assign _1675_ = ~subbytes_data_o[49];
  assign _1676_ = ~mixcol_data_o[49];
  assign _1677_ = ~data_i[49];
  assign _1678_ = _0459_ ? _1676_ : _1677_;
  assign _1679_ = _0455_ ? _1675_ : _1678_;
  assign _1680_ = _0470_ ? _1675_ : _1679_;
  assign _1681_ = _0469_ ? _1676_ : _1680_;
  assign _1682_ = subbytes_ready_o ? _1675_ : _1681_;
  assign _1683_ = _0468_ ? _1681_ : _1682_;
  assign _1684_ = _0463_ ? _1675_ : _1683_;
  assign _1685_ = _0450_ ? _1679_ : _1684_;
  assign _1686_ = _1685_ ^ _1674_;
  assign _1687_ = ~keysched_new_key_o[49];
  assign _1688_ = _1685_ ^ _1687_;
  assign _1689_ = _0479_ ? addroundkey_data_o[49] : _1688_;
  assign _1690_ = _0016_ ? addroundkey_data_o[49] : _1689_;
  assign next_addroundkey_data_reg[49] = _0004_ ? _1686_ : _1690_;
  assign _1691_ = ~key_i[4];
  assign _1692_ = ~subbytes_data_o[4];
  assign _1693_ = ~mixcol_data_o[4];
  assign _1694_ = ~data_i[4];
  assign _1695_ = _0459_ ? _1693_ : _1694_;
  assign _1696_ = _0455_ ? _1692_ : _1695_;
  assign _1697_ = _0470_ ? _1692_ : _1696_;
  assign _1698_ = _0469_ ? _1693_ : _1697_;
  assign _1699_ = subbytes_ready_o ? _1692_ : _1698_;
  assign _1700_ = _0468_ ? _1698_ : _1699_;
  assign _1701_ = _0463_ ? _1692_ : _1700_;
  assign _1702_ = _0450_ ? _1696_ : _1701_;
  assign _1703_ = _1702_ ^ _1691_;
  assign _1704_ = ~keysched_new_key_o[4];
  assign _1705_ = _1702_ ^ _1704_;
  assign _1706_ = _0479_ ? addroundkey_data_o[4] : _1705_;
  assign _1707_ = _0016_ ? addroundkey_data_o[4] : _1706_;
  assign next_addroundkey_data_reg[4] = _0004_ ? _1703_ : _1707_;
  assign _1708_ = ~key_i[50];
  assign _1709_ = ~subbytes_data_o[50];
  assign _1710_ = ~mixcol_data_o[50];
  assign _1711_ = ~data_i[50];
  assign _1712_ = _0459_ ? _1710_ : _1711_;
  assign _1713_ = _0455_ ? _1709_ : _1712_;
  assign _1714_ = _0470_ ? _1709_ : _1713_;
  assign _1715_ = _0469_ ? _1710_ : _1714_;
  assign _1716_ = subbytes_ready_o ? _1709_ : _1715_;
  assign _1717_ = _0468_ ? _1715_ : _1716_;
  assign _1718_ = _0463_ ? _1709_ : _1717_;
  assign _1719_ = _0450_ ? _1713_ : _1718_;
  assign _1720_ = _1719_ ^ _1708_;
  assign _1721_ = ~keysched_new_key_o[50];
  assign _1722_ = _1719_ ^ _1721_;
  assign _1723_ = _0479_ ? addroundkey_data_o[50] : _1722_;
  assign _1724_ = _0016_ ? addroundkey_data_o[50] : _1723_;
  assign next_addroundkey_data_reg[50] = _0004_ ? _1720_ : _1724_;
  assign _1725_ = ~key_i[51];
  assign _1726_ = ~subbytes_data_o[51];
  assign _1727_ = ~mixcol_data_o[51];
  assign _1728_ = ~data_i[51];
  assign _1729_ = _0459_ ? _1727_ : _1728_;
  assign _1730_ = _0455_ ? _1726_ : _1729_;
  assign _1731_ = _0470_ ? _1726_ : _1730_;
  assign _1732_ = _0469_ ? _1727_ : _1731_;
  assign _1733_ = subbytes_ready_o ? _1726_ : _1732_;
  assign _1734_ = _0468_ ? _1732_ : _1733_;
  assign _1735_ = _0463_ ? _1726_ : _1734_;
  assign _1736_ = _0450_ ? _1730_ : _1735_;
  assign _1737_ = _1736_ ^ _1725_;
  assign _1738_ = ~keysched_new_key_o[51];
  assign _1739_ = _1736_ ^ _1738_;
  assign _1740_ = _0479_ ? addroundkey_data_o[51] : _1739_;
  assign _1741_ = _0016_ ? addroundkey_data_o[51] : _1740_;
  assign next_addroundkey_data_reg[51] = _0004_ ? _1737_ : _1741_;
  assign _1742_ = ~key_i[52];
  assign _1743_ = ~subbytes_data_o[52];
  assign _1744_ = ~mixcol_data_o[52];
  assign _1745_ = ~data_i[52];
  assign _1746_ = _0459_ ? _1744_ : _1745_;
  assign _1747_ = _0455_ ? _1743_ : _1746_;
  assign _1748_ = _0470_ ? _1743_ : _1747_;
  assign _1749_ = _0469_ ? _1744_ : _1748_;
  assign _1750_ = subbytes_ready_o ? _1743_ : _1749_;
  assign _1751_ = _0468_ ? _1749_ : _1750_;
  assign _1752_ = _0463_ ? _1743_ : _1751_;
  assign _1753_ = _0450_ ? _1747_ : _1752_;
  assign _1754_ = _1753_ ^ _1742_;
  assign _1755_ = ~keysched_new_key_o[52];
  assign _1756_ = _1753_ ^ _1755_;
  assign _1757_ = _0479_ ? addroundkey_data_o[52] : _1756_;
  assign _1758_ = _0016_ ? addroundkey_data_o[52] : _1757_;
  assign next_addroundkey_data_reg[52] = _0004_ ? _1754_ : _1758_;
  assign _1759_ = ~key_i[53];
  assign _1760_ = ~subbytes_data_o[53];
  assign _1761_ = ~mixcol_data_o[53];
  assign _1762_ = ~data_i[53];
  assign _1763_ = _0459_ ? _1761_ : _1762_;
  assign _1764_ = _0455_ ? _1760_ : _1763_;
  assign _1765_ = _0470_ ? _1760_ : _1764_;
  assign _1766_ = _0469_ ? _1761_ : _1765_;
  assign _1767_ = subbytes_ready_o ? _1760_ : _1766_;
  assign _1768_ = _0468_ ? _1766_ : _1767_;
  assign _1769_ = _0463_ ? _1760_ : _1768_;
  assign _1770_ = _0450_ ? _1764_ : _1769_;
  assign _1771_ = _1770_ ^ _1759_;
  assign _1772_ = ~keysched_new_key_o[53];
  assign _1773_ = _1770_ ^ _1772_;
  assign _1774_ = _0479_ ? addroundkey_data_o[53] : _1773_;
  assign _1775_ = _0016_ ? addroundkey_data_o[53] : _1774_;
  assign next_addroundkey_data_reg[53] = _0004_ ? _1771_ : _1775_;
  assign _1776_ = ~key_i[54];
  assign _1777_ = ~subbytes_data_o[54];
  assign _1778_ = ~mixcol_data_o[54];
  assign _1779_ = ~data_i[54];
  assign _1780_ = _0459_ ? _1778_ : _1779_;
  assign _1781_ = _0455_ ? _1777_ : _1780_;
  assign _1782_ = _0470_ ? _1777_ : _1781_;
  assign _1783_ = _0469_ ? _1778_ : _1782_;
  assign _1784_ = subbytes_ready_o ? _1777_ : _1783_;
  assign _1785_ = _0468_ ? _1783_ : _1784_;
  assign _1786_ = _0463_ ? _1777_ : _1785_;
  assign _1787_ = _0450_ ? _1781_ : _1786_;
  assign _1788_ = _1787_ ^ _1776_;
  assign _1789_ = ~keysched_new_key_o[54];
  assign _1790_ = _1787_ ^ _1789_;
  assign _1791_ = _0479_ ? addroundkey_data_o[54] : _1790_;
  assign _1792_ = _0016_ ? addroundkey_data_o[54] : _1791_;
  assign next_addroundkey_data_reg[54] = _0004_ ? _1788_ : _1792_;
  assign _1793_ = ~key_i[55];
  assign _1794_ = ~subbytes_data_o[55];
  assign _1795_ = ~mixcol_data_o[55];
  assign _1796_ = ~data_i[55];
  assign _1797_ = _0459_ ? _1795_ : _1796_;
  assign _1798_ = _0455_ ? _1794_ : _1797_;
  assign _1799_ = _0470_ ? _1794_ : _1798_;
  assign _1800_ = _0469_ ? _1795_ : _1799_;
  assign _1801_ = subbytes_ready_o ? _1794_ : _1800_;
  assign _1802_ = _0468_ ? _1800_ : _1801_;
  assign _1803_ = _0463_ ? _1794_ : _1802_;
  assign _1804_ = _0450_ ? _1798_ : _1803_;
  assign _1805_ = _1804_ ^ _1793_;
  assign _1806_ = ~keysched_new_key_o[55];
  assign _1807_ = _1804_ ^ _1806_;
  assign _1808_ = _0479_ ? addroundkey_data_o[55] : _1807_;
  assign _1809_ = _0016_ ? addroundkey_data_o[55] : _1808_;
  assign next_addroundkey_data_reg[55] = _0004_ ? _1805_ : _1809_;
  assign _1810_ = ~key_i[56];
  assign _1811_ = ~subbytes_data_o[56];
  assign _1812_ = ~mixcol_data_o[56];
  assign _1813_ = ~data_i[56];
  assign _1814_ = _0459_ ? _1812_ : _1813_;
  assign _1815_ = _0455_ ? _1811_ : _1814_;
  assign _1816_ = _0470_ ? _1811_ : _1815_;
  assign _1817_ = _0469_ ? _1812_ : _1816_;
  assign _1818_ = subbytes_ready_o ? _1811_ : _1817_;
  assign _1819_ = _0468_ ? _1817_ : _1818_;
  assign _1820_ = _0463_ ? _1811_ : _1819_;
  assign _1821_ = _0450_ ? _1815_ : _1820_;
  assign _1822_ = _1821_ ^ _1810_;
  assign _1823_ = ~keysched_new_key_o[56];
  assign _1824_ = _1821_ ^ _1823_;
  assign _1825_ = _0479_ ? addroundkey_data_o[56] : _1824_;
  assign _1826_ = _0016_ ? addroundkey_data_o[56] : _1825_;
  assign next_addroundkey_data_reg[56] = _0004_ ? _1822_ : _1826_;
  assign _1827_ = ~key_i[57];
  assign _1828_ = ~subbytes_data_o[57];
  assign _1829_ = ~mixcol_data_o[57];
  assign _1830_ = ~data_i[57];
  assign _1831_ = _0459_ ? _1829_ : _1830_;
  assign _1832_ = _0455_ ? _1828_ : _1831_;
  assign _1833_ = _0470_ ? _1828_ : _1832_;
  assign _1834_ = _0469_ ? _1829_ : _1833_;
  assign _1835_ = subbytes_ready_o ? _1828_ : _1834_;
  assign _1836_ = _0468_ ? _1834_ : _1835_;
  assign _1837_ = _0463_ ? _1828_ : _1836_;
  assign _1838_ = _0450_ ? _1832_ : _1837_;
  assign _1839_ = _1838_ ^ _1827_;
  assign _1840_ = ~keysched_new_key_o[57];
  assign _1841_ = _1838_ ^ _1840_;
  assign _1842_ = _0479_ ? addroundkey_data_o[57] : _1841_;
  assign _1843_ = _0016_ ? addroundkey_data_o[57] : _1842_;
  assign next_addroundkey_data_reg[57] = _0004_ ? _1839_ : _1843_;
  assign _1844_ = ~key_i[58];
  assign _1845_ = ~subbytes_data_o[58];
  assign _1846_ = ~mixcol_data_o[58];
  assign _1847_ = ~data_i[58];
  assign _1848_ = _0459_ ? _1846_ : _1847_;
  assign _1849_ = _0455_ ? _1845_ : _1848_;
  assign _1850_ = _0470_ ? _1845_ : _1849_;
  assign _1851_ = _0469_ ? _1846_ : _1850_;
  assign _1852_ = subbytes_ready_o ? _1845_ : _1851_;
  assign _1853_ = _0468_ ? _1851_ : _1852_;
  assign _1854_ = _0463_ ? _1845_ : _1853_;
  assign _1855_ = _0450_ ? _1849_ : _1854_;
  assign _1856_ = _1855_ ^ _1844_;
  assign _1857_ = ~keysched_new_key_o[58];
  assign _1858_ = _1855_ ^ _1857_;
  assign _1859_ = _0479_ ? addroundkey_data_o[58] : _1858_;
  assign _1860_ = _0016_ ? addroundkey_data_o[58] : _1859_;
  assign next_addroundkey_data_reg[58] = _0004_ ? _1856_ : _1860_;
  assign _1861_ = ~key_i[59];
  assign _1862_ = ~subbytes_data_o[59];
  assign _1863_ = ~mixcol_data_o[59];
  assign _1864_ = ~data_i[59];
  assign _1865_ = _0459_ ? _1863_ : _1864_;
  assign _1866_ = _0455_ ? _1862_ : _1865_;
  assign _1867_ = _0470_ ? _1862_ : _1866_;
  assign _1868_ = _0469_ ? _1863_ : _1867_;
  assign _1869_ = subbytes_ready_o ? _1862_ : _1868_;
  assign _1870_ = _0468_ ? _1868_ : _1869_;
  assign _1871_ = _0463_ ? _1862_ : _1870_;
  assign _1872_ = _0450_ ? _1866_ : _1871_;
  assign _1873_ = _1872_ ^ _1861_;
  assign _1874_ = ~keysched_new_key_o[59];
  assign _1875_ = _1872_ ^ _1874_;
  assign _1876_ = _0479_ ? addroundkey_data_o[59] : _1875_;
  assign _1877_ = _0016_ ? addroundkey_data_o[59] : _1876_;
  assign next_addroundkey_data_reg[59] = _0004_ ? _1873_ : _1877_;
  assign _1878_ = ~key_i[5];
  assign _1879_ = ~subbytes_data_o[5];
  assign _1880_ = ~mixcol_data_o[5];
  assign _1881_ = ~data_i[5];
  assign _1882_ = _0459_ ? _1880_ : _1881_;
  assign _1883_ = _0455_ ? _1879_ : _1882_;
  assign _1884_ = _0470_ ? _1879_ : _1883_;
  assign _1885_ = _0469_ ? _1880_ : _1884_;
  assign _1886_ = subbytes_ready_o ? _1879_ : _1885_;
  assign _1887_ = _0468_ ? _1885_ : _1886_;
  assign _1888_ = _0463_ ? _1879_ : _1887_;
  assign _1889_ = _0450_ ? _1883_ : _1888_;
  assign _1890_ = _1889_ ^ _1878_;
  assign _1891_ = ~keysched_new_key_o[5];
  assign _1892_ = _1889_ ^ _1891_;
  assign _1893_ = _0479_ ? addroundkey_data_o[5] : _1892_;
  assign _1894_ = _0016_ ? addroundkey_data_o[5] : _1893_;
  assign next_addroundkey_data_reg[5] = _0004_ ? _1890_ : _1894_;
  assign _1895_ = ~key_i[60];
  assign _1896_ = ~subbytes_data_o[60];
  assign _1897_ = ~mixcol_data_o[60];
  assign _1898_ = ~data_i[60];
  assign _1899_ = _0459_ ? _1897_ : _1898_;
  assign _1900_ = _0455_ ? _1896_ : _1899_;
  assign _1901_ = _0470_ ? _1896_ : _1900_;
  assign _1902_ = _0469_ ? _1897_ : _1901_;
  assign _1903_ = subbytes_ready_o ? _1896_ : _1902_;
  assign _1904_ = _0468_ ? _1902_ : _1903_;
  assign _1905_ = _0463_ ? _1896_ : _1904_;
  assign _1906_ = _0450_ ? _1900_ : _1905_;
  assign _1907_ = _1906_ ^ _1895_;
  assign _1908_ = ~keysched_new_key_o[60];
  assign _1909_ = _1906_ ^ _1908_;
  assign _1910_ = _0479_ ? addroundkey_data_o[60] : _1909_;
  assign _1911_ = _0016_ ? addroundkey_data_o[60] : _1910_;
  assign next_addroundkey_data_reg[60] = _0004_ ? _1907_ : _1911_;
  assign _1912_ = ~key_i[61];
  assign _1913_ = ~subbytes_data_o[61];
  assign _1914_ = ~mixcol_data_o[61];
  assign _1915_ = ~data_i[61];
  assign _1916_ = _0459_ ? _1914_ : _1915_;
  assign _1917_ = _0455_ ? _1913_ : _1916_;
  assign _1918_ = _0470_ ? _1913_ : _1917_;
  assign _1919_ = _0469_ ? _1914_ : _1918_;
  assign _1920_ = subbytes_ready_o ? _1913_ : _1919_;
  assign _1921_ = _0468_ ? _1919_ : _1920_;
  assign _1922_ = _0463_ ? _1913_ : _1921_;
  assign _1923_ = _0450_ ? _1917_ : _1922_;
  assign _1924_ = _1923_ ^ _1912_;
  assign _1925_ = ~keysched_new_key_o[61];
  assign _1926_ = _1923_ ^ _1925_;
  assign _1927_ = _0479_ ? addroundkey_data_o[61] : _1926_;
  assign _1928_ = _0016_ ? addroundkey_data_o[61] : _1927_;
  assign next_addroundkey_data_reg[61] = _0004_ ? _1924_ : _1928_;
  assign _1929_ = ~key_i[62];
  assign _1930_ = ~subbytes_data_o[62];
  assign _1931_ = ~mixcol_data_o[62];
  assign _1932_ = ~data_i[62];
  assign _1933_ = _0459_ ? _1931_ : _1932_;
  assign _1934_ = _0455_ ? _1930_ : _1933_;
  assign _1935_ = _0470_ ? _1930_ : _1934_;
  assign _1936_ = _0469_ ? _1931_ : _1935_;
  assign _1937_ = subbytes_ready_o ? _1930_ : _1936_;
  assign _1938_ = _0468_ ? _1936_ : _1937_;
  assign _1939_ = _0463_ ? _1930_ : _1938_;
  assign _1940_ = _0450_ ? _1934_ : _1939_;
  assign _1941_ = _1940_ ^ _1929_;
  assign _1942_ = ~keysched_new_key_o[62];
  assign _1943_ = _1940_ ^ _1942_;
  assign _1944_ = _0479_ ? addroundkey_data_o[62] : _1943_;
  assign _1945_ = _0016_ ? addroundkey_data_o[62] : _1944_;
  assign next_addroundkey_data_reg[62] = _0004_ ? _1941_ : _1945_;
  assign _1946_ = ~key_i[63];
  assign _1947_ = ~subbytes_data_o[63];
  assign _1948_ = ~mixcol_data_o[63];
  assign _1949_ = ~data_i[63];
  assign _1950_ = _0459_ ? _1948_ : _1949_;
  assign _1951_ = _0455_ ? _1947_ : _1950_;
  assign _1952_ = _0470_ ? _1947_ : _1951_;
  assign _1953_ = _0469_ ? _1948_ : _1952_;
  assign _1954_ = subbytes_ready_o ? _1947_ : _1953_;
  assign _1955_ = _0468_ ? _1953_ : _1954_;
  assign _1956_ = _0463_ ? _1947_ : _1955_;
  assign _1957_ = _0450_ ? _1951_ : _1956_;
  assign _1958_ = _1957_ ^ _1946_;
  assign _1959_ = ~keysched_new_key_o[63];
  assign _1960_ = _1957_ ^ _1959_;
  assign _1961_ = _0479_ ? addroundkey_data_o[63] : _1960_;
  assign _1962_ = _0016_ ? addroundkey_data_o[63] : _1961_;
  assign next_addroundkey_data_reg[63] = _0004_ ? _1958_ : _1962_;
  assign _1963_ = ~key_i[64];
  assign _1964_ = ~subbytes_data_o[64];
  assign _1965_ = ~mixcol_data_o[64];
  assign _1966_ = ~data_i[64];
  assign _1967_ = _0459_ ? _1965_ : _1966_;
  assign _1968_ = _0455_ ? _1964_ : _1967_;
  assign _1969_ = _0470_ ? _1964_ : _1968_;
  assign _1970_ = _0469_ ? _1965_ : _1969_;
  assign _1971_ = subbytes_ready_o ? _1964_ : _1970_;
  assign _1972_ = _0468_ ? _1970_ : _1971_;
  assign _1973_ = _0463_ ? _1964_ : _1972_;
  assign _1974_ = _0450_ ? _1968_ : _1973_;
  assign _1975_ = _1974_ ^ _1963_;
  assign _1976_ = ~keysched_new_key_o[64];
  assign _1977_ = _1974_ ^ _1976_;
  assign _1978_ = _0479_ ? addroundkey_data_o[64] : _1977_;
  assign _1979_ = _0016_ ? addroundkey_data_o[64] : _1978_;
  assign next_addroundkey_data_reg[64] = _0004_ ? _1975_ : _1979_;
  assign _1980_ = ~key_i[65];
  assign _1981_ = ~subbytes_data_o[65];
  assign _1982_ = ~mixcol_data_o[65];
  assign _1983_ = ~data_i[65];
  assign _1984_ = _0459_ ? _1982_ : _1983_;
  assign _1985_ = _0455_ ? _1981_ : _1984_;
  assign _1986_ = _0470_ ? _1981_ : _1985_;
  assign _1987_ = _0469_ ? _1982_ : _1986_;
  assign _1988_ = subbytes_ready_o ? _1981_ : _1987_;
  assign _1989_ = _0468_ ? _1987_ : _1988_;
  assign _1990_ = _0463_ ? _1981_ : _1989_;
  assign _1991_ = _0450_ ? _1985_ : _1990_;
  assign _1992_ = _1991_ ^ _1980_;
  assign _1993_ = ~keysched_new_key_o[65];
  assign _1994_ = _1991_ ^ _1993_;
  assign _1995_ = _0479_ ? addroundkey_data_o[65] : _1994_;
  assign _1996_ = _0016_ ? addroundkey_data_o[65] : _1995_;
  assign next_addroundkey_data_reg[65] = _0004_ ? _1992_ : _1996_;
  assign _1997_ = ~key_i[66];
  assign _1998_ = ~subbytes_data_o[66];
  assign _1999_ = ~mixcol_data_o[66];
  assign _2000_ = ~data_i[66];
  assign _2001_ = _0459_ ? _1999_ : _2000_;
  assign _2002_ = _0455_ ? _1998_ : _2001_;
  assign _2003_ = _0470_ ? _1998_ : _2002_;
  assign _2004_ = _0469_ ? _1999_ : _2003_;
  assign _2005_ = subbytes_ready_o ? _1998_ : _2004_;
  assign _2006_ = _0468_ ? _2004_ : _2005_;
  assign _2007_ = _0463_ ? _1998_ : _2006_;
  assign _2008_ = _0450_ ? _2002_ : _2007_;
  assign _2009_ = _2008_ ^ _1997_;
  assign _2010_ = ~keysched_new_key_o[66];
  assign _2011_ = _2008_ ^ _2010_;
  assign _2012_ = _0479_ ? addroundkey_data_o[66] : _2011_;
  assign _2013_ = _0016_ ? addroundkey_data_o[66] : _2012_;
  assign next_addroundkey_data_reg[66] = _0004_ ? _2009_ : _2013_;
  assign _2014_ = ~key_i[67];
  assign _2015_ = ~subbytes_data_o[67];
  assign _2016_ = ~mixcol_data_o[67];
  assign _2017_ = ~data_i[67];
  assign _2018_ = _0459_ ? _2016_ : _2017_;
  assign _2019_ = _0455_ ? _2015_ : _2018_;
  assign _2020_ = _0470_ ? _2015_ : _2019_;
  assign _2021_ = _0469_ ? _2016_ : _2020_;
  assign _2022_ = subbytes_ready_o ? _2015_ : _2021_;
  assign _2023_ = _0468_ ? _2021_ : _2022_;
  assign _2024_ = _0463_ ? _2015_ : _2023_;
  assign _2025_ = _0450_ ? _2019_ : _2024_;
  assign _2026_ = _2025_ ^ _2014_;
  assign _2027_ = ~keysched_new_key_o[67];
  assign _2028_ = _2025_ ^ _2027_;
  assign _2029_ = _0479_ ? addroundkey_data_o[67] : _2028_;
  assign _2030_ = _0016_ ? addroundkey_data_o[67] : _2029_;
  assign next_addroundkey_data_reg[67] = _0004_ ? _2026_ : _2030_;
  assign _2031_ = ~key_i[68];
  assign _2032_ = ~subbytes_data_o[68];
  assign _2033_ = ~mixcol_data_o[68];
  assign _2034_ = ~data_i[68];
  assign _2035_ = _0459_ ? _2033_ : _2034_;
  assign _2036_ = _0455_ ? _2032_ : _2035_;
  assign _2037_ = _0470_ ? _2032_ : _2036_;
  assign _2038_ = _0469_ ? _2033_ : _2037_;
  assign _2039_ = subbytes_ready_o ? _2032_ : _2038_;
  assign _2040_ = _0468_ ? _2038_ : _2039_;
  assign _2041_ = _0463_ ? _2032_ : _2040_;
  assign _2042_ = _0450_ ? _2036_ : _2041_;
  assign _2043_ = _2042_ ^ _2031_;
  assign _2044_ = ~keysched_new_key_o[68];
  assign _2045_ = _2042_ ^ _2044_;
  assign _2046_ = _0479_ ? addroundkey_data_o[68] : _2045_;
  assign _2047_ = _0016_ ? addroundkey_data_o[68] : _2046_;
  assign next_addroundkey_data_reg[68] = _0004_ ? _2043_ : _2047_;
  assign _2048_ = ~key_i[69];
  assign _2049_ = ~subbytes_data_o[69];
  assign _2050_ = ~mixcol_data_o[69];
  assign _2051_ = ~data_i[69];
  assign _2052_ = _0459_ ? _2050_ : _2051_;
  assign _2053_ = _0455_ ? _2049_ : _2052_;
  assign _2054_ = _0470_ ? _2049_ : _2053_;
  assign _2055_ = _0469_ ? _2050_ : _2054_;
  assign _2056_ = subbytes_ready_o ? _2049_ : _2055_;
  assign _2057_ = _0468_ ? _2055_ : _2056_;
  assign _2058_ = _0463_ ? _2049_ : _2057_;
  assign _2059_ = _0450_ ? _2053_ : _2058_;
  assign _2060_ = _2059_ ^ _2048_;
  assign _2061_ = ~keysched_new_key_o[69];
  assign _2062_ = _2059_ ^ _2061_;
  assign _2063_ = _0479_ ? addroundkey_data_o[69] : _2062_;
  assign _2064_ = _0016_ ? addroundkey_data_o[69] : _2063_;
  assign next_addroundkey_data_reg[69] = _0004_ ? _2060_ : _2064_;
  assign _2065_ = ~key_i[6];
  assign _2066_ = ~subbytes_data_o[6];
  assign _2067_ = ~mixcol_data_o[6];
  assign _2068_ = ~data_i[6];
  assign _2069_ = _0459_ ? _2067_ : _2068_;
  assign _2070_ = _0455_ ? _2066_ : _2069_;
  assign _2071_ = _0470_ ? _2066_ : _2070_;
  assign _2072_ = _0469_ ? _2067_ : _2071_;
  assign _2073_ = subbytes_ready_o ? _2066_ : _2072_;
  assign _2074_ = _0468_ ? _2072_ : _2073_;
  assign _2075_ = _0463_ ? _2066_ : _2074_;
  assign _2076_ = _0450_ ? _2070_ : _2075_;
  assign _2077_ = _2076_ ^ _2065_;
  assign _2078_ = ~keysched_new_key_o[6];
  assign _2079_ = _2076_ ^ _2078_;
  assign _2080_ = _0479_ ? addroundkey_data_o[6] : _2079_;
  assign _2081_ = _0016_ ? addroundkey_data_o[6] : _2080_;
  assign next_addroundkey_data_reg[6] = _0004_ ? _2077_ : _2081_;
  assign _2082_ = ~key_i[70];
  assign _2083_ = ~subbytes_data_o[70];
  assign _2084_ = ~mixcol_data_o[70];
  assign _2085_ = ~data_i[70];
  assign _2086_ = _0459_ ? _2084_ : _2085_;
  assign _2087_ = _0455_ ? _2083_ : _2086_;
  assign _2088_ = _0470_ ? _2083_ : _2087_;
  assign _2089_ = _0469_ ? _2084_ : _2088_;
  assign _2090_ = subbytes_ready_o ? _2083_ : _2089_;
  assign _2091_ = _0468_ ? _2089_ : _2090_;
  assign _2092_ = _0463_ ? _2083_ : _2091_;
  assign _2093_ = _0450_ ? _2087_ : _2092_;
  assign _2094_ = _2093_ ^ _2082_;
  assign _2095_ = ~keysched_new_key_o[70];
  assign _2096_ = _2093_ ^ _2095_;
  assign _2097_ = _0479_ ? addroundkey_data_o[70] : _2096_;
  assign _2098_ = _0016_ ? addroundkey_data_o[70] : _2097_;
  assign next_addroundkey_data_reg[70] = _0004_ ? _2094_ : _2098_;
  assign _2099_ = ~key_i[71];
  assign _2100_ = ~subbytes_data_o[71];
  assign _2101_ = ~mixcol_data_o[71];
  assign _2102_ = ~data_i[71];
  assign _2103_ = _0459_ ? _2101_ : _2102_;
  assign _2104_ = _0455_ ? _2100_ : _2103_;
  assign _2105_ = _0470_ ? _2100_ : _2104_;
  assign _2106_ = _0469_ ? _2101_ : _2105_;
  assign _2107_ = subbytes_ready_o ? _2100_ : _2106_;
  assign _2108_ = _0468_ ? _2106_ : _2107_;
  assign _2109_ = _0463_ ? _2100_ : _2108_;
  assign _2110_ = _0450_ ? _2104_ : _2109_;
  assign _2111_ = _2110_ ^ _2099_;
  assign _2112_ = ~keysched_new_key_o[71];
  assign _2113_ = _2110_ ^ _2112_;
  assign _2114_ = _0479_ ? addroundkey_data_o[71] : _2113_;
  assign _2115_ = _0016_ ? addroundkey_data_o[71] : _2114_;
  assign next_addroundkey_data_reg[71] = _0004_ ? _2111_ : _2115_;
  assign _2116_ = ~key_i[72];
  assign _2117_ = ~subbytes_data_o[72];
  assign _2118_ = ~mixcol_data_o[72];
  assign _2119_ = ~data_i[72];
  assign _2120_ = _0459_ ? _2118_ : _2119_;
  assign _2121_ = _0455_ ? _2117_ : _2120_;
  assign _2122_ = _0470_ ? _2117_ : _2121_;
  assign _2123_ = _0469_ ? _2118_ : _2122_;
  assign _2124_ = subbytes_ready_o ? _2117_ : _2123_;
  assign _2125_ = _0468_ ? _2123_ : _2124_;
  assign _2126_ = _0463_ ? _2117_ : _2125_;
  assign _2127_ = _0450_ ? _2121_ : _2126_;
  assign _2128_ = _2127_ ^ _2116_;
  assign _2129_ = ~keysched_new_key_o[72];
  assign _2130_ = _2127_ ^ _2129_;
  assign _2131_ = _0479_ ? addroundkey_data_o[72] : _2130_;
  assign _2132_ = _0016_ ? addroundkey_data_o[72] : _2131_;
  assign next_addroundkey_data_reg[72] = _0004_ ? _2128_ : _2132_;
  assign _2133_ = ~key_i[73];
  assign _2134_ = ~subbytes_data_o[73];
  assign _2135_ = ~mixcol_data_o[73];
  assign _2136_ = ~data_i[73];
  assign _2137_ = _0459_ ? _2135_ : _2136_;
  assign _2138_ = _0455_ ? _2134_ : _2137_;
  assign _2139_ = _0470_ ? _2134_ : _2138_;
  assign _2140_ = _0469_ ? _2135_ : _2139_;
  assign _2141_ = subbytes_ready_o ? _2134_ : _2140_;
  assign _2142_ = _0468_ ? _2140_ : _2141_;
  assign _2143_ = _0463_ ? _2134_ : _2142_;
  assign _2144_ = _0450_ ? _2138_ : _2143_;
  assign _2145_ = _2144_ ^ _2133_;
  assign _2146_ = ~keysched_new_key_o[73];
  assign _2147_ = _2144_ ^ _2146_;
  assign _2148_ = _0479_ ? addroundkey_data_o[73] : _2147_;
  assign _2149_ = _0016_ ? addroundkey_data_o[73] : _2148_;
  assign next_addroundkey_data_reg[73] = _0004_ ? _2145_ : _2149_;
  assign _2150_ = ~key_i[74];
  assign _2151_ = ~subbytes_data_o[74];
  assign _2152_ = ~mixcol_data_o[74];
  assign _2153_ = ~data_i[74];
  assign _2154_ = _0459_ ? _2152_ : _2153_;
  assign _2155_ = _0455_ ? _2151_ : _2154_;
  assign _2156_ = _0470_ ? _2151_ : _2155_;
  assign _2157_ = _0469_ ? _2152_ : _2156_;
  assign _2158_ = subbytes_ready_o ? _2151_ : _2157_;
  assign _2159_ = _0468_ ? _2157_ : _2158_;
  assign _2160_ = _0463_ ? _2151_ : _2159_;
  assign _2161_ = _0450_ ? _2155_ : _2160_;
  assign _2162_ = _2161_ ^ _2150_;
  assign _2163_ = ~keysched_new_key_o[74];
  assign _2164_ = _2161_ ^ _2163_;
  assign _2165_ = _0479_ ? addroundkey_data_o[74] : _2164_;
  assign _2166_ = _0016_ ? addroundkey_data_o[74] : _2165_;
  assign next_addroundkey_data_reg[74] = _0004_ ? _2162_ : _2166_;
  assign _2167_ = ~key_i[75];
  assign _2168_ = ~subbytes_data_o[75];
  assign _2169_ = ~mixcol_data_o[75];
  assign _2170_ = ~data_i[75];
  assign _2171_ = _0459_ ? _2169_ : _2170_;
  assign _2172_ = _0455_ ? _2168_ : _2171_;
  assign _2173_ = _0470_ ? _2168_ : _2172_;
  assign _2174_ = _0469_ ? _2169_ : _2173_;
  assign _2175_ = subbytes_ready_o ? _2168_ : _2174_;
  assign _2176_ = _0468_ ? _2174_ : _2175_;
  assign _2177_ = _0463_ ? _2168_ : _2176_;
  assign _2178_ = _0450_ ? _2172_ : _2177_;
  assign _2179_ = _2178_ ^ _2167_;
  assign _2180_ = ~keysched_new_key_o[75];
  assign _2181_ = _2178_ ^ _2180_;
  assign _2182_ = _0479_ ? addroundkey_data_o[75] : _2181_;
  assign _2183_ = _0016_ ? addroundkey_data_o[75] : _2182_;
  assign next_addroundkey_data_reg[75] = _0004_ ? _2179_ : _2183_;
  assign _2184_ = ~key_i[76];
  assign _2185_ = ~subbytes_data_o[76];
  assign _2186_ = ~mixcol_data_o[76];
  assign _2187_ = ~data_i[76];
  assign _2188_ = _0459_ ? _2186_ : _2187_;
  assign _2189_ = _0455_ ? _2185_ : _2188_;
  assign _2190_ = _0470_ ? _2185_ : _2189_;
  assign _2191_ = _0469_ ? _2186_ : _2190_;
  assign _2192_ = subbytes_ready_o ? _2185_ : _2191_;
  assign _2193_ = _0468_ ? _2191_ : _2192_;
  assign _2194_ = _0463_ ? _2185_ : _2193_;
  assign _2195_ = _0450_ ? _2189_ : _2194_;
  assign _2196_ = _2195_ ^ _2184_;
  assign _2197_ = ~keysched_new_key_o[76];
  assign _2198_ = _2195_ ^ _2197_;
  assign _2199_ = _0479_ ? addroundkey_data_o[76] : _2198_;
  assign _2200_ = _0016_ ? addroundkey_data_o[76] : _2199_;
  assign next_addroundkey_data_reg[76] = _0004_ ? _2196_ : _2200_;
  assign _2201_ = ~key_i[77];
  assign _2202_ = ~subbytes_data_o[77];
  assign _2203_ = ~mixcol_data_o[77];
  assign _2204_ = ~data_i[77];
  assign _2205_ = _0459_ ? _2203_ : _2204_;
  assign _2206_ = _0455_ ? _2202_ : _2205_;
  assign _2207_ = _0470_ ? _2202_ : _2206_;
  assign _2208_ = _0469_ ? _2203_ : _2207_;
  assign _2209_ = subbytes_ready_o ? _2202_ : _2208_;
  assign _2210_ = _0468_ ? _2208_ : _2209_;
  assign _2211_ = _0463_ ? _2202_ : _2210_;
  assign _2212_ = _0450_ ? _2206_ : _2211_;
  assign _2213_ = _2212_ ^ _2201_;
  assign _2214_ = ~keysched_new_key_o[77];
  assign _2215_ = _2212_ ^ _2214_;
  assign _2216_ = _0479_ ? addroundkey_data_o[77] : _2215_;
  assign _2217_ = _0016_ ? addroundkey_data_o[77] : _2216_;
  assign next_addroundkey_data_reg[77] = _0004_ ? _2213_ : _2217_;
  assign _2218_ = ~key_i[78];
  assign _2219_ = ~subbytes_data_o[78];
  assign _2220_ = ~mixcol_data_o[78];
  assign _2221_ = ~data_i[78];
  assign _2222_ = _0459_ ? _2220_ : _2221_;
  assign _2223_ = _0455_ ? _2219_ : _2222_;
  assign _2224_ = _0470_ ? _2219_ : _2223_;
  assign _2225_ = _0469_ ? _2220_ : _2224_;
  assign _2226_ = subbytes_ready_o ? _2219_ : _2225_;
  assign _2227_ = _0468_ ? _2225_ : _2226_;
  assign _2228_ = _0463_ ? _2219_ : _2227_;
  assign _2229_ = _0450_ ? _2223_ : _2228_;
  assign _2230_ = _2229_ ^ _2218_;
  assign _2231_ = ~keysched_new_key_o[78];
  assign _2232_ = _2229_ ^ _2231_;
  assign _2233_ = _0479_ ? addroundkey_data_o[78] : _2232_;
  assign _2234_ = _0016_ ? addroundkey_data_o[78] : _2233_;
  assign next_addroundkey_data_reg[78] = _0004_ ? _2230_ : _2234_;
  assign _2235_ = ~key_i[79];
  assign _2236_ = ~subbytes_data_o[79];
  assign _2237_ = ~mixcol_data_o[79];
  assign _2238_ = ~data_i[79];
  assign _2239_ = _0459_ ? _2237_ : _2238_;
  assign _2240_ = _0455_ ? _2236_ : _2239_;
  assign _2241_ = _0470_ ? _2236_ : _2240_;
  assign _2242_ = _0469_ ? _2237_ : _2241_;
  assign _2243_ = subbytes_ready_o ? _2236_ : _2242_;
  assign _2244_ = _0468_ ? _2242_ : _2243_;
  assign _2245_ = _0463_ ? _2236_ : _2244_;
  assign _2246_ = _0450_ ? _2240_ : _2245_;
  assign _2247_ = _2246_ ^ _2235_;
  assign _2248_ = ~keysched_new_key_o[79];
  assign _2249_ = _2246_ ^ _2248_;
  assign _2250_ = _0479_ ? addroundkey_data_o[79] : _2249_;
  assign _2251_ = _0016_ ? addroundkey_data_o[79] : _2250_;
  assign next_addroundkey_data_reg[79] = _0004_ ? _2247_ : _2251_;
  assign _2252_ = ~key_i[7];
  assign _2253_ = ~subbytes_data_o[7];
  assign _2254_ = ~mixcol_data_o[7];
  assign _2255_ = ~data_i[7];
  assign _2256_ = _0459_ ? _2254_ : _2255_;
  assign _2257_ = _0455_ ? _2253_ : _2256_;
  assign _2258_ = _0470_ ? _2253_ : _2257_;
  assign _2259_ = _0469_ ? _2254_ : _2258_;
  assign _2260_ = subbytes_ready_o ? _2253_ : _2259_;
  assign _2261_ = _0468_ ? _2259_ : _2260_;
  assign _2262_ = _0463_ ? _2253_ : _2261_;
  assign _2263_ = _0450_ ? _2257_ : _2262_;
  assign _2264_ = _2263_ ^ _2252_;
  assign _2265_ = ~keysched_new_key_o[7];
  assign _2266_ = _2263_ ^ _2265_;
  assign _2267_ = _0479_ ? addroundkey_data_o[7] : _2266_;
  assign _2268_ = _0016_ ? addroundkey_data_o[7] : _2267_;
  assign next_addroundkey_data_reg[7] = _0004_ ? _2264_ : _2268_;
  assign _2269_ = ~key_i[80];
  assign _2270_ = ~subbytes_data_o[80];
  assign _2271_ = ~mixcol_data_o[80];
  assign _2272_ = ~data_i[80];
  assign _2273_ = _0459_ ? _2271_ : _2272_;
  assign _2274_ = _0455_ ? _2270_ : _2273_;
  assign _2275_ = _0470_ ? _2270_ : _2274_;
  assign _2276_ = _0469_ ? _2271_ : _2275_;
  assign _2277_ = subbytes_ready_o ? _2270_ : _2276_;
  assign _2278_ = _0468_ ? _2276_ : _2277_;
  assign _2279_ = _0463_ ? _2270_ : _2278_;
  assign _2280_ = _0450_ ? _2274_ : _2279_;
  assign _2281_ = _2280_ ^ _2269_;
  assign _2282_ = ~keysched_new_key_o[80];
  assign _2283_ = _2280_ ^ _2282_;
  assign _2284_ = _0479_ ? addroundkey_data_o[80] : _2283_;
  assign _2285_ = _0016_ ? addroundkey_data_o[80] : _2284_;
  assign next_addroundkey_data_reg[80] = _0004_ ? _2281_ : _2285_;
  assign _2286_ = ~key_i[81];
  assign _2287_ = ~subbytes_data_o[81];
  assign _2288_ = ~mixcol_data_o[81];
  assign _2289_ = ~data_i[81];
  assign _2290_ = _0459_ ? _2288_ : _2289_;
  assign _2291_ = _0455_ ? _2287_ : _2290_;
  assign _2292_ = _0470_ ? _2287_ : _2291_;
  assign _2293_ = _0469_ ? _2288_ : _2292_;
  assign _2294_ = subbytes_ready_o ? _2287_ : _2293_;
  assign _2295_ = _0468_ ? _2293_ : _2294_;
  assign _2296_ = _0463_ ? _2287_ : _2295_;
  assign _2297_ = _0450_ ? _2291_ : _2296_;
  assign _2298_ = _2297_ ^ _2286_;
  assign _2299_ = ~keysched_new_key_o[81];
  assign _2300_ = _2297_ ^ _2299_;
  assign _2301_ = _0479_ ? addroundkey_data_o[81] : _2300_;
  assign _2302_ = _0016_ ? addroundkey_data_o[81] : _2301_;
  assign next_addroundkey_data_reg[81] = _0004_ ? _2298_ : _2302_;
  assign _2303_ = ~key_i[82];
  assign _2304_ = ~subbytes_data_o[82];
  assign _2305_ = ~mixcol_data_o[82];
  assign _2306_ = ~data_i[82];
  assign _2307_ = _0459_ ? _2305_ : _2306_;
  assign _2308_ = _0455_ ? _2304_ : _2307_;
  assign _2309_ = _0470_ ? _2304_ : _2308_;
  assign _2310_ = _0469_ ? _2305_ : _2309_;
  assign _2311_ = subbytes_ready_o ? _2304_ : _2310_;
  assign _2312_ = _0468_ ? _2310_ : _2311_;
  assign _2313_ = _0463_ ? _2304_ : _2312_;
  assign _2314_ = _0450_ ? _2308_ : _2313_;
  assign _2315_ = _2314_ ^ _2303_;
  assign _2316_ = ~keysched_new_key_o[82];
  assign _2317_ = _2314_ ^ _2316_;
  assign _2318_ = _0479_ ? addroundkey_data_o[82] : _2317_;
  assign _2319_ = _0016_ ? addroundkey_data_o[82] : _2318_;
  assign next_addroundkey_data_reg[82] = _0004_ ? _2315_ : _2319_;
  assign _2320_ = ~key_i[83];
  assign _2321_ = ~subbytes_data_o[83];
  assign _2322_ = ~mixcol_data_o[83];
  assign _2323_ = ~data_i[83];
  assign _2324_ = _0459_ ? _2322_ : _2323_;
  assign _2325_ = _0455_ ? _2321_ : _2324_;
  assign _2326_ = _0470_ ? _2321_ : _2325_;
  assign _2327_ = _0469_ ? _2322_ : _2326_;
  assign _2328_ = subbytes_ready_o ? _2321_ : _2327_;
  assign _2329_ = _0468_ ? _2327_ : _2328_;
  assign _2330_ = _0463_ ? _2321_ : _2329_;
  assign _2331_ = _0450_ ? _2325_ : _2330_;
  assign _2332_ = _2331_ ^ _2320_;
  assign _2333_ = ~keysched_new_key_o[83];
  assign _2334_ = _2331_ ^ _2333_;
  assign _2335_ = _0479_ ? addroundkey_data_o[83] : _2334_;
  assign _2336_ = _0016_ ? addroundkey_data_o[83] : _2335_;
  assign next_addroundkey_data_reg[83] = _0004_ ? _2332_ : _2336_;
  assign _2337_ = ~key_i[84];
  assign _2338_ = ~subbytes_data_o[84];
  assign _2339_ = ~mixcol_data_o[84];
  assign _2340_ = ~data_i[84];
  assign _2341_ = _0459_ ? _2339_ : _2340_;
  assign _2342_ = _0455_ ? _2338_ : _2341_;
  assign _2343_ = _0470_ ? _2338_ : _2342_;
  assign _2344_ = _0469_ ? _2339_ : _2343_;
  assign _2345_ = subbytes_ready_o ? _2338_ : _2344_;
  assign _2346_ = _0468_ ? _2344_ : _2345_;
  assign _2347_ = _0463_ ? _2338_ : _2346_;
  assign _2348_ = _0450_ ? _2342_ : _2347_;
  assign _2349_ = _2348_ ^ _2337_;
  assign _2350_ = ~keysched_new_key_o[84];
  assign _2351_ = _2348_ ^ _2350_;
  assign _2352_ = _0479_ ? addroundkey_data_o[84] : _2351_;
  assign _2353_ = _0016_ ? addroundkey_data_o[84] : _2352_;
  assign next_addroundkey_data_reg[84] = _0004_ ? _2349_ : _2353_;
  assign _2354_ = ~key_i[85];
  assign _2355_ = ~subbytes_data_o[85];
  assign _2356_ = ~mixcol_data_o[85];
  assign _2357_ = ~data_i[85];
  assign _2358_ = _0459_ ? _2356_ : _2357_;
  assign _2359_ = _0455_ ? _2355_ : _2358_;
  assign _2360_ = _0470_ ? _2355_ : _2359_;
  assign _2361_ = _0469_ ? _2356_ : _2360_;
  assign _2362_ = subbytes_ready_o ? _2355_ : _2361_;
  assign _2363_ = _0468_ ? _2361_ : _2362_;
  assign _2364_ = _0463_ ? _2355_ : _2363_;
  assign _2365_ = _0450_ ? _2359_ : _2364_;
  assign _2366_ = _2365_ ^ _2354_;
  assign _2367_ = ~keysched_new_key_o[85];
  assign _2368_ = _2365_ ^ _2367_;
  assign _2369_ = _0479_ ? addroundkey_data_o[85] : _2368_;
  assign _2370_ = _0016_ ? addroundkey_data_o[85] : _2369_;
  assign next_addroundkey_data_reg[85] = _0004_ ? _2366_ : _2370_;
  assign _2371_ = ~key_i[86];
  assign _2372_ = ~subbytes_data_o[86];
  assign _2373_ = ~mixcol_data_o[86];
  assign _2374_ = ~data_i[86];
  assign _2375_ = _0459_ ? _2373_ : _2374_;
  assign _2376_ = _0455_ ? _2372_ : _2375_;
  assign _2377_ = _0470_ ? _2372_ : _2376_;
  assign _2378_ = _0469_ ? _2373_ : _2377_;
  assign _2379_ = subbytes_ready_o ? _2372_ : _2378_;
  assign _2380_ = _0468_ ? _2378_ : _2379_;
  assign _2381_ = _0463_ ? _2372_ : _2380_;
  assign _2382_ = _0450_ ? _2376_ : _2381_;
  assign _2383_ = _2382_ ^ _2371_;
  assign _2384_ = ~keysched_new_key_o[86];
  assign _2385_ = _2382_ ^ _2384_;
  assign _2386_ = _0479_ ? addroundkey_data_o[86] : _2385_;
  assign _2387_ = _0016_ ? addroundkey_data_o[86] : _2386_;
  assign next_addroundkey_data_reg[86] = _0004_ ? _2383_ : _2387_;
  assign _2388_ = ~key_i[87];
  assign _2389_ = ~subbytes_data_o[87];
  assign _2390_ = ~mixcol_data_o[87];
  assign _2391_ = ~data_i[87];
  assign _2392_ = _0459_ ? _2390_ : _2391_;
  assign _2393_ = _0455_ ? _2389_ : _2392_;
  assign _2394_ = _0470_ ? _2389_ : _2393_;
  assign _2395_ = _0469_ ? _2390_ : _2394_;
  assign _2396_ = subbytes_ready_o ? _2389_ : _2395_;
  assign _2397_ = _0468_ ? _2395_ : _2396_;
  assign _2398_ = _0463_ ? _2389_ : _2397_;
  assign _2399_ = _0450_ ? _2393_ : _2398_;
  assign _2400_ = _2399_ ^ _2388_;
  assign _2401_ = ~keysched_new_key_o[87];
  assign _2402_ = _2399_ ^ _2401_;
  assign _2403_ = _0479_ ? addroundkey_data_o[87] : _2402_;
  assign _2404_ = _0016_ ? addroundkey_data_o[87] : _2403_;
  assign next_addroundkey_data_reg[87] = _0004_ ? _2400_ : _2404_;
  assign _2405_ = ~key_i[88];
  assign _2406_ = ~subbytes_data_o[88];
  assign _2407_ = ~mixcol_data_o[88];
  assign _2408_ = ~data_i[88];
  assign _2409_ = _0459_ ? _2407_ : _2408_;
  assign _2410_ = _0455_ ? _2406_ : _2409_;
  assign _2411_ = _0470_ ? _2406_ : _2410_;
  assign _2412_ = _0469_ ? _2407_ : _2411_;
  assign _2413_ = subbytes_ready_o ? _2406_ : _2412_;
  assign _2414_ = _0468_ ? _2412_ : _2413_;
  assign _2415_ = _0463_ ? _2406_ : _2414_;
  assign _2416_ = _0450_ ? _2410_ : _2415_;
  assign _2417_ = _2416_ ^ _2405_;
  assign _2418_ = ~keysched_new_key_o[88];
  assign _2419_ = _2416_ ^ _2418_;
  assign _2420_ = _0479_ ? addroundkey_data_o[88] : _2419_;
  assign _2421_ = _0016_ ? addroundkey_data_o[88] : _2420_;
  assign next_addroundkey_data_reg[88] = _0004_ ? _2417_ : _2421_;
  assign _2422_ = ~key_i[89];
  assign _2423_ = ~subbytes_data_o[89];
  assign _2424_ = ~mixcol_data_o[89];
  assign _2425_ = ~data_i[89];
  assign _2426_ = _0459_ ? _2424_ : _2425_;
  assign _2427_ = _0455_ ? _2423_ : _2426_;
  assign _2428_ = _0470_ ? _2423_ : _2427_;
  assign _2429_ = _0469_ ? _2424_ : _2428_;
  assign _2430_ = subbytes_ready_o ? _2423_ : _2429_;
  assign _2431_ = _0468_ ? _2429_ : _2430_;
  assign _2432_ = _0463_ ? _2423_ : _2431_;
  assign _2433_ = _0450_ ? _2427_ : _2432_;
  assign _2434_ = _2433_ ^ _2422_;
  assign _2435_ = ~keysched_new_key_o[89];
  assign _2436_ = _2433_ ^ _2435_;
  assign _2437_ = _0479_ ? addroundkey_data_o[89] : _2436_;
  assign _2438_ = _0016_ ? addroundkey_data_o[89] : _2437_;
  assign next_addroundkey_data_reg[89] = _0004_ ? _2434_ : _2438_;
  assign _2439_ = ~key_i[8];
  assign _2440_ = ~subbytes_data_o[8];
  assign _2441_ = ~mixcol_data_o[8];
  assign _2442_ = ~data_i[8];
  assign _2443_ = _0459_ ? _2441_ : _2442_;
  assign _2444_ = _0455_ ? _2440_ : _2443_;
  assign _2445_ = _0470_ ? _2440_ : _2444_;
  assign _2446_ = _0469_ ? _2441_ : _2445_;
  assign _2447_ = subbytes_ready_o ? _2440_ : _2446_;
  assign _2448_ = _0468_ ? _2446_ : _2447_;
  assign _2449_ = _0463_ ? _2440_ : _2448_;
  assign _2450_ = _0450_ ? _2444_ : _2449_;
  assign _2451_ = _2450_ ^ _2439_;
  assign _2452_ = ~keysched_new_key_o[8];
  assign _2453_ = _2450_ ^ _2452_;
  assign _2454_ = _0479_ ? addroundkey_data_o[8] : _2453_;
  assign _2455_ = _0016_ ? addroundkey_data_o[8] : _2454_;
  assign next_addroundkey_data_reg[8] = _0004_ ? _2451_ : _2455_;
  assign _2456_ = ~key_i[90];
  assign _2457_ = ~subbytes_data_o[90];
  assign _2458_ = ~mixcol_data_o[90];
  assign _2459_ = ~data_i[90];
  assign _2460_ = _0459_ ? _2458_ : _2459_;
  assign _2461_ = _0455_ ? _2457_ : _2460_;
  assign _2462_ = _0470_ ? _2457_ : _2461_;
  assign _2463_ = _0469_ ? _2458_ : _2462_;
  assign _2464_ = subbytes_ready_o ? _2457_ : _2463_;
  assign _2465_ = _0468_ ? _2463_ : _2464_;
  assign _2466_ = _0463_ ? _2457_ : _2465_;
  assign _2467_ = _0450_ ? _2461_ : _2466_;
  assign _2468_ = _2467_ ^ _2456_;
  assign _2469_ = ~keysched_new_key_o[90];
  assign _2470_ = _2467_ ^ _2469_;
  assign _2471_ = _0479_ ? addroundkey_data_o[90] : _2470_;
  assign _2472_ = _0016_ ? addroundkey_data_o[90] : _2471_;
  assign next_addroundkey_data_reg[90] = _0004_ ? _2468_ : _2472_;
  assign _2473_ = ~key_i[91];
  assign _2474_ = ~subbytes_data_o[91];
  assign _2475_ = ~mixcol_data_o[91];
  assign _2476_ = ~data_i[91];
  assign _2477_ = _0459_ ? _2475_ : _2476_;
  assign _2478_ = _0455_ ? _2474_ : _2477_;
  assign _2479_ = _0470_ ? _2474_ : _2478_;
  assign _2480_ = _0469_ ? _2475_ : _2479_;
  assign _2481_ = subbytes_ready_o ? _2474_ : _2480_;
  assign _2482_ = _0468_ ? _2480_ : _2481_;
  assign _2483_ = _0463_ ? _2474_ : _2482_;
  assign _2484_ = _0450_ ? _2478_ : _2483_;
  assign _2485_ = _2484_ ^ _2473_;
  assign _2486_ = ~keysched_new_key_o[91];
  assign _2487_ = _2484_ ^ _2486_;
  assign _2488_ = _0479_ ? addroundkey_data_o[91] : _2487_;
  assign _2489_ = _0016_ ? addroundkey_data_o[91] : _2488_;
  assign next_addroundkey_data_reg[91] = _0004_ ? _2485_ : _2489_;
  assign _2490_ = ~key_i[92];
  assign _2491_ = ~subbytes_data_o[92];
  assign _2492_ = ~mixcol_data_o[92];
  assign _2493_ = ~data_i[92];
  assign _2494_ = _0459_ ? _2492_ : _2493_;
  assign _2495_ = _0455_ ? _2491_ : _2494_;
  assign _2496_ = _0470_ ? _2491_ : _2495_;
  assign _2497_ = _0469_ ? _2492_ : _2496_;
  assign _2498_ = subbytes_ready_o ? _2491_ : _2497_;
  assign _2499_ = _0468_ ? _2497_ : _2498_;
  assign _2500_ = _0463_ ? _2491_ : _2499_;
  assign _2501_ = _0450_ ? _2495_ : _2500_;
  assign _2502_ = _2501_ ^ _2490_;
  assign _2503_ = ~keysched_new_key_o[92];
  assign _2504_ = _2501_ ^ _2503_;
  assign _2505_ = _0479_ ? addroundkey_data_o[92] : _2504_;
  assign _2506_ = _0016_ ? addroundkey_data_o[92] : _2505_;
  assign next_addroundkey_data_reg[92] = _0004_ ? _2502_ : _2506_;
  assign _2507_ = ~key_i[93];
  assign _2508_ = ~subbytes_data_o[93];
  assign _2509_ = ~mixcol_data_o[93];
  assign _2510_ = ~data_i[93];
  assign _2511_ = _0459_ ? _2509_ : _2510_;
  assign _2512_ = _0455_ ? _2508_ : _2511_;
  assign _2513_ = _0470_ ? _2508_ : _2512_;
  assign _2514_ = _0469_ ? _2509_ : _2513_;
  assign _2515_ = subbytes_ready_o ? _2508_ : _2514_;
  assign _2516_ = _0468_ ? _2514_ : _2515_;
  assign _2517_ = _0463_ ? _2508_ : _2516_;
  assign _2518_ = _0450_ ? _2512_ : _2517_;
  assign _2519_ = _2518_ ^ _2507_;
  assign _2520_ = ~keysched_new_key_o[93];
  assign _2521_ = _2518_ ^ _2520_;
  assign _2522_ = _0479_ ? addroundkey_data_o[93] : _2521_;
  assign _2523_ = _0016_ ? addroundkey_data_o[93] : _2522_;
  assign next_addroundkey_data_reg[93] = _0004_ ? _2519_ : _2523_;
  assign _2524_ = ~key_i[94];
  assign _2525_ = ~subbytes_data_o[94];
  assign _2526_ = ~mixcol_data_o[94];
  assign _2527_ = ~data_i[94];
  assign _2528_ = _0459_ ? _2526_ : _2527_;
  assign _2529_ = _0455_ ? _2525_ : _2528_;
  assign _2530_ = _0470_ ? _2525_ : _2529_;
  assign _2531_ = _0469_ ? _2526_ : _2530_;
  assign _2532_ = subbytes_ready_o ? _2525_ : _2531_;
  assign _2533_ = _0468_ ? _2531_ : _2532_;
  assign _2534_ = _0463_ ? _2525_ : _2533_;
  assign _2535_ = _0450_ ? _2529_ : _2534_;
  assign _2536_ = _2535_ ^ _2524_;
  assign _2537_ = ~keysched_new_key_o[94];
  assign _2538_ = _2535_ ^ _2537_;
  assign _2539_ = _0479_ ? addroundkey_data_o[94] : _2538_;
  assign _2540_ = _0016_ ? addroundkey_data_o[94] : _2539_;
  assign next_addroundkey_data_reg[94] = _0004_ ? _2536_ : _2540_;
  assign _2541_ = ~key_i[95];
  assign _2542_ = ~subbytes_data_o[95];
  assign _2543_ = ~mixcol_data_o[95];
  assign _2544_ = ~data_i[95];
  assign _2545_ = _0459_ ? _2543_ : _2544_;
  assign _2546_ = _0455_ ? _2542_ : _2545_;
  assign _2547_ = _0470_ ? _2542_ : _2546_;
  assign _2548_ = _0469_ ? _2543_ : _2547_;
  assign _2549_ = subbytes_ready_o ? _2542_ : _2548_;
  assign _2550_ = _0468_ ? _2548_ : _2549_;
  assign _2551_ = _0463_ ? _2542_ : _2550_;
  assign _2552_ = _0450_ ? _2546_ : _2551_;
  assign _2553_ = _2552_ ^ _2541_;
  assign _2554_ = ~keysched_new_key_o[95];
  assign _2555_ = _2552_ ^ _2554_;
  assign _2556_ = _0479_ ? addroundkey_data_o[95] : _2555_;
  assign _2557_ = _0016_ ? addroundkey_data_o[95] : _2556_;
  assign next_addroundkey_data_reg[95] = _0004_ ? _2553_ : _2557_;
  assign _2558_ = ~key_i[96];
  assign _2559_ = ~subbytes_data_o[96];
  assign _2560_ = ~mixcol_data_o[96];
  assign _2561_ = ~data_i[96];
  assign _2562_ = _0459_ ? _2560_ : _2561_;
  assign _2563_ = _0455_ ? _2559_ : _2562_;
  assign _2564_ = _0470_ ? _2559_ : _2563_;
  assign _2565_ = _0469_ ? _2560_ : _2564_;
  assign _2566_ = subbytes_ready_o ? _2559_ : _2565_;
  assign _2567_ = _0468_ ? _2565_ : _2566_;
  assign _2568_ = _0463_ ? _2559_ : _2567_;
  assign _2569_ = _0450_ ? _2563_ : _2568_;
  assign _2570_ = _2569_ ^ _2558_;
  assign _2571_ = ~keysched_new_key_o[96];
  assign _2572_ = _2569_ ^ _2571_;
  assign _2573_ = _0479_ ? addroundkey_data_o[96] : _2572_;
  assign _2574_ = _0016_ ? addroundkey_data_o[96] : _2573_;
  assign next_addroundkey_data_reg[96] = _0004_ ? _2570_ : _2574_;
  assign _2575_ = ~key_i[97];
  assign _2576_ = ~subbytes_data_o[97];
  assign _2577_ = ~mixcol_data_o[97];
  assign _2578_ = ~data_i[97];
  assign _2579_ = _0459_ ? _2577_ : _2578_;
  assign _2580_ = _0455_ ? _2576_ : _2579_;
  assign _2581_ = _0470_ ? _2576_ : _2580_;
  assign _2582_ = _0469_ ? _2577_ : _2581_;
  assign _2583_ = subbytes_ready_o ? _2576_ : _2582_;
  assign _2584_ = _0468_ ? _2582_ : _2583_;
  assign _2585_ = _0463_ ? _2576_ : _2584_;
  assign _2586_ = _0450_ ? _2580_ : _2585_;
  assign _2587_ = _2586_ ^ _2575_;
  assign _2588_ = ~keysched_new_key_o[97];
  assign _2589_ = _2586_ ^ _2588_;
  assign _2590_ = _0479_ ? addroundkey_data_o[97] : _2589_;
  assign _2591_ = _0016_ ? addroundkey_data_o[97] : _2590_;
  assign next_addroundkey_data_reg[97] = _0004_ ? _2587_ : _2591_;
  assign _2592_ = ~key_i[98];
  assign _2593_ = ~subbytes_data_o[98];
  assign _2594_ = ~mixcol_data_o[98];
  assign _2595_ = ~data_i[98];
  assign _2596_ = _0459_ ? _2594_ : _2595_;
  assign _2597_ = _0455_ ? _2593_ : _2596_;
  assign _2598_ = _0470_ ? _2593_ : _2597_;
  assign _2599_ = _0469_ ? _2594_ : _2598_;
  assign _2600_ = subbytes_ready_o ? _2593_ : _2599_;
  assign _2601_ = _0468_ ? _2599_ : _2600_;
  assign _2602_ = _0463_ ? _2593_ : _2601_;
  assign _2603_ = _0450_ ? _2597_ : _2602_;
  assign _2604_ = _2603_ ^ _2592_;
  assign _2605_ = ~keysched_new_key_o[98];
  assign _2606_ = _2603_ ^ _2605_;
  assign _2607_ = _0479_ ? addroundkey_data_o[98] : _2606_;
  assign _2608_ = _0016_ ? addroundkey_data_o[98] : _2607_;
  assign next_addroundkey_data_reg[98] = _0004_ ? _2604_ : _2608_;
  assign _2609_ = ~key_i[99];
  assign _2610_ = ~subbytes_data_o[99];
  assign _2611_ = ~mixcol_data_o[99];
  assign _2612_ = ~data_i[99];
  assign _2613_ = _0459_ ? _2611_ : _2612_;
  assign _2614_ = _0455_ ? _2610_ : _2613_;
  assign _2615_ = _0470_ ? _2610_ : _2614_;
  assign _2616_ = _0469_ ? _2611_ : _2615_;
  assign _2617_ = subbytes_ready_o ? _2610_ : _2616_;
  assign _2618_ = _0468_ ? _2616_ : _2617_;
  assign _2619_ = _0463_ ? _2610_ : _2618_;
  assign _2620_ = _0450_ ? _2614_ : _2619_;
  assign _2621_ = _2620_ ^ _2609_;
  assign _2622_ = ~keysched_new_key_o[99];
  assign _2623_ = _2620_ ^ _2622_;
  assign _2624_ = _0479_ ? addroundkey_data_o[99] : _2623_;
  assign _2625_ = _0016_ ? addroundkey_data_o[99] : _2624_;
  assign next_addroundkey_data_reg[99] = _0004_ ? _2621_ : _2625_;
  assign _2626_ = ~key_i[9];
  assign _2627_ = ~subbytes_data_o[9];
  assign _2628_ = ~mixcol_data_o[9];
  assign _2629_ = ~data_i[9];
  assign _2630_ = _0459_ ? _2628_ : _2629_;
  assign _2631_ = _0455_ ? _2627_ : _2630_;
  assign _2632_ = _0470_ ? _2627_ : _2631_;
  assign _2633_ = _0469_ ? _2628_ : _2632_;
  assign _2634_ = subbytes_ready_o ? _2627_ : _2633_;
  assign _2635_ = _0468_ ? _2633_ : _2634_;
  assign _2636_ = _0463_ ? _2627_ : _2635_;
  assign _2637_ = _0450_ ? _2631_ : _2636_;
  assign _2638_ = _2637_ ^ _2626_;
  assign _2639_ = ~keysched_new_key_o[9];
  assign _2640_ = _2637_ ^ _2639_;
  assign _2641_ = _0479_ ? addroundkey_data_o[9] : _2640_;
  assign _2642_ = _0016_ ? addroundkey_data_o[9] : _2641_;
  assign next_addroundkey_data_reg[9] = _0004_ ? _2638_ : _2642_;
  assign _2643_ = ~_0029_;
  assign _2644_ = _0420_ & _2643_;
  assign _2645_ = _2644_ & _0478_;
  assign next_addroundkey_ready_o = _2645_ | _0004_;
  assign sbox_decrypt_i = keysched_sbox_access_o ? keysched_sbox_decrypt_o : subbytes_sbox_decrypt_o;
  assign sbox_data_i[0] = keysched_sbox_access_o ? keysched_sbox_data_o[0] : subbytes_sbox_data_o[0];
  assign sbox_data_i[1] = keysched_sbox_access_o ? keysched_sbox_data_o[1] : subbytes_sbox_data_o[1];
  assign sbox_data_i[2] = keysched_sbox_access_o ? keysched_sbox_data_o[2] : subbytes_sbox_data_o[2];
  assign sbox_data_i[3] = keysched_sbox_access_o ? keysched_sbox_data_o[3] : subbytes_sbox_data_o[3];
  assign sbox_data_i[4] = keysched_sbox_access_o ? keysched_sbox_data_o[4] : subbytes_sbox_data_o[4];
  assign sbox_data_i[5] = keysched_sbox_access_o ? keysched_sbox_data_o[5] : subbytes_sbox_data_o[5];
  assign sbox_data_i[6] = keysched_sbox_access_o ? keysched_sbox_data_o[6] : subbytes_sbox_data_o[6];
  assign sbox_data_i[7] = keysched_sbox_access_o ? keysched_sbox_data_o[7] : subbytes_sbox_data_o[7];
  assign subbytes_data_i[0] = _0455_ ? mixcol_data_o[0] : addroundkey_data_o[0];
  assign subbytes_data_i[100] = _0455_ ? mixcol_data_o[100] : addroundkey_data_o[100];
  assign subbytes_data_i[101] = _0455_ ? mixcol_data_o[101] : addroundkey_data_o[101];
  assign subbytes_data_i[102] = _0455_ ? mixcol_data_o[102] : addroundkey_data_o[102];
  assign subbytes_data_i[103] = _0455_ ? mixcol_data_o[103] : addroundkey_data_o[103];
  assign subbytes_data_i[104] = _0455_ ? mixcol_data_o[104] : addroundkey_data_o[104];
  assign subbytes_data_i[105] = _0455_ ? mixcol_data_o[105] : addroundkey_data_o[105];
  assign subbytes_data_i[106] = _0455_ ? mixcol_data_o[106] : addroundkey_data_o[106];
  assign subbytes_data_i[107] = _0455_ ? mixcol_data_o[107] : addroundkey_data_o[107];
  assign subbytes_data_i[108] = _0455_ ? mixcol_data_o[108] : addroundkey_data_o[108];
  assign subbytes_data_i[109] = _0455_ ? mixcol_data_o[109] : addroundkey_data_o[109];
  assign subbytes_data_i[10] = _0455_ ? mixcol_data_o[10] : addroundkey_data_o[10];
  assign subbytes_data_i[110] = _0455_ ? mixcol_data_o[110] : addroundkey_data_o[110];
  assign subbytes_data_i[111] = _0455_ ? mixcol_data_o[111] : addroundkey_data_o[111];
  assign subbytes_data_i[112] = _0455_ ? mixcol_data_o[112] : addroundkey_data_o[112];
  assign subbytes_data_i[113] = _0455_ ? mixcol_data_o[113] : addroundkey_data_o[113];
  assign subbytes_data_i[114] = _0455_ ? mixcol_data_o[114] : addroundkey_data_o[114];
  assign subbytes_data_i[115] = _0455_ ? mixcol_data_o[115] : addroundkey_data_o[115];
  assign subbytes_data_i[116] = _0455_ ? mixcol_data_o[116] : addroundkey_data_o[116];
  assign subbytes_data_i[117] = _0455_ ? mixcol_data_o[117] : addroundkey_data_o[117];
  assign subbytes_data_i[118] = _0455_ ? mixcol_data_o[118] : addroundkey_data_o[118];
  assign subbytes_data_i[119] = _0455_ ? mixcol_data_o[119] : addroundkey_data_o[119];
  assign subbytes_data_i[11] = _0455_ ? mixcol_data_o[11] : addroundkey_data_o[11];
  assign subbytes_data_i[120] = _0455_ ? mixcol_data_o[120] : addroundkey_data_o[120];
  assign subbytes_data_i[121] = _0455_ ? mixcol_data_o[121] : addroundkey_data_o[121];
  assign subbytes_data_i[122] = _0455_ ? mixcol_data_o[122] : addroundkey_data_o[122];
  assign subbytes_data_i[123] = _0455_ ? mixcol_data_o[123] : addroundkey_data_o[123];
  assign subbytes_data_i[124] = _0455_ ? mixcol_data_o[124] : addroundkey_data_o[124];
  assign subbytes_data_i[125] = _0455_ ? mixcol_data_o[125] : addroundkey_data_o[125];
  assign subbytes_data_i[126] = _0455_ ? mixcol_data_o[126] : addroundkey_data_o[126];
  assign subbytes_data_i[127] = _0455_ ? mixcol_data_o[127] : addroundkey_data_o[127];
  assign subbytes_data_i[12] = _0455_ ? mixcol_data_o[12] : addroundkey_data_o[12];
  assign subbytes_data_i[13] = _0455_ ? mixcol_data_o[13] : addroundkey_data_o[13];
  assign subbytes_data_i[14] = _0455_ ? mixcol_data_o[14] : addroundkey_data_o[14];
  assign subbytes_data_i[15] = _0455_ ? mixcol_data_o[15] : addroundkey_data_o[15];
  assign subbytes_data_i[16] = _0455_ ? mixcol_data_o[16] : addroundkey_data_o[16];
  assign subbytes_data_i[17] = _0455_ ? mixcol_data_o[17] : addroundkey_data_o[17];
  assign subbytes_data_i[18] = _0455_ ? mixcol_data_o[18] : addroundkey_data_o[18];
  assign subbytes_data_i[19] = _0455_ ? mixcol_data_o[19] : addroundkey_data_o[19];
  assign subbytes_data_i[1] = _0455_ ? mixcol_data_o[1] : addroundkey_data_o[1];
  assign subbytes_data_i[20] = _0455_ ? mixcol_data_o[20] : addroundkey_data_o[20];
  assign subbytes_data_i[21] = _0455_ ? mixcol_data_o[21] : addroundkey_data_o[21];
  assign subbytes_data_i[22] = _0455_ ? mixcol_data_o[22] : addroundkey_data_o[22];
  assign subbytes_data_i[23] = _0455_ ? mixcol_data_o[23] : addroundkey_data_o[23];
  assign subbytes_data_i[24] = _0455_ ? mixcol_data_o[24] : addroundkey_data_o[24];
  assign subbytes_data_i[25] = _0455_ ? mixcol_data_o[25] : addroundkey_data_o[25];
  assign subbytes_data_i[26] = _0455_ ? mixcol_data_o[26] : addroundkey_data_o[26];
  assign subbytes_data_i[27] = _0455_ ? mixcol_data_o[27] : addroundkey_data_o[27];
  assign subbytes_data_i[28] = _0455_ ? mixcol_data_o[28] : addroundkey_data_o[28];
  assign subbytes_data_i[29] = _0455_ ? mixcol_data_o[29] : addroundkey_data_o[29];
  assign subbytes_data_i[2] = _0455_ ? mixcol_data_o[2] : addroundkey_data_o[2];
  assign subbytes_data_i[30] = _0455_ ? mixcol_data_o[30] : addroundkey_data_o[30];
  assign subbytes_data_i[31] = _0455_ ? mixcol_data_o[31] : addroundkey_data_o[31];
  assign subbytes_data_i[32] = _0455_ ? mixcol_data_o[32] : addroundkey_data_o[32];
  assign subbytes_data_i[33] = _0455_ ? mixcol_data_o[33] : addroundkey_data_o[33];
  assign subbytes_data_i[34] = _0455_ ? mixcol_data_o[34] : addroundkey_data_o[34];
  assign subbytes_data_i[35] = _0455_ ? mixcol_data_o[35] : addroundkey_data_o[35];
  assign subbytes_data_i[36] = _0455_ ? mixcol_data_o[36] : addroundkey_data_o[36];
  assign subbytes_data_i[37] = _0455_ ? mixcol_data_o[37] : addroundkey_data_o[37];
  assign subbytes_data_i[38] = _0455_ ? mixcol_data_o[38] : addroundkey_data_o[38];
  assign subbytes_data_i[39] = _0455_ ? mixcol_data_o[39] : addroundkey_data_o[39];
  assign subbytes_data_i[3] = _0455_ ? mixcol_data_o[3] : addroundkey_data_o[3];
  assign subbytes_data_i[40] = _0455_ ? mixcol_data_o[40] : addroundkey_data_o[40];
  assign subbytes_data_i[41] = _0455_ ? mixcol_data_o[41] : addroundkey_data_o[41];
  assign subbytes_data_i[42] = _0455_ ? mixcol_data_o[42] : addroundkey_data_o[42];
  assign subbytes_data_i[43] = _0455_ ? mixcol_data_o[43] : addroundkey_data_o[43];
  assign subbytes_data_i[44] = _0455_ ? mixcol_data_o[44] : addroundkey_data_o[44];
  assign subbytes_data_i[45] = _0455_ ? mixcol_data_o[45] : addroundkey_data_o[45];
  assign subbytes_data_i[46] = _0455_ ? mixcol_data_o[46] : addroundkey_data_o[46];
  assign subbytes_data_i[47] = _0455_ ? mixcol_data_o[47] : addroundkey_data_o[47];
  assign subbytes_data_i[48] = _0455_ ? mixcol_data_o[48] : addroundkey_data_o[48];
  assign subbytes_data_i[49] = _0455_ ? mixcol_data_o[49] : addroundkey_data_o[49];
  assign subbytes_data_i[4] = _0455_ ? mixcol_data_o[4] : addroundkey_data_o[4];
  assign subbytes_data_i[50] = _0455_ ? mixcol_data_o[50] : addroundkey_data_o[50];
  assign subbytes_data_i[51] = _0455_ ? mixcol_data_o[51] : addroundkey_data_o[51];
  assign subbytes_data_i[52] = _0455_ ? mixcol_data_o[52] : addroundkey_data_o[52];
  assign subbytes_data_i[53] = _0455_ ? mixcol_data_o[53] : addroundkey_data_o[53];
  assign subbytes_data_i[54] = _0455_ ? mixcol_data_o[54] : addroundkey_data_o[54];
  assign subbytes_data_i[55] = _0455_ ? mixcol_data_o[55] : addroundkey_data_o[55];
  assign subbytes_data_i[56] = _0455_ ? mixcol_data_o[56] : addroundkey_data_o[56];
  assign subbytes_data_i[57] = _0455_ ? mixcol_data_o[57] : addroundkey_data_o[57];
  assign subbytes_data_i[58] = _0455_ ? mixcol_data_o[58] : addroundkey_data_o[58];
  assign subbytes_data_i[59] = _0455_ ? mixcol_data_o[59] : addroundkey_data_o[59];
  assign subbytes_data_i[5] = _0455_ ? mixcol_data_o[5] : addroundkey_data_o[5];
  assign subbytes_data_i[60] = _0455_ ? mixcol_data_o[60] : addroundkey_data_o[60];
  assign subbytes_data_i[61] = _0455_ ? mixcol_data_o[61] : addroundkey_data_o[61];
  assign subbytes_data_i[62] = _0455_ ? mixcol_data_o[62] : addroundkey_data_o[62];
  assign subbytes_data_i[63] = _0455_ ? mixcol_data_o[63] : addroundkey_data_o[63];
  assign subbytes_data_i[64] = _0455_ ? mixcol_data_o[64] : addroundkey_data_o[64];
  assign subbytes_data_i[65] = _0455_ ? mixcol_data_o[65] : addroundkey_data_o[65];
  assign subbytes_data_i[66] = _0455_ ? mixcol_data_o[66] : addroundkey_data_o[66];
  assign subbytes_data_i[67] = _0455_ ? mixcol_data_o[67] : addroundkey_data_o[67];
  assign subbytes_data_i[68] = _0455_ ? mixcol_data_o[68] : addroundkey_data_o[68];
  assign subbytes_data_i[69] = _0455_ ? mixcol_data_o[69] : addroundkey_data_o[69];
  assign subbytes_data_i[6] = _0455_ ? mixcol_data_o[6] : addroundkey_data_o[6];
  assign subbytes_data_i[70] = _0455_ ? mixcol_data_o[70] : addroundkey_data_o[70];
  assign subbytes_data_i[71] = _0455_ ? mixcol_data_o[71] : addroundkey_data_o[71];
  assign subbytes_data_i[72] = _0455_ ? mixcol_data_o[72] : addroundkey_data_o[72];
  assign subbytes_data_i[73] = _0455_ ? mixcol_data_o[73] : addroundkey_data_o[73];
  assign subbytes_data_i[74] = _0455_ ? mixcol_data_o[74] : addroundkey_data_o[74];
  assign subbytes_data_i[75] = _0455_ ? mixcol_data_o[75] : addroundkey_data_o[75];
  assign subbytes_data_i[76] = _0455_ ? mixcol_data_o[76] : addroundkey_data_o[76];
  assign subbytes_data_i[77] = _0455_ ? mixcol_data_o[77] : addroundkey_data_o[77];
  assign subbytes_data_i[78] = _0455_ ? mixcol_data_o[78] : addroundkey_data_o[78];
  assign subbytes_data_i[79] = _0455_ ? mixcol_data_o[79] : addroundkey_data_o[79];
  assign subbytes_data_i[7] = _0455_ ? mixcol_data_o[7] : addroundkey_data_o[7];
  assign subbytes_data_i[80] = _0455_ ? mixcol_data_o[80] : addroundkey_data_o[80];
  assign subbytes_data_i[81] = _0455_ ? mixcol_data_o[81] : addroundkey_data_o[81];
  assign subbytes_data_i[82] = _0455_ ? mixcol_data_o[82] : addroundkey_data_o[82];
  assign subbytes_data_i[83] = _0455_ ? mixcol_data_o[83] : addroundkey_data_o[83];
  assign subbytes_data_i[84] = _0455_ ? mixcol_data_o[84] : addroundkey_data_o[84];
  assign subbytes_data_i[85] = _0455_ ? mixcol_data_o[85] : addroundkey_data_o[85];
  assign subbytes_data_i[86] = _0455_ ? mixcol_data_o[86] : addroundkey_data_o[86];
  assign subbytes_data_i[87] = _0455_ ? mixcol_data_o[87] : addroundkey_data_o[87];
  assign subbytes_data_i[88] = _0455_ ? mixcol_data_o[88] : addroundkey_data_o[88];
  assign subbytes_data_i[89] = _0455_ ? mixcol_data_o[89] : addroundkey_data_o[89];
  assign subbytes_data_i[8] = _0455_ ? mixcol_data_o[8] : addroundkey_data_o[8];
  assign subbytes_data_i[90] = _0455_ ? mixcol_data_o[90] : addroundkey_data_o[90];
  assign subbytes_data_i[91] = _0455_ ? mixcol_data_o[91] : addroundkey_data_o[91];
  assign subbytes_data_i[92] = _0455_ ? mixcol_data_o[92] : addroundkey_data_o[92];
  assign subbytes_data_i[93] = _0455_ ? mixcol_data_o[93] : addroundkey_data_o[93];
  assign subbytes_data_i[94] = _0455_ ? mixcol_data_o[94] : addroundkey_data_o[94];
  assign subbytes_data_i[95] = _0455_ ? mixcol_data_o[95] : addroundkey_data_o[95];
  assign subbytes_data_i[96] = _0455_ ? mixcol_data_o[96] : addroundkey_data_o[96];
  assign subbytes_data_i[97] = _0455_ ? mixcol_data_o[97] : addroundkey_data_o[97];
  assign subbytes_data_i[98] = _0455_ ? mixcol_data_o[98] : addroundkey_data_o[98];
  assign subbytes_data_i[99] = _0455_ ? mixcol_data_o[99] : addroundkey_data_o[99];
  assign subbytes_data_i[9] = _0455_ ? mixcol_data_o[9] : addroundkey_data_o[9];
  assign mixcol_data_i[0] = _0455_ ? addroundkey_data_o[0] : subbytes_data_o[0];
  assign mixcol_data_i[100] = _0455_ ? addroundkey_data_o[100] : subbytes_data_o[100];
  assign mixcol_data_i[101] = _0455_ ? addroundkey_data_o[101] : subbytes_data_o[101];
  assign mixcol_data_i[102] = _0455_ ? addroundkey_data_o[102] : subbytes_data_o[102];
  assign mixcol_data_i[103] = _0455_ ? addroundkey_data_o[103] : subbytes_data_o[103];
  assign mixcol_data_i[104] = _0455_ ? addroundkey_data_o[104] : subbytes_data_o[104];
  assign mixcol_data_i[105] = _0455_ ? addroundkey_data_o[105] : subbytes_data_o[105];
  assign mixcol_data_i[106] = _0455_ ? addroundkey_data_o[106] : subbytes_data_o[106];
  assign mixcol_data_i[107] = _0455_ ? addroundkey_data_o[107] : subbytes_data_o[107];
  assign mixcol_data_i[108] = _0455_ ? addroundkey_data_o[108] : subbytes_data_o[108];
  assign mixcol_data_i[109] = _0455_ ? addroundkey_data_o[109] : subbytes_data_o[109];
  assign mixcol_data_i[10] = _0455_ ? addroundkey_data_o[10] : subbytes_data_o[10];
  assign mixcol_data_i[110] = _0455_ ? addroundkey_data_o[110] : subbytes_data_o[110];
  assign mixcol_data_i[111] = _0455_ ? addroundkey_data_o[111] : subbytes_data_o[111];
  assign mixcol_data_i[112] = _0455_ ? addroundkey_data_o[112] : subbytes_data_o[112];
  assign mixcol_data_i[113] = _0455_ ? addroundkey_data_o[113] : subbytes_data_o[113];
  assign mixcol_data_i[114] = _0455_ ? addroundkey_data_o[114] : subbytes_data_o[114];
  assign mixcol_data_i[115] = _0455_ ? addroundkey_data_o[115] : subbytes_data_o[115];
  assign mixcol_data_i[116] = _0455_ ? addroundkey_data_o[116] : subbytes_data_o[116];
  assign mixcol_data_i[117] = _0455_ ? addroundkey_data_o[117] : subbytes_data_o[117];
  assign mixcol_data_i[118] = _0455_ ? addroundkey_data_o[118] : subbytes_data_o[118];
  assign mixcol_data_i[119] = _0455_ ? addroundkey_data_o[119] : subbytes_data_o[119];
  assign mixcol_data_i[11] = _0455_ ? addroundkey_data_o[11] : subbytes_data_o[11];
  assign mixcol_data_i[120] = _0455_ ? addroundkey_data_o[120] : subbytes_data_o[120];
  assign mixcol_data_i[121] = _0455_ ? addroundkey_data_o[121] : subbytes_data_o[121];
  assign mixcol_data_i[122] = _0455_ ? addroundkey_data_o[122] : subbytes_data_o[122];
  assign mixcol_data_i[123] = _0455_ ? addroundkey_data_o[123] : subbytes_data_o[123];
  assign mixcol_data_i[124] = _0455_ ? addroundkey_data_o[124] : subbytes_data_o[124];
  assign mixcol_data_i[125] = _0455_ ? addroundkey_data_o[125] : subbytes_data_o[125];
  assign mixcol_data_i[126] = _0455_ ? addroundkey_data_o[126] : subbytes_data_o[126];
  assign mixcol_data_i[127] = _0455_ ? addroundkey_data_o[127] : subbytes_data_o[127];
  assign mixcol_data_i[12] = _0455_ ? addroundkey_data_o[12] : subbytes_data_o[12];
  assign mixcol_data_i[13] = _0455_ ? addroundkey_data_o[13] : subbytes_data_o[13];
  assign mixcol_data_i[14] = _0455_ ? addroundkey_data_o[14] : subbytes_data_o[14];
  assign mixcol_data_i[15] = _0455_ ? addroundkey_data_o[15] : subbytes_data_o[15];
  assign mixcol_data_i[16] = _0455_ ? addroundkey_data_o[16] : subbytes_data_o[16];
  assign mixcol_data_i[17] = _0455_ ? addroundkey_data_o[17] : subbytes_data_o[17];
  assign mixcol_data_i[18] = _0455_ ? addroundkey_data_o[18] : subbytes_data_o[18];
  assign mixcol_data_i[19] = _0455_ ? addroundkey_data_o[19] : subbytes_data_o[19];
  assign mixcol_data_i[1] = _0455_ ? addroundkey_data_o[1] : subbytes_data_o[1];
  assign mixcol_data_i[20] = _0455_ ? addroundkey_data_o[20] : subbytes_data_o[20];
  assign mixcol_data_i[21] = _0455_ ? addroundkey_data_o[21] : subbytes_data_o[21];
  assign mixcol_data_i[22] = _0455_ ? addroundkey_data_o[22] : subbytes_data_o[22];
  assign mixcol_data_i[23] = _0455_ ? addroundkey_data_o[23] : subbytes_data_o[23];
  assign mixcol_data_i[24] = _0455_ ? addroundkey_data_o[24] : subbytes_data_o[24];
  assign mixcol_data_i[25] = _0455_ ? addroundkey_data_o[25] : subbytes_data_o[25];
  assign mixcol_data_i[26] = _0455_ ? addroundkey_data_o[26] : subbytes_data_o[26];
  assign mixcol_data_i[27] = _0455_ ? addroundkey_data_o[27] : subbytes_data_o[27];
  assign mixcol_data_i[28] = _0455_ ? addroundkey_data_o[28] : subbytes_data_o[28];
  assign mixcol_data_i[29] = _0455_ ? addroundkey_data_o[29] : subbytes_data_o[29];
  assign mixcol_data_i[2] = _0455_ ? addroundkey_data_o[2] : subbytes_data_o[2];
  assign mixcol_data_i[30] = _0455_ ? addroundkey_data_o[30] : subbytes_data_o[30];
  assign mixcol_data_i[31] = _0455_ ? addroundkey_data_o[31] : subbytes_data_o[31];
  assign mixcol_data_i[32] = _0455_ ? addroundkey_data_o[32] : subbytes_data_o[32];
  assign mixcol_data_i[33] = _0455_ ? addroundkey_data_o[33] : subbytes_data_o[33];
  assign mixcol_data_i[34] = _0455_ ? addroundkey_data_o[34] : subbytes_data_o[34];
  assign mixcol_data_i[35] = _0455_ ? addroundkey_data_o[35] : subbytes_data_o[35];
  assign mixcol_data_i[36] = _0455_ ? addroundkey_data_o[36] : subbytes_data_o[36];
  assign mixcol_data_i[37] = _0455_ ? addroundkey_data_o[37] : subbytes_data_o[37];
  assign mixcol_data_i[38] = _0455_ ? addroundkey_data_o[38] : subbytes_data_o[38];
  assign mixcol_data_i[39] = _0455_ ? addroundkey_data_o[39] : subbytes_data_o[39];
  assign mixcol_data_i[3] = _0455_ ? addroundkey_data_o[3] : subbytes_data_o[3];
  assign mixcol_data_i[40] = _0455_ ? addroundkey_data_o[40] : subbytes_data_o[40];
  assign mixcol_data_i[41] = _0455_ ? addroundkey_data_o[41] : subbytes_data_o[41];
  assign mixcol_data_i[42] = _0455_ ? addroundkey_data_o[42] : subbytes_data_o[42];
  assign mixcol_data_i[43] = _0455_ ? addroundkey_data_o[43] : subbytes_data_o[43];
  assign mixcol_data_i[44] = _0455_ ? addroundkey_data_o[44] : subbytes_data_o[44];
  assign mixcol_data_i[45] = _0455_ ? addroundkey_data_o[45] : subbytes_data_o[45];
  assign mixcol_data_i[46] = _0455_ ? addroundkey_data_o[46] : subbytes_data_o[46];
  assign mixcol_data_i[47] = _0455_ ? addroundkey_data_o[47] : subbytes_data_o[47];
  assign mixcol_data_i[48] = _0455_ ? addroundkey_data_o[48] : subbytes_data_o[48];
  assign mixcol_data_i[49] = _0455_ ? addroundkey_data_o[49] : subbytes_data_o[49];
  assign mixcol_data_i[4] = _0455_ ? addroundkey_data_o[4] : subbytes_data_o[4];
  assign mixcol_data_i[50] = _0455_ ? addroundkey_data_o[50] : subbytes_data_o[50];
  assign mixcol_data_i[51] = _0455_ ? addroundkey_data_o[51] : subbytes_data_o[51];
  assign mixcol_data_i[52] = _0455_ ? addroundkey_data_o[52] : subbytes_data_o[52];
  assign mixcol_data_i[53] = _0455_ ? addroundkey_data_o[53] : subbytes_data_o[53];
  assign mixcol_data_i[54] = _0455_ ? addroundkey_data_o[54] : subbytes_data_o[54];
  assign mixcol_data_i[55] = _0455_ ? addroundkey_data_o[55] : subbytes_data_o[55];
  assign mixcol_data_i[56] = _0455_ ? addroundkey_data_o[56] : subbytes_data_o[56];
  assign mixcol_data_i[57] = _0455_ ? addroundkey_data_o[57] : subbytes_data_o[57];
  assign mixcol_data_i[58] = _0455_ ? addroundkey_data_o[58] : subbytes_data_o[58];
  assign mixcol_data_i[59] = _0455_ ? addroundkey_data_o[59] : subbytes_data_o[59];
  assign mixcol_data_i[5] = _0455_ ? addroundkey_data_o[5] : subbytes_data_o[5];
  assign mixcol_data_i[60] = _0455_ ? addroundkey_data_o[60] : subbytes_data_o[60];
  assign mixcol_data_i[61] = _0455_ ? addroundkey_data_o[61] : subbytes_data_o[61];
  assign mixcol_data_i[62] = _0455_ ? addroundkey_data_o[62] : subbytes_data_o[62];
  assign mixcol_data_i[63] = _0455_ ? addroundkey_data_o[63] : subbytes_data_o[63];
  assign mixcol_data_i[64] = _0455_ ? addroundkey_data_o[64] : subbytes_data_o[64];
  assign mixcol_data_i[65] = _0455_ ? addroundkey_data_o[65] : subbytes_data_o[65];
  assign mixcol_data_i[66] = _0455_ ? addroundkey_data_o[66] : subbytes_data_o[66];
  assign mixcol_data_i[67] = _0455_ ? addroundkey_data_o[67] : subbytes_data_o[67];
  assign mixcol_data_i[68] = _0455_ ? addroundkey_data_o[68] : subbytes_data_o[68];
  assign mixcol_data_i[69] = _0455_ ? addroundkey_data_o[69] : subbytes_data_o[69];
  assign mixcol_data_i[6] = _0455_ ? addroundkey_data_o[6] : subbytes_data_o[6];
  assign mixcol_data_i[70] = _0455_ ? addroundkey_data_o[70] : subbytes_data_o[70];
  assign mixcol_data_i[71] = _0455_ ? addroundkey_data_o[71] : subbytes_data_o[71];
  assign mixcol_data_i[72] = _0455_ ? addroundkey_data_o[72] : subbytes_data_o[72];
  assign mixcol_data_i[73] = _0455_ ? addroundkey_data_o[73] : subbytes_data_o[73];
  assign mixcol_data_i[74] = _0455_ ? addroundkey_data_o[74] : subbytes_data_o[74];
  assign mixcol_data_i[75] = _0455_ ? addroundkey_data_o[75] : subbytes_data_o[75];
  assign mixcol_data_i[76] = _0455_ ? addroundkey_data_o[76] : subbytes_data_o[76];
  assign mixcol_data_i[77] = _0455_ ? addroundkey_data_o[77] : subbytes_data_o[77];
  assign mixcol_data_i[78] = _0455_ ? addroundkey_data_o[78] : subbytes_data_o[78];
  assign mixcol_data_i[79] = _0455_ ? addroundkey_data_o[79] : subbytes_data_o[79];
  assign mixcol_data_i[7] = _0455_ ? addroundkey_data_o[7] : subbytes_data_o[7];
  assign mixcol_data_i[80] = _0455_ ? addroundkey_data_o[80] : subbytes_data_o[80];
  assign mixcol_data_i[81] = _0455_ ? addroundkey_data_o[81] : subbytes_data_o[81];
  assign mixcol_data_i[82] = _0455_ ? addroundkey_data_o[82] : subbytes_data_o[82];
  assign mixcol_data_i[83] = _0455_ ? addroundkey_data_o[83] : subbytes_data_o[83];
  assign mixcol_data_i[84] = _0455_ ? addroundkey_data_o[84] : subbytes_data_o[84];
  assign mixcol_data_i[85] = _0455_ ? addroundkey_data_o[85] : subbytes_data_o[85];
  assign mixcol_data_i[86] = _0455_ ? addroundkey_data_o[86] : subbytes_data_o[86];
  assign mixcol_data_i[87] = _0455_ ? addroundkey_data_o[87] : subbytes_data_o[87];
  assign mixcol_data_i[88] = _0455_ ? addroundkey_data_o[88] : subbytes_data_o[88];
  assign mixcol_data_i[89] = _0455_ ? addroundkey_data_o[89] : subbytes_data_o[89];
  assign mixcol_data_i[8] = _0455_ ? addroundkey_data_o[8] : subbytes_data_o[8];
  assign mixcol_data_i[90] = _0455_ ? addroundkey_data_o[90] : subbytes_data_o[90];
  assign mixcol_data_i[91] = _0455_ ? addroundkey_data_o[91] : subbytes_data_o[91];
  assign mixcol_data_i[92] = _0455_ ? addroundkey_data_o[92] : subbytes_data_o[92];
  assign mixcol_data_i[93] = _0455_ ? addroundkey_data_o[93] : subbytes_data_o[93];
  assign mixcol_data_i[94] = _0455_ ? addroundkey_data_o[94] : subbytes_data_o[94];
  assign mixcol_data_i[95] = _0455_ ? addroundkey_data_o[95] : subbytes_data_o[95];
  assign mixcol_data_i[96] = _0455_ ? addroundkey_data_o[96] : subbytes_data_o[96];
  assign mixcol_data_i[97] = _0455_ ? addroundkey_data_o[97] : subbytes_data_o[97];
  assign mixcol_data_i[98] = _0455_ ? addroundkey_data_o[98] : subbytes_data_o[98];
  assign mixcol_data_i[99] = _0455_ ? addroundkey_data_o[99] : subbytes_data_o[99];
  assign mixcol_data_i[9] = _0455_ ? addroundkey_data_o[9] : subbytes_data_o[9];
  assign _2646_ = addroundkey_ready_o & decrypt_i;
  assign _2647_ = _2646_ & _0454_;
  assign _2648_ = subbytes_ready_o & _0458_;
  assign _2649_ = _2648_ | _2647_;
  assign _2650_ = _2649_ & _0450_;
  assign _2651_ = _0468_ & state;
  assign _2652_ = _2651_ & _2649_;
  assign mixcol_start_i = _2652_ | _2650_;
  assign _2653_ = _0470_ | first_round_reg;
  assign _2654_ = _2653_ | _0469_;
  assign _2655_ = _0468_ ? _2654_ : subbytes_ready_o;
  assign _2656_ = ~addroundkey_ready_o;
  assign _2657_ = _0463_ & _2656_;
  assign _2658_ = _2657_ & _2655_;
  assign _2659_ = _2655_ & _0462_;
  assign _2660_ = _2659_ | _2658_;
  assign next_addroundkey_start_i = _0450_ ? first_round_reg : _2660_;
  assign _2661_ = state & addroundkey_ready_o;
  assign next_ready_o = _2661_ & _0463_;
  assign _2662_ = ~_0454_;
  assign _2663_ = _2646_ & _2662_;
  assign _2664_ = decrypt_i ? mixcol_ready_o : addroundkey_ready_o;
  assign _2665_ = _2664_ | _2663_;
  assign _2666_ = _2665_ & _0450_;
  assign _2667_ = _0462_ & state;
  assign _2668_ = _2667_ & _2665_;
  assign subbytes_start_i = _2668_ | _2666_;
  assign next_first_round_reg = _0450_ & load_i;
  assign _2669_ = ~load_i;
  assign _2670_ = _2669_ & round[0];
  assign _2671_ = _0470_ ^ round[0];
  assign _2672_ = _0469_ ? _0019_ : _2671_;
  assign _2673_ = subbytes_ready_o ? _0019_ : _2672_;
  assign _2674_ = _0468_ ? _2672_ : _2673_;
  assign _2675_ = _2674_ & _2657_;
  assign _2676_ = _2674_ & _0462_;
  assign _2677_ = _2676_ | _2675_;
  assign next_round[0] = _0450_ ? _2670_ : _2677_;
  assign _2678_ = load_i ? decrypt_i : round[1];
  assign _2679_ = round[1] ^ round[0];
  assign _2680_ = ~_0470_;
  assign _2681_ = round[1] ^ _0019_;
  assign _2682_ = _2680_ ? round[1] : _2681_;
  assign _2683_ = _0469_ ? _2679_ : _2682_;
  assign _2684_ = subbytes_ready_o ? _2679_ : _2683_;
  assign _2685_ = _0468_ ? _2683_ : _2684_;
  assign _2686_ = _2685_ & _2657_;
  assign _2687_ = _2685_ & _0462_;
  assign _2688_ = _2687_ | _2686_;
  assign next_round[1] = _0450_ ? _2678_ : _2688_;
  assign _2689_ = _2669_ & round[2];
  assign _2690_ = round[1] & round[0];
  assign _2691_ = _2690_ ^ round[2];
  assign _2692_ = _0000_ ^ _0024_;
  assign _2693_ = _2680_ ? round[2] : _2692_;
  assign _2694_ = _0469_ ? _2691_ : _2693_;
  assign _2695_ = subbytes_ready_o ? _2691_ : _2694_;
  assign _2696_ = _0468_ ? _2694_ : _2695_;
  assign next_round[2] = _0450_ ? _2689_ : _2696_;
  assign _2697_ = load_i ? decrypt_i : round[3];
  assign _2698_ = _2690_ & round[2];
  assign _2699_ = _2698_ ^ round[3];
  assign _2700_ = _0000_ | round[2];
  assign _2701_ = _2700_ ^ _0022_;
  assign _2702_ = _2680_ ? round[3] : _2701_;
  assign _2703_ = _0469_ ? _2699_ : _2702_;
  assign _2704_ = subbytes_ready_o ? _2699_ : _2703_;
  assign _2705_ = _0468_ ? _2703_ : _2704_;
  assign _2706_ = _2705_ & _0462_;
  assign _2707_ = _2706_ | _2686_;
  assign next_round[3] = _0450_ ? _2697_ : _2707_;
  assign _2708_ = state & _2656_;
  assign _2709_ = _0462_ ? state : _2708_;
  assign next_state = _0450_ ? load_i : _2709_;
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[0] <= 0;
    else
      addroundkey_data_o[0] <= next_addroundkey_data_reg[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[100] <= 0;
    else
      addroundkey_data_o[100] <= next_addroundkey_data_reg[100];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[101] <= 0;
    else
      addroundkey_data_o[101] <= next_addroundkey_data_reg[101];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[102] <= 0;
    else
      addroundkey_data_o[102] <= next_addroundkey_data_reg[102];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[103] <= 0;
    else
      addroundkey_data_o[103] <= next_addroundkey_data_reg[103];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[104] <= 0;
    else
      addroundkey_data_o[104] <= next_addroundkey_data_reg[104];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[105] <= 0;
    else
      addroundkey_data_o[105] <= next_addroundkey_data_reg[105];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[106] <= 0;
    else
      addroundkey_data_o[106] <= next_addroundkey_data_reg[106];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[107] <= 0;
    else
      addroundkey_data_o[107] <= next_addroundkey_data_reg[107];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[108] <= 0;
    else
      addroundkey_data_o[108] <= next_addroundkey_data_reg[108];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[109] <= 0;
    else
      addroundkey_data_o[109] <= next_addroundkey_data_reg[109];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[10] <= 0;
    else
      addroundkey_data_o[10] <= next_addroundkey_data_reg[10];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[110] <= 0;
    else
      addroundkey_data_o[110] <= next_addroundkey_data_reg[110];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[111] <= 0;
    else
      addroundkey_data_o[111] <= next_addroundkey_data_reg[111];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[112] <= 0;
    else
      addroundkey_data_o[112] <= next_addroundkey_data_reg[112];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[113] <= 0;
    else
      addroundkey_data_o[113] <= next_addroundkey_data_reg[113];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[114] <= 0;
    else
      addroundkey_data_o[114] <= next_addroundkey_data_reg[114];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[115] <= 0;
    else
      addroundkey_data_o[115] <= next_addroundkey_data_reg[115];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[116] <= 0;
    else
      addroundkey_data_o[116] <= next_addroundkey_data_reg[116];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[117] <= 0;
    else
      addroundkey_data_o[117] <= next_addroundkey_data_reg[117];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[118] <= 0;
    else
      addroundkey_data_o[118] <= next_addroundkey_data_reg[118];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[119] <= 0;
    else
      addroundkey_data_o[119] <= next_addroundkey_data_reg[119];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[11] <= 0;
    else
      addroundkey_data_o[11] <= next_addroundkey_data_reg[11];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[120] <= 0;
    else
      addroundkey_data_o[120] <= next_addroundkey_data_reg[120];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[121] <= 0;
    else
      addroundkey_data_o[121] <= next_addroundkey_data_reg[121];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[122] <= 0;
    else
      addroundkey_data_o[122] <= next_addroundkey_data_reg[122];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[123] <= 0;
    else
      addroundkey_data_o[123] <= next_addroundkey_data_reg[123];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[124] <= 0;
    else
      addroundkey_data_o[124] <= next_addroundkey_data_reg[124];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[125] <= 0;
    else
      addroundkey_data_o[125] <= next_addroundkey_data_reg[125];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[126] <= 0;
    else
      addroundkey_data_o[126] <= next_addroundkey_data_reg[126];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[127] <= 0;
    else
      addroundkey_data_o[127] <= next_addroundkey_data_reg[127];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[12] <= 0;
    else
      addroundkey_data_o[12] <= next_addroundkey_data_reg[12];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[13] <= 0;
    else
      addroundkey_data_o[13] <= next_addroundkey_data_reg[13];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[14] <= 0;
    else
      addroundkey_data_o[14] <= next_addroundkey_data_reg[14];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[15] <= 0;
    else
      addroundkey_data_o[15] <= next_addroundkey_data_reg[15];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[16] <= 0;
    else
      addroundkey_data_o[16] <= next_addroundkey_data_reg[16];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[17] <= 0;
    else
      addroundkey_data_o[17] <= next_addroundkey_data_reg[17];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[18] <= 0;
    else
      addroundkey_data_o[18] <= next_addroundkey_data_reg[18];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[19] <= 0;
    else
      addroundkey_data_o[19] <= next_addroundkey_data_reg[19];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[1] <= 0;
    else
      addroundkey_data_o[1] <= next_addroundkey_data_reg[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[20] <= 0;
    else
      addroundkey_data_o[20] <= next_addroundkey_data_reg[20];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[21] <= 0;
    else
      addroundkey_data_o[21] <= next_addroundkey_data_reg[21];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[22] <= 0;
    else
      addroundkey_data_o[22] <= next_addroundkey_data_reg[22];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[23] <= 0;
    else
      addroundkey_data_o[23] <= next_addroundkey_data_reg[23];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[24] <= 0;
    else
      addroundkey_data_o[24] <= next_addroundkey_data_reg[24];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[25] <= 0;
    else
      addroundkey_data_o[25] <= next_addroundkey_data_reg[25];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[26] <= 0;
    else
      addroundkey_data_o[26] <= next_addroundkey_data_reg[26];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[27] <= 0;
    else
      addroundkey_data_o[27] <= next_addroundkey_data_reg[27];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[28] <= 0;
    else
      addroundkey_data_o[28] <= next_addroundkey_data_reg[28];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[29] <= 0;
    else
      addroundkey_data_o[29] <= next_addroundkey_data_reg[29];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[2] <= 0;
    else
      addroundkey_data_o[2] <= next_addroundkey_data_reg[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[30] <= 0;
    else
      addroundkey_data_o[30] <= next_addroundkey_data_reg[30];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[31] <= 0;
    else
      addroundkey_data_o[31] <= next_addroundkey_data_reg[31];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[32] <= 0;
    else
      addroundkey_data_o[32] <= next_addroundkey_data_reg[32];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[33] <= 0;
    else
      addroundkey_data_o[33] <= next_addroundkey_data_reg[33];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[34] <= 0;
    else
      addroundkey_data_o[34] <= next_addroundkey_data_reg[34];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[35] <= 0;
    else
      addroundkey_data_o[35] <= next_addroundkey_data_reg[35];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[36] <= 0;
    else
      addroundkey_data_o[36] <= next_addroundkey_data_reg[36];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[37] <= 0;
    else
      addroundkey_data_o[37] <= next_addroundkey_data_reg[37];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[38] <= 0;
    else
      addroundkey_data_o[38] <= next_addroundkey_data_reg[38];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[39] <= 0;
    else
      addroundkey_data_o[39] <= next_addroundkey_data_reg[39];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[3] <= 0;
    else
      addroundkey_data_o[3] <= next_addroundkey_data_reg[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[40] <= 0;
    else
      addroundkey_data_o[40] <= next_addroundkey_data_reg[40];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[41] <= 0;
    else
      addroundkey_data_o[41] <= next_addroundkey_data_reg[41];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[42] <= 0;
    else
      addroundkey_data_o[42] <= next_addroundkey_data_reg[42];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[43] <= 0;
    else
      addroundkey_data_o[43] <= next_addroundkey_data_reg[43];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[44] <= 0;
    else
      addroundkey_data_o[44] <= next_addroundkey_data_reg[44];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[45] <= 0;
    else
      addroundkey_data_o[45] <= next_addroundkey_data_reg[45];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[46] <= 0;
    else
      addroundkey_data_o[46] <= next_addroundkey_data_reg[46];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[47] <= 0;
    else
      addroundkey_data_o[47] <= next_addroundkey_data_reg[47];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[48] <= 0;
    else
      addroundkey_data_o[48] <= next_addroundkey_data_reg[48];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[49] <= 0;
    else
      addroundkey_data_o[49] <= next_addroundkey_data_reg[49];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[4] <= 0;
    else
      addroundkey_data_o[4] <= next_addroundkey_data_reg[4];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[50] <= 0;
    else
      addroundkey_data_o[50] <= next_addroundkey_data_reg[50];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[51] <= 0;
    else
      addroundkey_data_o[51] <= next_addroundkey_data_reg[51];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[52] <= 0;
    else
      addroundkey_data_o[52] <= next_addroundkey_data_reg[52];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[53] <= 0;
    else
      addroundkey_data_o[53] <= next_addroundkey_data_reg[53];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[54] <= 0;
    else
      addroundkey_data_o[54] <= next_addroundkey_data_reg[54];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[55] <= 0;
    else
      addroundkey_data_o[55] <= next_addroundkey_data_reg[55];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[56] <= 0;
    else
      addroundkey_data_o[56] <= next_addroundkey_data_reg[56];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[57] <= 0;
    else
      addroundkey_data_o[57] <= next_addroundkey_data_reg[57];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[58] <= 0;
    else
      addroundkey_data_o[58] <= next_addroundkey_data_reg[58];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[59] <= 0;
    else
      addroundkey_data_o[59] <= next_addroundkey_data_reg[59];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[5] <= 0;
    else
      addroundkey_data_o[5] <= next_addroundkey_data_reg[5];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[60] <= 0;
    else
      addroundkey_data_o[60] <= next_addroundkey_data_reg[60];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[61] <= 0;
    else
      addroundkey_data_o[61] <= next_addroundkey_data_reg[61];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[62] <= 0;
    else
      addroundkey_data_o[62] <= next_addroundkey_data_reg[62];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[63] <= 0;
    else
      addroundkey_data_o[63] <= next_addroundkey_data_reg[63];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[64] <= 0;
    else
      addroundkey_data_o[64] <= next_addroundkey_data_reg[64];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[65] <= 0;
    else
      addroundkey_data_o[65] <= next_addroundkey_data_reg[65];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[66] <= 0;
    else
      addroundkey_data_o[66] <= next_addroundkey_data_reg[66];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[67] <= 0;
    else
      addroundkey_data_o[67] <= next_addroundkey_data_reg[67];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[68] <= 0;
    else
      addroundkey_data_o[68] <= next_addroundkey_data_reg[68];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[69] <= 0;
    else
      addroundkey_data_o[69] <= next_addroundkey_data_reg[69];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[6] <= 0;
    else
      addroundkey_data_o[6] <= next_addroundkey_data_reg[6];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[70] <= 0;
    else
      addroundkey_data_o[70] <= next_addroundkey_data_reg[70];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[71] <= 0;
    else
      addroundkey_data_o[71] <= next_addroundkey_data_reg[71];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[72] <= 0;
    else
      addroundkey_data_o[72] <= next_addroundkey_data_reg[72];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[73] <= 0;
    else
      addroundkey_data_o[73] <= next_addroundkey_data_reg[73];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[74] <= 0;
    else
      addroundkey_data_o[74] <= next_addroundkey_data_reg[74];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[75] <= 0;
    else
      addroundkey_data_o[75] <= next_addroundkey_data_reg[75];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[76] <= 0;
    else
      addroundkey_data_o[76] <= next_addroundkey_data_reg[76];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[77] <= 0;
    else
      addroundkey_data_o[77] <= next_addroundkey_data_reg[77];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[78] <= 0;
    else
      addroundkey_data_o[78] <= next_addroundkey_data_reg[78];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[79] <= 0;
    else
      addroundkey_data_o[79] <= next_addroundkey_data_reg[79];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[7] <= 0;
    else
      addroundkey_data_o[7] <= next_addroundkey_data_reg[7];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[80] <= 0;
    else
      addroundkey_data_o[80] <= next_addroundkey_data_reg[80];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[81] <= 0;
    else
      addroundkey_data_o[81] <= next_addroundkey_data_reg[81];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[82] <= 0;
    else
      addroundkey_data_o[82] <= next_addroundkey_data_reg[82];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[83] <= 0;
    else
      addroundkey_data_o[83] <= next_addroundkey_data_reg[83];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[84] <= 0;
    else
      addroundkey_data_o[84] <= next_addroundkey_data_reg[84];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[85] <= 0;
    else
      addroundkey_data_o[85] <= next_addroundkey_data_reg[85];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[86] <= 0;
    else
      addroundkey_data_o[86] <= next_addroundkey_data_reg[86];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[87] <= 0;
    else
      addroundkey_data_o[87] <= next_addroundkey_data_reg[87];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[88] <= 0;
    else
      addroundkey_data_o[88] <= next_addroundkey_data_reg[88];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[89] <= 0;
    else
      addroundkey_data_o[89] <= next_addroundkey_data_reg[89];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[8] <= 0;
    else
      addroundkey_data_o[8] <= next_addroundkey_data_reg[8];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[90] <= 0;
    else
      addroundkey_data_o[90] <= next_addroundkey_data_reg[90];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[91] <= 0;
    else
      addroundkey_data_o[91] <= next_addroundkey_data_reg[91];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[92] <= 0;
    else
      addroundkey_data_o[92] <= next_addroundkey_data_reg[92];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[93] <= 0;
    else
      addroundkey_data_o[93] <= next_addroundkey_data_reg[93];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[94] <= 0;
    else
      addroundkey_data_o[94] <= next_addroundkey_data_reg[94];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[95] <= 0;
    else
      addroundkey_data_o[95] <= next_addroundkey_data_reg[95];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[96] <= 0;
    else
      addroundkey_data_o[96] <= next_addroundkey_data_reg[96];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[97] <= 0;
    else
      addroundkey_data_o[97] <= next_addroundkey_data_reg[97];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[98] <= 0;
    else
      addroundkey_data_o[98] <= next_addroundkey_data_reg[98];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[99] <= 0;
    else
      addroundkey_data_o[99] <= next_addroundkey_data_reg[99];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_data_o[9] <= 0;
    else
      addroundkey_data_o[9] <= next_addroundkey_data_reg[9];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_ready_o <= 0;
    else
      addroundkey_ready_o <= next_addroundkey_ready_o;
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_round[0] <= 0;
    else
      addroundkey_round[0] <= next_addroundkey_round[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_round[1] <= 0;
    else
      addroundkey_round[1] <= next_addroundkey_round[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_round[2] <= 0;
    else
      addroundkey_round[2] <= next_addroundkey_round[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_round[3] <= 0;
    else
      addroundkey_round[3] <= next_addroundkey_round[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      addroundkey_start_i <= 0;
    else
      addroundkey_start_i <= next_addroundkey_start_i;
  always @(posedge clk or negedge reset)
    if (!reset)
      first_round_reg <= 0;
    else
      first_round_reg <= next_first_round_reg;
  always @(posedge clk or negedge reset)
    if (!reset)
      ready_o <= 0;
    else
      ready_o <= next_ready_o;
  always @(posedge clk or negedge reset)
    if (!reset)
      round[0] <= 0;
    else
      round[0] <= next_round[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      round[1] <= 0;
    else
      round[1] <= next_round[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      round[2] <= 0;
    else
      round[2] <= next_round[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      round[3] <= 0;
    else
      round[3] <= next_round[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      state <= 0;
    else
      state <= next_state;
  keysched ks1 (
    .clk(clk),
    .last_key_i(keysched_last_key_i),
    .new_key_o(keysched_new_key_o),
    .ready_o(keysched_ready_o),
    .reset(reset),
    .round_i(keysched_round_i),
    .sbox_access_o(keysched_sbox_access_o),
    .sbox_data_i(sbox_data_o),
    .sbox_data_o(keysched_sbox_data_o),
    .sbox_decrypt_o(keysched_sbox_decrypt_o),
    .start_i(keysched_start_i)
  );
  mixcolum mix1 (
    .clk(clk),
    .data_i(mixcol_data_i),
    .data_o(mixcol_data_o),
    .decrypt_i(decrypt_i),
    .ready_o(mixcol_ready_o),
    .reset(reset),
    .start_i(mixcol_start_i)
  );
  sbox sbox1 (
    .clk(clk),
    .data_i(sbox_data_i),
    .data_o(sbox_data_o),
    .decrypt_i(sbox_decrypt_i),
    .reset(reset)
  );
  subbytes sub1 (
    .clk(clk),
    .data_i(subbytes_data_i),
    .data_o(subbytes_data_o),
    .decrypt_i(decrypt_i),
    .ready_o(subbytes_ready_o),
    .reset(reset),
    .sbox_data_i(sbox_data_o),
    .sbox_data_o(subbytes_sbox_data_o),
    .sbox_decrypt_o(subbytes_sbox_decrypt_o),
    .start_i(subbytes_start_i)
  );
  assign addroundkey_data_reg = addroundkey_data_o;
  assign data_o = addroundkey_data_o;
endmodule

module byte_mixcolum(a, b, c, d, outx, outy);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  input [7:0] a;
  input [7:0] b;
  input [7:0] c;
  input [7:0] d;
  output [7:0] outx;
  wire [7:0] outx_var;
  output [7:0] outy;
  assign _019_ = d[0] ^ c[0];
  assign _020_ = _019_ ^ b[0];
  assign _021_ = a[7] ^ b[7];
  assign outx[0] = _021_ ^ _020_;
  assign _022_ = d[1] ^ c[1];
  assign _023_ = _022_ ^ b[1];
  assign _024_ = a[0] ^ b[0];
  assign _025_ = _024_ ^ _021_;
  assign outx[1] = _025_ ^ _023_;
  assign _026_ = d[2] ^ c[2];
  assign _027_ = _026_ ^ b[2];
  assign _028_ = a[1] ^ b[1];
  assign outx[2] = _028_ ^ _027_;
  assign _029_ = d[3] ^ c[3];
  assign _030_ = _029_ ^ b[3];
  assign _031_ = a[2] ^ b[2];
  assign _032_ = _031_ ^ _021_;
  assign outx[3] = _032_ ^ _030_;
  assign _033_ = d[4] ^ c[4];
  assign _034_ = _033_ ^ b[4];
  assign _035_ = a[3] ^ b[3];
  assign _036_ = _035_ ^ _021_;
  assign outx[4] = _036_ ^ _034_;
  assign _037_ = d[5] ^ c[5];
  assign _038_ = _037_ ^ b[5];
  assign _039_ = a[4] ^ b[4];
  assign outx[5] = _039_ ^ _038_;
  assign _040_ = d[6] ^ c[6];
  assign _041_ = _040_ ^ b[6];
  assign _042_ = a[5] ^ b[5];
  assign outx[6] = _042_ ^ _041_;
  assign _043_ = d[7] ^ c[7];
  assign _044_ = _043_ ^ b[7];
  assign _045_ = a[6] ^ b[6];
  assign outx[7] = _045_ ^ _044_;
  assign _046_ = c[6] ^ a[6];
  assign _047_ = _046_ ^ _042_;
  assign _048_ = _047_ ^ _037_;
  assign outy[0] = _048_ ^ outx[0];
  assign _049_ = c[7] ^ a[7];
  assign _050_ = _049_ ^ _045_;
  assign _051_ = _050_ ^ _040_;
  assign _052_ = _051_ ^ _048_;
  assign outy[1] = _052_ ^ outx[1];
  assign _053_ = c[0] ^ a[0];
  assign _054_ = _053_ ^ _021_;
  assign _055_ = _054_ ^ _043_;
  assign _056_ = _055_ ^ _051_;
  assign outy[2] = _056_ ^ outx[2];
  assign _057_ = c[1] ^ a[1];
  assign _058_ = _057_ ^ _025_;
  assign _059_ = _043_ ^ _019_;
  assign _000_ = _059_ ^ _058_;
  assign _001_ = _000_ ^ _048_;
  assign outy[3] = _001_ ^ outx[3];
  assign _002_ = c[2] ^ a[2];
  assign _003_ = _002_ ^ _028_;
  assign _004_ = _003_ ^ _022_;
  assign _005_ = _004_ ^ _051_;
  assign _006_ = _005_ ^ _048_;
  assign outy[4] = _006_ ^ outx[4];
  assign _007_ = c[3] ^ a[3];
  assign _008_ = _007_ ^ _032_;
  assign _009_ = _043_ ^ _026_;
  assign _010_ = _009_ ^ _008_;
  assign _011_ = _010_ ^ _051_;
  assign outy[5] = _011_ ^ outx[5];
  assign _012_ = c[4] ^ a[4];
  assign _013_ = _012_ ^ _036_;
  assign _014_ = _043_ ^ _029_;
  assign _015_ = _014_ ^ _013_;
  assign outy[6] = _015_ ^ outx[6];
  assign _016_ = c[5] ^ a[5];
  assign _017_ = _016_ ^ _039_;
  assign _018_ = _017_ ^ _033_;
  assign outy[7] = _018_ ^ outx[7];
  assign outx_var = outx;
endmodule

module keysched(clk, reset, start_i, round_i, last_key_i, new_key_o, ready_o, sbox_access_o, sbox_data_o, sbox_data_i, sbox_decrypt_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire [127:0] K_var;
  input clk;
  reg [31:0] col;
  wire [31:0] col_t;
  reg [127:0] key_reg;
  input [127:0] last_key_i;
  output [127:0] new_key_o;
  wire [31:0] next_col;
  wire [127:0] next_key_reg;
  wire next_ready_o;
  wire [2:0] next_state;
  output ready_o;
  reg ready_o;
  input reset;
  input [3:0] round_i;
  output sbox_access_o;
  input [7:0] sbox_data_i;
  output [7:0] sbox_data_o;
  output sbox_decrypt_o;
  input start_i;
  reg [2:0] state;
  assign _0194_ = ~state[2];
  assign _0195_ = state[1] | state[0];
  assign _0196_ = _0195_ | _0194_;
  assign _0197_ = last_key_i[96] ^ col[0];
  assign _0198_ = _0197_ ^ last_key_i[64];
  assign _0199_ = _0198_ ^ last_key_i[32];
  assign _0200_ = _0199_ ^ last_key_i[0];
  assign next_key_reg[0] = _0196_ ? key_reg[0] : _0200_;
  assign _0201_ = last_key_i[100] ^ col[4];
  assign next_key_reg[100] = _0196_ ? key_reg[100] : _0201_;
  assign _0202_ = last_key_i[101] ^ col[5];
  assign next_key_reg[101] = _0196_ ? key_reg[101] : _0202_;
  assign _0203_ = last_key_i[102] ^ col[6];
  assign next_key_reg[102] = _0196_ ? key_reg[102] : _0203_;
  assign _0204_ = last_key_i[103] ^ col[7];
  assign next_key_reg[103] = _0196_ ? key_reg[103] : _0204_;
  assign _0205_ = ~col[8];
  assign _0206_ = _0195_ | state[2];
  assign _0207_ = _0205_ | start_i;
  assign _0208_ = _0207_ | _0206_;
  assign _0209_ = ~sbox_data_i[0];
  assign _0210_ = _0196_ | _0209_;
  assign _0211_ = _0210_ & _0208_;
  assign _0212_ = _0195_ ? _0205_ : _0211_;
  assign _0213_ = _0212_ ^ last_key_i[104];
  assign _0214_ = ~_0213_;
  assign next_key_reg[104] = _0196_ ? key_reg[104] : _0214_;
  assign _0215_ = ~col[9];
  assign _0216_ = _0215_ | start_i;
  assign _0217_ = _0216_ | _0206_;
  assign _0218_ = ~sbox_data_i[1];
  assign _0219_ = _0196_ | _0218_;
  assign _0220_ = _0219_ & _0217_;
  assign _0221_ = _0195_ ? _0215_ : _0220_;
  assign _0222_ = _0221_ ^ last_key_i[105];
  assign _0223_ = ~_0222_;
  assign next_key_reg[105] = _0196_ ? key_reg[105] : _0223_;
  assign _0224_ = ~col[10];
  assign _0225_ = _0224_ | start_i;
  assign _0226_ = _0225_ | _0206_;
  assign _0227_ = ~sbox_data_i[2];
  assign _0228_ = _0196_ | _0227_;
  assign _0229_ = _0228_ & _0226_;
  assign _0230_ = _0195_ ? _0224_ : _0229_;
  assign _0231_ = _0230_ ^ last_key_i[106];
  assign _0232_ = ~_0231_;
  assign next_key_reg[106] = _0196_ ? key_reg[106] : _0232_;
  assign _0233_ = ~col[11];
  assign _0234_ = _0233_ | start_i;
  assign _0235_ = _0234_ | _0206_;
  assign _0236_ = ~sbox_data_i[3];
  assign _0237_ = _0196_ | _0236_;
  assign _0238_ = _0237_ & _0235_;
  assign _0239_ = _0195_ ? _0233_ : _0238_;
  assign _0240_ = _0239_ ^ last_key_i[107];
  assign _0241_ = ~_0240_;
  assign next_key_reg[107] = _0196_ ? key_reg[107] : _0241_;
  assign _0242_ = ~col[12];
  assign _0243_ = _0242_ | start_i;
  assign _0244_ = _0243_ | _0206_;
  assign _0245_ = ~sbox_data_i[4];
  assign _0246_ = _0196_ | _0245_;
  assign _0247_ = _0246_ & _0244_;
  assign _0248_ = _0195_ ? _0242_ : _0247_;
  assign _0249_ = _0248_ ^ last_key_i[108];
  assign _0250_ = ~_0249_;
  assign next_key_reg[108] = _0196_ ? key_reg[108] : _0250_;
  assign _0251_ = ~col[13];
  assign _0252_ = _0251_ | start_i;
  assign _0253_ = _0252_ | _0206_;
  assign _0254_ = ~sbox_data_i[5];
  assign _0255_ = _0196_ | _0254_;
  assign _0256_ = _0255_ & _0253_;
  assign _0257_ = _0195_ ? _0251_ : _0256_;
  assign _0258_ = _0257_ ^ last_key_i[109];
  assign _0259_ = ~_0258_;
  assign next_key_reg[109] = _0196_ ? key_reg[109] : _0259_;
  assign _0260_ = _0231_ ^ last_key_i[74];
  assign _0261_ = ~_0260_;
  assign _0262_ = _0261_ ^ last_key_i[42];
  assign _0263_ = _0262_ ^ last_key_i[10];
  assign next_key_reg[10] = _0196_ ? key_reg[10] : _0263_;
  assign _0264_ = ~col[14];
  assign _0265_ = _0264_ | start_i;
  assign _0266_ = _0265_ | _0206_;
  assign _0267_ = ~sbox_data_i[6];
  assign _0268_ = _0196_ | _0267_;
  assign _0269_ = _0268_ & _0266_;
  assign _0270_ = _0195_ ? _0264_ : _0269_;
  assign _0271_ = _0270_ ^ last_key_i[110];
  assign _0272_ = ~_0271_;
  assign next_key_reg[110] = _0196_ ? key_reg[110] : _0272_;
  assign _0273_ = ~col[15];
  assign _0274_ = _0273_ | start_i;
  assign _0275_ = _0274_ | _0206_;
  assign _0276_ = ~sbox_data_i[7];
  assign _0277_ = _0196_ | _0276_;
  assign _0278_ = _0277_ & _0275_;
  assign _0279_ = _0195_ ? _0273_ : _0278_;
  assign _0280_ = _0279_ ^ last_key_i[111];
  assign _0281_ = ~_0280_;
  assign next_key_reg[111] = _0196_ ? key_reg[111] : _0281_;
  assign _0282_ = last_key_i[112] ^ col[16];
  assign next_key_reg[112] = _0196_ ? key_reg[112] : _0282_;
  assign _0283_ = last_key_i[113] ^ col[17];
  assign next_key_reg[113] = _0196_ ? key_reg[113] : _0283_;
  assign _0284_ = last_key_i[114] ^ col[18];
  assign next_key_reg[114] = _0196_ ? key_reg[114] : _0284_;
  assign _0285_ = last_key_i[115] ^ col[19];
  assign next_key_reg[115] = _0196_ ? key_reg[115] : _0285_;
  assign _0286_ = last_key_i[116] ^ col[20];
  assign next_key_reg[116] = _0196_ ? key_reg[116] : _0286_;
  assign _0287_ = last_key_i[117] ^ col[21];
  assign next_key_reg[117] = _0196_ ? key_reg[117] : _0287_;
  assign _0288_ = last_key_i[118] ^ col[22];
  assign next_key_reg[118] = _0196_ ? key_reg[118] : _0288_;
  assign _0289_ = last_key_i[119] ^ col[23];
  assign next_key_reg[119] = _0196_ ? key_reg[119] : _0289_;
  assign _0290_ = _0240_ ^ last_key_i[75];
  assign _0291_ = ~_0290_;
  assign _0292_ = _0291_ ^ last_key_i[43];
  assign _0293_ = _0292_ ^ last_key_i[11];
  assign next_key_reg[11] = _0196_ ? key_reg[11] : _0293_;
  assign _0294_ = last_key_i[120] ^ col[24];
  assign _0295_ = ~round_i[3];
  assign _0296_ = ~round_i[2];
  assign _0297_ = ~round_i[0];
  assign _0298_ = round_i[1] & _0297_;
  assign _0299_ = _0298_ & _0296_;
  assign _0300_ = _0299_ & _0295_;
  assign _0301_ = ~round_i[1];
  assign _0302_ = _0301_ & round_i[0];
  assign _0303_ = _0302_ & _0296_;
  assign _0304_ = round_i[1] & round_i[0];
  assign _0305_ = _0295_ & _0296_;
  assign _0306_ = _0305_ & _0304_;
  assign _0307_ = _0301_ & _0297_;
  assign _0308_ = _0295_ & round_i[2];
  assign _0309_ = _0308_ & _0307_;
  assign _0310_ = _0303_ & round_i[3];
  assign _0311_ = _0299_ & round_i[3];
  assign _0312_ = _0311_ | _0310_;
  assign _0313_ = _0308_ & _0302_;
  assign _0314_ = _0308_ & _0298_;
  assign _0315_ = _0308_ & _0304_;
  assign _0316_ = round_i[3] & _0296_;
  assign _0317_ = _0316_ & _0307_;
  assign _0318_ = _0303_ ^ _0294_;
  assign next_key_reg[120] = _0196_ ? key_reg[120] : _0318_;
  assign _0319_ = last_key_i[121] ^ col[25];
  assign _0320_ = _0312_ | _0300_;
  assign _0321_ = _0320_ ^ _0319_;
  assign next_key_reg[121] = _0196_ ? key_reg[121] : _0321_;
  assign _0322_ = last_key_i[122] ^ col[26];
  assign _0323_ = _0311_ | _0306_;
  assign _0324_ = _0323_ ^ _0322_;
  assign next_key_reg[122] = _0196_ ? key_reg[122] : _0324_;
  assign _0325_ = last_key_i[123] ^ col[27];
  assign _0326_ = _0310_ | _0309_;
  assign _0327_ = _0326_ ^ _0325_;
  assign next_key_reg[123] = _0196_ ? key_reg[123] : _0327_;
  assign _0328_ = last_key_i[124] ^ col[28];
  assign _0329_ = _0313_ | _0312_;
  assign _0330_ = _0329_ ^ _0328_;
  assign next_key_reg[124] = _0196_ ? key_reg[124] : _0330_;
  assign _0331_ = last_key_i[125] ^ col[29];
  assign _0332_ = _0314_ | _0311_;
  assign _0333_ = _0332_ ^ _0331_;
  assign next_key_reg[125] = _0196_ ? key_reg[125] : _0333_;
  assign _0334_ = last_key_i[126] ^ col[30];
  assign _0335_ = _0315_ ^ _0334_;
  assign next_key_reg[126] = _0196_ ? key_reg[126] : _0335_;
  assign _0336_ = last_key_i[127] ^ col[31];
  assign _0337_ = _0317_ ^ _0336_;
  assign next_key_reg[127] = _0196_ ? key_reg[127] : _0337_;
  assign _0338_ = _0249_ ^ last_key_i[76];
  assign _0339_ = ~_0338_;
  assign _0340_ = _0339_ ^ last_key_i[44];
  assign _0341_ = _0340_ ^ last_key_i[12];
  assign next_key_reg[12] = _0196_ ? key_reg[12] : _0341_;
  assign _0342_ = _0258_ ^ last_key_i[77];
  assign _0343_ = ~_0342_;
  assign _0344_ = _0343_ ^ last_key_i[45];
  assign _0345_ = _0344_ ^ last_key_i[13];
  assign next_key_reg[13] = _0196_ ? key_reg[13] : _0345_;
  assign _0346_ = _0271_ ^ last_key_i[78];
  assign _0347_ = ~_0346_;
  assign _0348_ = _0347_ ^ last_key_i[46];
  assign _0349_ = _0348_ ^ last_key_i[14];
  assign next_key_reg[14] = _0196_ ? key_reg[14] : _0349_;
  assign _0350_ = _0280_ ^ last_key_i[79];
  assign _0351_ = ~_0350_;
  assign _0352_ = _0351_ ^ last_key_i[47];
  assign _0353_ = _0352_ ^ last_key_i[15];
  assign next_key_reg[15] = _0196_ ? key_reg[15] : _0353_;
  assign _0354_ = _0282_ ^ last_key_i[80];
  assign _0355_ = _0354_ ^ last_key_i[48];
  assign _0356_ = _0355_ ^ last_key_i[16];
  assign next_key_reg[16] = _0196_ ? key_reg[16] : _0356_;
  assign _0357_ = _0283_ ^ last_key_i[81];
  assign _0358_ = _0357_ ^ last_key_i[49];
  assign _0359_ = _0358_ ^ last_key_i[17];
  assign next_key_reg[17] = _0196_ ? key_reg[17] : _0359_;
  assign _0360_ = _0284_ ^ last_key_i[82];
  assign _0361_ = _0360_ ^ last_key_i[50];
  assign _0362_ = _0361_ ^ last_key_i[18];
  assign next_key_reg[18] = _0196_ ? key_reg[18] : _0362_;
  assign _0363_ = _0285_ ^ last_key_i[83];
  assign _0364_ = _0363_ ^ last_key_i[51];
  assign _0365_ = _0364_ ^ last_key_i[19];
  assign next_key_reg[19] = _0196_ ? key_reg[19] : _0365_;
  assign _0366_ = last_key_i[97] ^ col[1];
  assign _0367_ = _0366_ ^ last_key_i[65];
  assign _0368_ = _0367_ ^ last_key_i[33];
  assign _0369_ = _0368_ ^ last_key_i[1];
  assign next_key_reg[1] = _0196_ ? key_reg[1] : _0369_;
  assign _0370_ = _0286_ ^ last_key_i[84];
  assign _0371_ = _0370_ ^ last_key_i[52];
  assign _0372_ = _0371_ ^ last_key_i[20];
  assign next_key_reg[20] = _0196_ ? key_reg[20] : _0372_;
  assign _0373_ = _0287_ ^ last_key_i[85];
  assign _0374_ = _0373_ ^ last_key_i[53];
  assign _0375_ = _0374_ ^ last_key_i[21];
  assign next_key_reg[21] = _0196_ ? key_reg[21] : _0375_;
  assign _0376_ = _0288_ ^ last_key_i[86];
  assign _0377_ = _0376_ ^ last_key_i[54];
  assign _0378_ = _0377_ ^ last_key_i[22];
  assign next_key_reg[22] = _0196_ ? key_reg[22] : _0378_;
  assign _0379_ = _0289_ ^ last_key_i[87];
  assign _0380_ = _0379_ ^ last_key_i[55];
  assign _0381_ = _0380_ ^ last_key_i[23];
  assign next_key_reg[23] = _0196_ ? key_reg[23] : _0381_;
  assign _0382_ = _0318_ ^ last_key_i[88];
  assign _0383_ = _0382_ ^ last_key_i[56];
  assign _0384_ = _0383_ ^ last_key_i[24];
  assign next_key_reg[24] = _0196_ ? key_reg[24] : _0384_;
  assign _0385_ = _0321_ ^ last_key_i[89];
  assign _0386_ = _0385_ ^ last_key_i[57];
  assign _0387_ = _0386_ ^ last_key_i[25];
  assign next_key_reg[25] = _0196_ ? key_reg[25] : _0387_;
  assign _0388_ = _0324_ ^ last_key_i[90];
  assign _0389_ = _0388_ ^ last_key_i[58];
  assign _0390_ = _0389_ ^ last_key_i[26];
  assign next_key_reg[26] = _0196_ ? key_reg[26] : _0390_;
  assign _0391_ = _0327_ ^ last_key_i[91];
  assign _0392_ = _0391_ ^ last_key_i[59];
  assign _0393_ = _0392_ ^ last_key_i[27];
  assign next_key_reg[27] = _0196_ ? key_reg[27] : _0393_;
  assign _0394_ = _0330_ ^ last_key_i[92];
  assign _0395_ = _0394_ ^ last_key_i[60];
  assign _0396_ = _0395_ ^ last_key_i[28];
  assign next_key_reg[28] = _0196_ ? key_reg[28] : _0396_;
  assign _0397_ = _0333_ ^ last_key_i[93];
  assign _0398_ = _0397_ ^ last_key_i[61];
  assign _0399_ = _0398_ ^ last_key_i[29];
  assign next_key_reg[29] = _0196_ ? key_reg[29] : _0399_;
  assign _0400_ = last_key_i[98] ^ col[2];
  assign _0401_ = _0400_ ^ last_key_i[66];
  assign _0402_ = _0401_ ^ last_key_i[34];
  assign _0403_ = _0402_ ^ last_key_i[2];
  assign next_key_reg[2] = _0196_ ? key_reg[2] : _0403_;
  assign _0404_ = _0335_ ^ last_key_i[94];
  assign _0405_ = _0404_ ^ last_key_i[62];
  assign _0406_ = _0405_ ^ last_key_i[30];
  assign next_key_reg[30] = _0196_ ? key_reg[30] : _0406_;
  assign _0407_ = _0337_ ^ last_key_i[95];
  assign _0408_ = _0407_ ^ last_key_i[63];
  assign _0409_ = _0408_ ^ last_key_i[31];
  assign next_key_reg[31] = _0196_ ? key_reg[31] : _0409_;
  assign next_key_reg[32] = _0196_ ? key_reg[32] : _0199_;
  assign next_key_reg[33] = _0196_ ? key_reg[33] : _0368_;
  assign next_key_reg[34] = _0196_ ? key_reg[34] : _0402_;
  assign _0410_ = last_key_i[99] ^ col[3];
  assign _0411_ = _0410_ ^ last_key_i[67];
  assign _0412_ = _0411_ ^ last_key_i[35];
  assign next_key_reg[35] = _0196_ ? key_reg[35] : _0412_;
  assign _0413_ = _0201_ ^ last_key_i[68];
  assign _0414_ = _0413_ ^ last_key_i[36];
  assign next_key_reg[36] = _0196_ ? key_reg[36] : _0414_;
  assign _0415_ = _0202_ ^ last_key_i[69];
  assign _0416_ = _0415_ ^ last_key_i[37];
  assign next_key_reg[37] = _0196_ ? key_reg[37] : _0416_;
  assign _0417_ = _0203_ ^ last_key_i[70];
  assign _0418_ = _0417_ ^ last_key_i[38];
  assign next_key_reg[38] = _0196_ ? key_reg[38] : _0418_;
  assign _0419_ = _0204_ ^ last_key_i[71];
  assign _0420_ = _0419_ ^ last_key_i[39];
  assign next_key_reg[39] = _0196_ ? key_reg[39] : _0420_;
  assign _0421_ = _0412_ ^ last_key_i[3];
  assign next_key_reg[3] = _0196_ ? key_reg[3] : _0421_;
  assign _0422_ = _0213_ ^ last_key_i[72];
  assign _0423_ = ~_0422_;
  assign _0424_ = _0423_ ^ last_key_i[40];
  assign next_key_reg[40] = _0196_ ? key_reg[40] : _0424_;
  assign _0425_ = _0222_ ^ last_key_i[73];
  assign _0426_ = ~_0425_;
  assign _0427_ = _0426_ ^ last_key_i[41];
  assign next_key_reg[41] = _0196_ ? key_reg[41] : _0427_;
  assign next_key_reg[42] = _0196_ ? key_reg[42] : _0262_;
  assign next_key_reg[43] = _0196_ ? key_reg[43] : _0292_;
  assign next_key_reg[44] = _0196_ ? key_reg[44] : _0340_;
  assign next_key_reg[45] = _0196_ ? key_reg[45] : _0344_;
  assign next_key_reg[46] = _0196_ ? key_reg[46] : _0348_;
  assign next_key_reg[47] = _0196_ ? key_reg[47] : _0352_;
  assign next_key_reg[48] = _0196_ ? key_reg[48] : _0355_;
  assign next_key_reg[49] = _0196_ ? key_reg[49] : _0358_;
  assign _0428_ = _0414_ ^ last_key_i[4];
  assign next_key_reg[4] = _0196_ ? key_reg[4] : _0428_;
  assign next_key_reg[50] = _0196_ ? key_reg[50] : _0361_;
  assign next_key_reg[51] = _0196_ ? key_reg[51] : _0364_;
  assign next_key_reg[52] = _0196_ ? key_reg[52] : _0371_;
  assign next_key_reg[53] = _0196_ ? key_reg[53] : _0374_;
  assign next_key_reg[54] = _0196_ ? key_reg[54] : _0377_;
  assign next_key_reg[55] = _0196_ ? key_reg[55] : _0380_;
  assign next_key_reg[56] = _0196_ ? key_reg[56] : _0383_;
  assign next_key_reg[57] = _0196_ ? key_reg[57] : _0386_;
  assign next_key_reg[58] = _0196_ ? key_reg[58] : _0389_;
  assign next_key_reg[59] = _0196_ ? key_reg[59] : _0392_;
  assign _0429_ = _0416_ ^ last_key_i[5];
  assign next_key_reg[5] = _0196_ ? key_reg[5] : _0429_;
  assign next_key_reg[60] = _0196_ ? key_reg[60] : _0395_;
  assign next_key_reg[61] = _0196_ ? key_reg[61] : _0398_;
  assign next_key_reg[62] = _0196_ ? key_reg[62] : _0405_;
  assign next_key_reg[63] = _0196_ ? key_reg[63] : _0408_;
  assign next_key_reg[64] = _0196_ ? key_reg[64] : _0198_;
  assign next_key_reg[65] = _0196_ ? key_reg[65] : _0367_;
  assign next_key_reg[66] = _0196_ ? key_reg[66] : _0401_;
  assign next_key_reg[67] = _0196_ ? key_reg[67] : _0411_;
  assign next_key_reg[68] = _0196_ ? key_reg[68] : _0413_;
  assign next_key_reg[69] = _0196_ ? key_reg[69] : _0415_;
  assign _0430_ = _0418_ ^ last_key_i[6];
  assign next_key_reg[6] = _0196_ ? key_reg[6] : _0430_;
  assign next_key_reg[70] = _0196_ ? key_reg[70] : _0417_;
  assign next_key_reg[71] = _0196_ ? key_reg[71] : _0419_;
  assign next_key_reg[72] = _0196_ ? key_reg[72] : _0423_;
  assign next_key_reg[73] = _0196_ ? key_reg[73] : _0426_;
  assign next_key_reg[74] = _0196_ ? key_reg[74] : _0261_;
  assign next_key_reg[75] = _0196_ ? key_reg[75] : _0291_;
  assign next_key_reg[76] = _0196_ ? key_reg[76] : _0339_;
  assign next_key_reg[77] = _0196_ ? key_reg[77] : _0343_;
  assign next_key_reg[78] = _0196_ ? key_reg[78] : _0347_;
  assign next_key_reg[79] = _0196_ ? key_reg[79] : _0351_;
  assign _0431_ = _0420_ ^ last_key_i[7];
  assign next_key_reg[7] = _0196_ ? key_reg[7] : _0431_;
  assign next_key_reg[80] = _0196_ ? key_reg[80] : _0354_;
  assign next_key_reg[81] = _0196_ ? key_reg[81] : _0357_;
  assign next_key_reg[82] = _0196_ ? key_reg[82] : _0360_;
  assign next_key_reg[83] = _0196_ ? key_reg[83] : _0363_;
  assign next_key_reg[84] = _0196_ ? key_reg[84] : _0370_;
  assign next_key_reg[85] = _0196_ ? key_reg[85] : _0373_;
  assign next_key_reg[86] = _0196_ ? key_reg[86] : _0376_;
  assign next_key_reg[87] = _0196_ ? key_reg[87] : _0379_;
  assign next_key_reg[88] = _0196_ ? key_reg[88] : _0382_;
  assign next_key_reg[89] = _0196_ ? key_reg[89] : _0385_;
  assign _0432_ = _0424_ ^ last_key_i[8];
  assign next_key_reg[8] = _0196_ ? key_reg[8] : _0432_;
  assign next_key_reg[90] = _0196_ ? key_reg[90] : _0388_;
  assign next_key_reg[91] = _0196_ ? key_reg[91] : _0391_;
  assign next_key_reg[92] = _0196_ ? key_reg[92] : _0394_;
  assign next_key_reg[93] = _0196_ ? key_reg[93] : _0397_;
  assign next_key_reg[94] = _0196_ ? key_reg[94] : _0404_;
  assign next_key_reg[95] = _0196_ ? key_reg[95] : _0407_;
  assign next_key_reg[96] = _0196_ ? key_reg[96] : _0197_;
  assign next_key_reg[97] = _0196_ ? key_reg[97] : _0366_;
  assign next_key_reg[98] = _0196_ ? key_reg[98] : _0400_;
  assign next_key_reg[99] = _0196_ ? key_reg[99] : _0410_;
  assign _0433_ = _0427_ ^ last_key_i[9];
  assign next_key_reg[9] = _0196_ ? key_reg[9] : _0433_;
  assign next_ready_o = ~_0196_;
  assign _0434_ = ~state[1];
  assign _0435_ = _0434_ & state[0];
  assign _0436_ = _0435_ & _0194_;
  assign _0437_ = _0436_ | next_ready_o;
  assign _0438_ = ~state[0];
  assign _0439_ = state[1] & _0438_;
  assign _0440_ = _0439_ & _0194_;
  assign _0441_ = state[1] & state[0];
  assign _0442_ = _0441_ & _0194_;
  assign _0443_ = _0442_ | _0440_;
  assign _0444_ = _0443_ | _0437_;
  assign _0445_ = ~_0444_;
  assign _0446_ = _0436_ & sbox_data_i[0];
  assign _0447_ = _0440_ & col[0];
  assign _0448_ = _0447_ | _0446_;
  assign _0449_ = _0442_ & col[0];
  assign _0450_ = next_ready_o & col[0];
  assign _0451_ = _0450_ | _0449_;
  assign _0452_ = _0451_ | _0448_;
  assign next_col[0] = _0445_ ? col[0] : _0452_;
  assign _0453_ = ~_0230_;
  assign _0454_ = _0453_ & next_ready_o;
  assign _0455_ = _0442_ & col[10];
  assign _0456_ = _0436_ & col[10];
  assign _0457_ = _0440_ & col[10];
  assign _0458_ = _0457_ | _0456_;
  assign _0459_ = _0458_ | _0455_;
  assign _0460_ = _0459_ | _0454_;
  assign next_col[10] = _0445_ ? col[10] : _0460_;
  assign _0461_ = ~_0239_;
  assign _0462_ = _0461_ & next_ready_o;
  assign _0463_ = _0442_ & col[11];
  assign _0464_ = _0436_ & col[11];
  assign _0465_ = _0440_ & col[11];
  assign _0466_ = _0465_ | _0464_;
  assign _0467_ = _0466_ | _0463_;
  assign _0468_ = _0467_ | _0462_;
  assign next_col[11] = _0445_ ? col[11] : _0468_;
  assign _0469_ = ~_0248_;
  assign _0470_ = _0469_ & next_ready_o;
  assign _0471_ = _0442_ & col[12];
  assign _0472_ = _0436_ & col[12];
  assign _0473_ = _0440_ & col[12];
  assign _0474_ = _0473_ | _0472_;
  assign _0475_ = _0474_ | _0471_;
  assign _0476_ = _0475_ | _0470_;
  assign next_col[12] = _0445_ ? col[12] : _0476_;
  assign _0477_ = ~_0257_;
  assign _0478_ = _0477_ & next_ready_o;
  assign _0479_ = _0442_ & col[13];
  assign _0480_ = _0436_ & col[13];
  assign _0481_ = _0440_ & col[13];
  assign _0482_ = _0481_ | _0480_;
  assign _0483_ = _0482_ | _0479_;
  assign _0484_ = _0483_ | _0478_;
  assign next_col[13] = _0445_ ? col[13] : _0484_;
  assign _0485_ = ~_0270_;
  assign _0486_ = _0485_ & next_ready_o;
  assign _0487_ = _0442_ & col[14];
  assign _0488_ = _0436_ & col[14];
  assign _0489_ = _0440_ & col[14];
  assign _0490_ = _0489_ | _0488_;
  assign _0491_ = _0490_ | _0487_;
  assign _0492_ = _0491_ | _0486_;
  assign next_col[14] = _0445_ ? col[14] : _0492_;
  assign _0493_ = ~_0279_;
  assign _0494_ = _0493_ & next_ready_o;
  assign _0495_ = _0442_ & col[15];
  assign _0496_ = _0436_ & col[15];
  assign _0497_ = _0440_ & col[15];
  assign _0498_ = _0497_ | _0496_;
  assign _0499_ = _0498_ | _0495_;
  assign _0500_ = _0499_ | _0494_;
  assign next_col[15] = _0445_ ? col[15] : _0500_;
  assign _0501_ = _0436_ & col[16];
  assign _0502_ = _0440_ & col[16];
  assign _0503_ = _0502_ | _0501_;
  assign _0504_ = _0442_ & sbox_data_i[0];
  assign _0505_ = next_ready_o & col[16];
  assign _0506_ = _0505_ | _0504_;
  assign _0507_ = _0506_ | _0503_;
  assign next_col[16] = _0445_ ? col[16] : _0507_;
  assign _0508_ = _0436_ & col[17];
  assign _0509_ = _0440_ & col[17];
  assign _0510_ = _0509_ | _0508_;
  assign _0511_ = _0442_ & sbox_data_i[1];
  assign _0512_ = next_ready_o & col[17];
  assign _0513_ = _0512_ | _0511_;
  assign _0514_ = _0513_ | _0510_;
  assign next_col[17] = _0445_ ? col[17] : _0514_;
  assign _0515_ = _0436_ & col[18];
  assign _0516_ = _0440_ & col[18];
  assign _0517_ = _0516_ | _0515_;
  assign _0518_ = _0442_ & sbox_data_i[2];
  assign _0519_ = next_ready_o & col[18];
  assign _0520_ = _0519_ | _0518_;
  assign _0521_ = _0520_ | _0517_;
  assign next_col[18] = _0445_ ? col[18] : _0521_;
  assign _0522_ = _0436_ & col[19];
  assign _0523_ = _0440_ & col[19];
  assign _0524_ = _0523_ | _0522_;
  assign _0525_ = _0442_ & sbox_data_i[3];
  assign _0526_ = next_ready_o & col[19];
  assign _0527_ = _0526_ | _0525_;
  assign _0528_ = _0527_ | _0524_;
  assign next_col[19] = _0445_ ? col[19] : _0528_;
  assign _0529_ = _0436_ & sbox_data_i[1];
  assign _0530_ = _0440_ & col[1];
  assign _0531_ = _0530_ | _0529_;
  assign _0532_ = _0442_ & col[1];
  assign _0533_ = next_ready_o & col[1];
  assign _0534_ = _0533_ | _0532_;
  assign _0535_ = _0534_ | _0531_;
  assign next_col[1] = _0445_ ? col[1] : _0535_;
  assign _0536_ = _0436_ & col[20];
  assign _0537_ = _0440_ & col[20];
  assign _0538_ = _0537_ | _0536_;
  assign _0539_ = _0442_ & sbox_data_i[4];
  assign _0540_ = next_ready_o & col[20];
  assign _0541_ = _0540_ | _0539_;
  assign _0542_ = _0541_ | _0538_;
  assign next_col[20] = _0445_ ? col[20] : _0542_;
  assign _0543_ = _0436_ & col[21];
  assign _0544_ = _0440_ & col[21];
  assign _0545_ = _0544_ | _0543_;
  assign _0546_ = _0442_ & sbox_data_i[5];
  assign _0547_ = next_ready_o & col[21];
  assign _0548_ = _0547_ | _0546_;
  assign _0549_ = _0548_ | _0545_;
  assign next_col[21] = _0445_ ? col[21] : _0549_;
  assign _0550_ = _0436_ & col[22];
  assign _0551_ = _0440_ & col[22];
  assign _0552_ = _0551_ | _0550_;
  assign _0553_ = _0442_ & sbox_data_i[6];
  assign _0554_ = next_ready_o & col[22];
  assign _0000_ = _0554_ | _0553_;
  assign _0001_ = _0000_ | _0552_;
  assign next_col[22] = _0445_ ? col[22] : _0001_;
  assign _0002_ = _0436_ & col[23];
  assign _0003_ = _0440_ & col[23];
  assign _0004_ = _0003_ | _0002_;
  assign _0005_ = _0442_ & sbox_data_i[7];
  assign _0006_ = next_ready_o & col[23];
  assign _0007_ = _0006_ | _0005_;
  assign _0008_ = _0007_ | _0004_;
  assign next_col[23] = _0445_ ? col[23] : _0008_;
  assign _0009_ = _0436_ & col[24];
  assign _0010_ = _0440_ & sbox_data_i[0];
  assign _0011_ = _0010_ | _0009_;
  assign _0012_ = _0442_ & col[24];
  assign _0013_ = next_ready_o & col[24];
  assign _0014_ = _0013_ | _0012_;
  assign _0015_ = _0014_ | _0011_;
  assign next_col[24] = _0445_ ? col[24] : _0015_;
  assign _0016_ = _0436_ & col[25];
  assign _0017_ = _0440_ & sbox_data_i[1];
  assign _0018_ = _0017_ | _0016_;
  assign _0019_ = _0442_ & col[25];
  assign _0020_ = next_ready_o & col[25];
  assign _0021_ = _0020_ | _0019_;
  assign _0022_ = _0021_ | _0018_;
  assign next_col[25] = _0445_ ? col[25] : _0022_;
  assign _0023_ = _0436_ & col[26];
  assign _0024_ = _0440_ & sbox_data_i[2];
  assign _0025_ = _0024_ | _0023_;
  assign _0026_ = _0442_ & col[26];
  assign _0027_ = next_ready_o & col[26];
  assign _0028_ = _0027_ | _0026_;
  assign _0029_ = _0028_ | _0025_;
  assign next_col[26] = _0445_ ? col[26] : _0029_;
  assign _0030_ = _0436_ & col[27];
  assign _0031_ = _0440_ & sbox_data_i[3];
  assign _0032_ = _0031_ | _0030_;
  assign _0033_ = _0442_ & col[27];
  assign _0034_ = next_ready_o & col[27];
  assign _0035_ = _0034_ | _0033_;
  assign _0036_ = _0035_ | _0032_;
  assign next_col[27] = _0445_ ? col[27] : _0036_;
  assign _0037_ = _0436_ & col[28];
  assign _0038_ = _0440_ & sbox_data_i[4];
  assign _0039_ = _0038_ | _0037_;
  assign _0040_ = _0442_ & col[28];
  assign _0041_ = next_ready_o & col[28];
  assign _0042_ = _0041_ | _0040_;
  assign _0043_ = _0042_ | _0039_;
  assign next_col[28] = _0445_ ? col[28] : _0043_;
  assign _0044_ = _0436_ & col[29];
  assign _0045_ = _0440_ & sbox_data_i[5];
  assign _0046_ = _0045_ | _0044_;
  assign _0047_ = _0442_ & col[29];
  assign _0048_ = next_ready_o & col[29];
  assign _0049_ = _0048_ | _0047_;
  assign _0050_ = _0049_ | _0046_;
  assign next_col[29] = _0445_ ? col[29] : _0050_;
  assign _0051_ = _0436_ & sbox_data_i[2];
  assign _0052_ = _0440_ & col[2];
  assign _0053_ = _0052_ | _0051_;
  assign _0054_ = _0442_ & col[2];
  assign _0055_ = next_ready_o & col[2];
  assign _0056_ = _0055_ | _0054_;
  assign _0057_ = _0056_ | _0053_;
  assign next_col[2] = _0445_ ? col[2] : _0057_;
  assign _0058_ = _0436_ & col[30];
  assign _0059_ = _0440_ & sbox_data_i[6];
  assign _0060_ = _0059_ | _0058_;
  assign _0061_ = _0442_ & col[30];
  assign _0062_ = next_ready_o & col[30];
  assign _0063_ = _0062_ | _0061_;
  assign _0064_ = _0063_ | _0060_;
  assign next_col[30] = _0445_ ? col[30] : _0064_;
  assign _0065_ = _0436_ & col[31];
  assign _0066_ = _0440_ & sbox_data_i[7];
  assign _0067_ = _0066_ | _0065_;
  assign _0068_ = _0442_ & col[31];
  assign _0069_ = next_ready_o & col[31];
  assign _0070_ = _0069_ | _0068_;
  assign _0071_ = _0070_ | _0067_;
  assign next_col[31] = _0445_ ? col[31] : _0071_;
  assign _0072_ = _0436_ & sbox_data_i[3];
  assign _0073_ = _0440_ & col[3];
  assign _0074_ = _0073_ | _0072_;
  assign _0075_ = _0442_ & col[3];
  assign _0076_ = next_ready_o & col[3];
  assign _0077_ = _0076_ | _0075_;
  assign _0078_ = _0077_ | _0074_;
  assign next_col[3] = _0445_ ? col[3] : _0078_;
  assign _0079_ = _0436_ & sbox_data_i[4];
  assign _0080_ = _0440_ & col[4];
  assign _0081_ = _0080_ | _0079_;
  assign _0082_ = _0442_ & col[4];
  assign _0083_ = next_ready_o & col[4];
  assign _0084_ = _0083_ | _0082_;
  assign _0085_ = _0084_ | _0081_;
  assign next_col[4] = _0445_ ? col[4] : _0085_;
  assign _0086_ = _0436_ & sbox_data_i[5];
  assign _0087_ = _0440_ & col[5];
  assign _0088_ = _0087_ | _0086_;
  assign _0089_ = _0442_ & col[5];
  assign _0090_ = next_ready_o & col[5];
  assign _0091_ = _0090_ | _0089_;
  assign _0092_ = _0091_ | _0088_;
  assign next_col[5] = _0445_ ? col[5] : _0092_;
  assign _0093_ = _0436_ & sbox_data_i[6];
  assign _0094_ = _0440_ & col[6];
  assign _0095_ = _0094_ | _0093_;
  assign _0096_ = _0442_ & col[6];
  assign _0097_ = next_ready_o & col[6];
  assign _0098_ = _0097_ | _0096_;
  assign _0099_ = _0098_ | _0095_;
  assign next_col[6] = _0445_ ? col[6] : _0099_;
  assign _0100_ = _0436_ & sbox_data_i[7];
  assign _0101_ = _0440_ & col[7];
  assign _0102_ = _0101_ | _0100_;
  assign _0103_ = _0442_ & col[7];
  assign _0104_ = next_ready_o & col[7];
  assign _0105_ = _0104_ | _0103_;
  assign _0106_ = _0105_ | _0102_;
  assign next_col[7] = _0445_ ? col[7] : _0106_;
  assign _0107_ = ~_0212_;
  assign _0108_ = _0107_ & next_ready_o;
  assign _0109_ = _0442_ & col[8];
  assign _0110_ = _0436_ & col[8];
  assign _0111_ = _0440_ & col[8];
  assign _0112_ = _0111_ | _0110_;
  assign _0113_ = _0112_ | _0109_;
  assign _0114_ = _0113_ | _0108_;
  assign next_col[8] = _0445_ ? col[8] : _0114_;
  assign _0115_ = ~_0221_;
  assign _0116_ = _0115_ & next_ready_o;
  assign _0117_ = _0442_ & col[9];
  assign _0118_ = _0436_ & col[9];
  assign _0119_ = _0440_ & col[9];
  assign _0120_ = _0119_ | _0118_;
  assign _0121_ = _0120_ | _0117_;
  assign _0122_ = _0121_ | _0116_;
  assign next_col[9] = _0445_ ? col[9] : _0122_;
  assign _0123_ = ~_0206_;
  assign _0124_ = state[0] | start_i;
  assign _0125_ = _0124_ & _0123_;
  assign _0126_ = _0125_ | _0440_;
  assign next_state[0] = _0126_ & _0194_;
  assign _0127_ = _0440_ | _0436_;
  assign next_state[1] = _0127_ & _0194_;
  assign next_state[2] = _0442_ & _0194_;
  assign _0128_ = _0444_ | _0123_;
  assign _0129_ = _0125_ | _0444_;
  assign sbox_access_o = _0129_ & _0128_;
  assign _0130_ = last_key_i[24] & start_i;
  assign _0131_ = _0130_ & _0123_;
  assign _0132_ = _0436_ & last_key_i[16];
  assign _0133_ = _0132_ | _0131_;
  assign _0134_ = _0440_ & last_key_i[8];
  assign _0135_ = _0442_ & last_key_i[0];
  assign _0136_ = _0135_ | _0134_;
  assign _0137_ = _0136_ | _0133_;
  assign sbox_data_o[0] = _0137_ & _0194_;
  assign _0138_ = last_key_i[25] & start_i;
  assign _0139_ = _0138_ & _0123_;
  assign _0140_ = _0436_ & last_key_i[17];
  assign _0141_ = _0140_ | _0139_;
  assign _0142_ = _0440_ & last_key_i[9];
  assign _0143_ = _0442_ & last_key_i[1];
  assign _0144_ = _0143_ | _0142_;
  assign _0145_ = _0144_ | _0141_;
  assign sbox_data_o[1] = _0145_ & _0194_;
  assign _0146_ = last_key_i[26] & start_i;
  assign _0147_ = _0146_ & _0123_;
  assign _0148_ = _0436_ & last_key_i[18];
  assign _0149_ = _0148_ | _0147_;
  assign _0150_ = _0440_ & last_key_i[10];
  assign _0151_ = _0442_ & last_key_i[2];
  assign _0152_ = _0151_ | _0150_;
  assign _0153_ = _0152_ | _0149_;
  assign sbox_data_o[2] = _0153_ & _0194_;
  assign _0154_ = last_key_i[27] & start_i;
  assign _0155_ = _0154_ & _0123_;
  assign _0156_ = _0436_ & last_key_i[19];
  assign _0157_ = _0156_ | _0155_;
  assign _0158_ = _0440_ & last_key_i[11];
  assign _0159_ = _0442_ & last_key_i[3];
  assign _0160_ = _0159_ | _0158_;
  assign _0161_ = _0160_ | _0157_;
  assign sbox_data_o[3] = _0161_ & _0194_;
  assign _0162_ = last_key_i[28] & start_i;
  assign _0163_ = _0162_ & _0123_;
  assign _0164_ = _0436_ & last_key_i[20];
  assign _0165_ = _0164_ | _0163_;
  assign _0166_ = _0440_ & last_key_i[12];
  assign _0167_ = _0442_ & last_key_i[4];
  assign _0168_ = _0167_ | _0166_;
  assign _0169_ = _0168_ | _0165_;
  assign sbox_data_o[4] = _0169_ & _0194_;
  assign _0170_ = last_key_i[29] & start_i;
  assign _0171_ = _0170_ & _0123_;
  assign _0172_ = _0436_ & last_key_i[21];
  assign _0173_ = _0172_ | _0171_;
  assign _0174_ = _0440_ & last_key_i[13];
  assign _0175_ = _0442_ & last_key_i[5];
  assign _0176_ = _0175_ | _0174_;
  assign _0177_ = _0176_ | _0173_;
  assign sbox_data_o[5] = _0177_ & _0194_;
  assign _0178_ = last_key_i[30] & start_i;
  assign _0179_ = _0178_ & _0123_;
  assign _0180_ = _0436_ & last_key_i[22];
  assign _0181_ = _0180_ | _0179_;
  assign _0182_ = _0440_ & last_key_i[14];
  assign _0183_ = _0442_ & last_key_i[6];
  assign _0184_ = _0183_ | _0182_;
  assign _0185_ = _0184_ | _0181_;
  assign sbox_data_o[6] = _0185_ & _0194_;
  assign _0186_ = last_key_i[31] & start_i;
  assign _0187_ = _0186_ & _0123_;
  assign _0188_ = _0436_ & last_key_i[23];
  assign _0189_ = _0188_ | _0187_;
  assign _0190_ = _0440_ & last_key_i[15];
  assign _0191_ = _0442_ & last_key_i[7];
  assign _0192_ = _0191_ | _0190_;
  assign _0193_ = _0192_ | _0189_;
  assign sbox_data_o[7] = _0193_ & _0194_;
  always @(posedge clk or negedge reset)
    if (!reset)
      col[0] <= 0;
    else
      col[0] <= next_col[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[10] <= 0;
    else
      col[10] <= next_col[10];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[11] <= 0;
    else
      col[11] <= next_col[11];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[12] <= 0;
    else
      col[12] <= next_col[12];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[13] <= 0;
    else
      col[13] <= next_col[13];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[14] <= 0;
    else
      col[14] <= next_col[14];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[15] <= 0;
    else
      col[15] <= next_col[15];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[16] <= 0;
    else
      col[16] <= next_col[16];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[17] <= 0;
    else
      col[17] <= next_col[17];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[18] <= 0;
    else
      col[18] <= next_col[18];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[19] <= 0;
    else
      col[19] <= next_col[19];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[1] <= 0;
    else
      col[1] <= next_col[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[20] <= 0;
    else
      col[20] <= next_col[20];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[21] <= 0;
    else
      col[21] <= next_col[21];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[22] <= 0;
    else
      col[22] <= next_col[22];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[23] <= 0;
    else
      col[23] <= next_col[23];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[24] <= 0;
    else
      col[24] <= next_col[24];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[25] <= 0;
    else
      col[25] <= next_col[25];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[26] <= 0;
    else
      col[26] <= next_col[26];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[27] <= 0;
    else
      col[27] <= next_col[27];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[28] <= 0;
    else
      col[28] <= next_col[28];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[29] <= 0;
    else
      col[29] <= next_col[29];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[2] <= 0;
    else
      col[2] <= next_col[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[30] <= 0;
    else
      col[30] <= next_col[30];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[31] <= 0;
    else
      col[31] <= next_col[31];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[3] <= 0;
    else
      col[3] <= next_col[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[4] <= 0;
    else
      col[4] <= next_col[4];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[5] <= 0;
    else
      col[5] <= next_col[5];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[6] <= 0;
    else
      col[6] <= next_col[6];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[7] <= 0;
    else
      col[7] <= next_col[7];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[8] <= 0;
    else
      col[8] <= next_col[8];
  always @(posedge clk or negedge reset)
    if (!reset)
      col[9] <= 0;
    else
      col[9] <= next_col[9];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[0] <= 0;
    else
      key_reg[0] <= next_key_reg[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[100] <= 0;
    else
      key_reg[100] <= next_key_reg[100];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[101] <= 0;
    else
      key_reg[101] <= next_key_reg[101];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[102] <= 0;
    else
      key_reg[102] <= next_key_reg[102];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[103] <= 0;
    else
      key_reg[103] <= next_key_reg[103];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[104] <= 0;
    else
      key_reg[104] <= next_key_reg[104];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[105] <= 0;
    else
      key_reg[105] <= next_key_reg[105];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[106] <= 0;
    else
      key_reg[106] <= next_key_reg[106];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[107] <= 0;
    else
      key_reg[107] <= next_key_reg[107];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[108] <= 0;
    else
      key_reg[108] <= next_key_reg[108];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[109] <= 0;
    else
      key_reg[109] <= next_key_reg[109];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[10] <= 0;
    else
      key_reg[10] <= next_key_reg[10];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[110] <= 0;
    else
      key_reg[110] <= next_key_reg[110];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[111] <= 0;
    else
      key_reg[111] <= next_key_reg[111];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[112] <= 0;
    else
      key_reg[112] <= next_key_reg[112];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[113] <= 0;
    else
      key_reg[113] <= next_key_reg[113];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[114] <= 0;
    else
      key_reg[114] <= next_key_reg[114];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[115] <= 0;
    else
      key_reg[115] <= next_key_reg[115];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[116] <= 0;
    else
      key_reg[116] <= next_key_reg[116];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[117] <= 0;
    else
      key_reg[117] <= next_key_reg[117];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[118] <= 0;
    else
      key_reg[118] <= next_key_reg[118];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[119] <= 0;
    else
      key_reg[119] <= next_key_reg[119];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[11] <= 0;
    else
      key_reg[11] <= next_key_reg[11];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[120] <= 0;
    else
      key_reg[120] <= next_key_reg[120];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[121] <= 0;
    else
      key_reg[121] <= next_key_reg[121];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[122] <= 0;
    else
      key_reg[122] <= next_key_reg[122];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[123] <= 0;
    else
      key_reg[123] <= next_key_reg[123];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[124] <= 0;
    else
      key_reg[124] <= next_key_reg[124];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[125] <= 0;
    else
      key_reg[125] <= next_key_reg[125];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[126] <= 0;
    else
      key_reg[126] <= next_key_reg[126];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[127] <= 0;
    else
      key_reg[127] <= next_key_reg[127];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[12] <= 0;
    else
      key_reg[12] <= next_key_reg[12];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[13] <= 0;
    else
      key_reg[13] <= next_key_reg[13];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[14] <= 0;
    else
      key_reg[14] <= next_key_reg[14];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[15] <= 0;
    else
      key_reg[15] <= next_key_reg[15];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[16] <= 0;
    else
      key_reg[16] <= next_key_reg[16];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[17] <= 0;
    else
      key_reg[17] <= next_key_reg[17];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[18] <= 0;
    else
      key_reg[18] <= next_key_reg[18];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[19] <= 0;
    else
      key_reg[19] <= next_key_reg[19];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[1] <= 0;
    else
      key_reg[1] <= next_key_reg[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[20] <= 0;
    else
      key_reg[20] <= next_key_reg[20];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[21] <= 0;
    else
      key_reg[21] <= next_key_reg[21];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[22] <= 0;
    else
      key_reg[22] <= next_key_reg[22];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[23] <= 0;
    else
      key_reg[23] <= next_key_reg[23];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[24] <= 0;
    else
      key_reg[24] <= next_key_reg[24];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[25] <= 0;
    else
      key_reg[25] <= next_key_reg[25];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[26] <= 0;
    else
      key_reg[26] <= next_key_reg[26];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[27] <= 0;
    else
      key_reg[27] <= next_key_reg[27];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[28] <= 0;
    else
      key_reg[28] <= next_key_reg[28];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[29] <= 0;
    else
      key_reg[29] <= next_key_reg[29];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[2] <= 0;
    else
      key_reg[2] <= next_key_reg[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[30] <= 0;
    else
      key_reg[30] <= next_key_reg[30];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[31] <= 0;
    else
      key_reg[31] <= next_key_reg[31];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[32] <= 0;
    else
      key_reg[32] <= next_key_reg[32];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[33] <= 0;
    else
      key_reg[33] <= next_key_reg[33];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[34] <= 0;
    else
      key_reg[34] <= next_key_reg[34];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[35] <= 0;
    else
      key_reg[35] <= next_key_reg[35];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[36] <= 0;
    else
      key_reg[36] <= next_key_reg[36];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[37] <= 0;
    else
      key_reg[37] <= next_key_reg[37];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[38] <= 0;
    else
      key_reg[38] <= next_key_reg[38];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[39] <= 0;
    else
      key_reg[39] <= next_key_reg[39];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[3] <= 0;
    else
      key_reg[3] <= next_key_reg[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[40] <= 0;
    else
      key_reg[40] <= next_key_reg[40];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[41] <= 0;
    else
      key_reg[41] <= next_key_reg[41];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[42] <= 0;
    else
      key_reg[42] <= next_key_reg[42];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[43] <= 0;
    else
      key_reg[43] <= next_key_reg[43];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[44] <= 0;
    else
      key_reg[44] <= next_key_reg[44];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[45] <= 0;
    else
      key_reg[45] <= next_key_reg[45];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[46] <= 0;
    else
      key_reg[46] <= next_key_reg[46];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[47] <= 0;
    else
      key_reg[47] <= next_key_reg[47];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[48] <= 0;
    else
      key_reg[48] <= next_key_reg[48];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[49] <= 0;
    else
      key_reg[49] <= next_key_reg[49];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[4] <= 0;
    else
      key_reg[4] <= next_key_reg[4];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[50] <= 0;
    else
      key_reg[50] <= next_key_reg[50];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[51] <= 0;
    else
      key_reg[51] <= next_key_reg[51];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[52] <= 0;
    else
      key_reg[52] <= next_key_reg[52];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[53] <= 0;
    else
      key_reg[53] <= next_key_reg[53];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[54] <= 0;
    else
      key_reg[54] <= next_key_reg[54];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[55] <= 0;
    else
      key_reg[55] <= next_key_reg[55];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[56] <= 0;
    else
      key_reg[56] <= next_key_reg[56];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[57] <= 0;
    else
      key_reg[57] <= next_key_reg[57];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[58] <= 0;
    else
      key_reg[58] <= next_key_reg[58];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[59] <= 0;
    else
      key_reg[59] <= next_key_reg[59];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[5] <= 0;
    else
      key_reg[5] <= next_key_reg[5];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[60] <= 0;
    else
      key_reg[60] <= next_key_reg[60];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[61] <= 0;
    else
      key_reg[61] <= next_key_reg[61];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[62] <= 0;
    else
      key_reg[62] <= next_key_reg[62];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[63] <= 0;
    else
      key_reg[63] <= next_key_reg[63];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[64] <= 0;
    else
      key_reg[64] <= next_key_reg[64];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[65] <= 0;
    else
      key_reg[65] <= next_key_reg[65];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[66] <= 0;
    else
      key_reg[66] <= next_key_reg[66];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[67] <= 0;
    else
      key_reg[67] <= next_key_reg[67];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[68] <= 0;
    else
      key_reg[68] <= next_key_reg[68];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[69] <= 0;
    else
      key_reg[69] <= next_key_reg[69];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[6] <= 0;
    else
      key_reg[6] <= next_key_reg[6];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[70] <= 0;
    else
      key_reg[70] <= next_key_reg[70];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[71] <= 0;
    else
      key_reg[71] <= next_key_reg[71];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[72] <= 0;
    else
      key_reg[72] <= next_key_reg[72];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[73] <= 0;
    else
      key_reg[73] <= next_key_reg[73];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[74] <= 0;
    else
      key_reg[74] <= next_key_reg[74];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[75] <= 0;
    else
      key_reg[75] <= next_key_reg[75];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[76] <= 0;
    else
      key_reg[76] <= next_key_reg[76];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[77] <= 0;
    else
      key_reg[77] <= next_key_reg[77];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[78] <= 0;
    else
      key_reg[78] <= next_key_reg[78];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[79] <= 0;
    else
      key_reg[79] <= next_key_reg[79];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[7] <= 0;
    else
      key_reg[7] <= next_key_reg[7];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[80] <= 0;
    else
      key_reg[80] <= next_key_reg[80];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[81] <= 0;
    else
      key_reg[81] <= next_key_reg[81];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[82] <= 0;
    else
      key_reg[82] <= next_key_reg[82];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[83] <= 0;
    else
      key_reg[83] <= next_key_reg[83];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[84] <= 0;
    else
      key_reg[84] <= next_key_reg[84];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[85] <= 0;
    else
      key_reg[85] <= next_key_reg[85];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[86] <= 0;
    else
      key_reg[86] <= next_key_reg[86];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[87] <= 0;
    else
      key_reg[87] <= next_key_reg[87];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[88] <= 0;
    else
      key_reg[88] <= next_key_reg[88];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[89] <= 0;
    else
      key_reg[89] <= next_key_reg[89];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[8] <= 0;
    else
      key_reg[8] <= next_key_reg[8];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[90] <= 0;
    else
      key_reg[90] <= next_key_reg[90];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[91] <= 0;
    else
      key_reg[91] <= next_key_reg[91];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[92] <= 0;
    else
      key_reg[92] <= next_key_reg[92];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[93] <= 0;
    else
      key_reg[93] <= next_key_reg[93];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[94] <= 0;
    else
      key_reg[94] <= next_key_reg[94];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[95] <= 0;
    else
      key_reg[95] <= next_key_reg[95];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[96] <= 0;
    else
      key_reg[96] <= next_key_reg[96];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[97] <= 0;
    else
      key_reg[97] <= next_key_reg[97];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[98] <= 0;
    else
      key_reg[98] <= next_key_reg[98];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[99] <= 0;
    else
      key_reg[99] <= next_key_reg[99];
  always @(posedge clk or negedge reset)
    if (!reset)
      key_reg[9] <= 0;
    else
      key_reg[9] <= next_key_reg[9];
  always @(posedge clk or negedge reset)
    if (!reset)
      ready_o <= 0;
    else
      ready_o <= next_ready_o;
  always @(posedge clk or negedge reset)
    if (!reset)
      state[0] <= 0;
    else
      state[0] <= next_state[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[1] <= 0;
    else
      state[1] <= next_state[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[2] <= 0;
    else
      state[2] <= next_state[2];
  assign K_var = last_key_i;
  assign { col_t[23:16], col_t[7:0] } = { sbox_data_i, sbox_data_i };
  assign new_key_o = key_reg;
  assign sbox_decrypt_o = 1'b0;
endmodule

module mixcolum(clk, reset, decrypt_i, start_i, data_i, ready_o, data_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  input clk;
  input [127:0] data_i;
  wire [127:0] data_i_var;
  output [127:0] data_o;
  reg [127:0] data_o;
  wire [127:0] data_o_reg;
  wire [127:0] data_reg;
  input decrypt_i;
  wire [31:0] mix_word;
  wire [127:0] next_data_o;
  wire [127:0] next_data_reg;
  wire next_ready_o;
  wire [1:0] next_state;
  wire [31:0] outx;
  wire [31:0] outy;
  output ready_o;
  reg ready_o;
  input reset;
  input start_i;
  reg [1:0] state;
  assign next_ready_o = state[1] & state[0];
  assign _0512_ = decrypt_i ? outy[0] : outx[0];
  assign next_data_o[0] = next_ready_o ? _0512_ : data_o[0];
  assign next_data_o[100] = next_ready_o ? data_reg[100] : data_o[100];
  assign next_data_o[101] = next_ready_o ? data_reg[101] : data_o[101];
  assign next_data_o[102] = next_ready_o ? data_reg[102] : data_o[102];
  assign next_data_o[103] = next_ready_o ? data_reg[103] : data_o[103];
  assign next_data_o[104] = next_ready_o ? data_reg[104] : data_o[104];
  assign next_data_o[105] = next_ready_o ? data_reg[105] : data_o[105];
  assign next_data_o[106] = next_ready_o ? data_reg[106] : data_o[106];
  assign next_data_o[107] = next_ready_o ? data_reg[107] : data_o[107];
  assign next_data_o[108] = next_ready_o ? data_reg[108] : data_o[108];
  assign next_data_o[109] = next_ready_o ? data_reg[109] : data_o[109];
  assign _0513_ = decrypt_i ? outy[10] : outx[10];
  assign next_data_o[10] = next_ready_o ? _0513_ : data_o[10];
  assign next_data_o[110] = next_ready_o ? data_reg[110] : data_o[110];
  assign next_data_o[111] = next_ready_o ? data_reg[111] : data_o[111];
  assign next_data_o[112] = next_ready_o ? data_reg[112] : data_o[112];
  assign next_data_o[113] = next_ready_o ? data_reg[113] : data_o[113];
  assign next_data_o[114] = next_ready_o ? data_reg[114] : data_o[114];
  assign next_data_o[115] = next_ready_o ? data_reg[115] : data_o[115];
  assign next_data_o[116] = next_ready_o ? data_reg[116] : data_o[116];
  assign next_data_o[117] = next_ready_o ? data_reg[117] : data_o[117];
  assign next_data_o[118] = next_ready_o ? data_reg[118] : data_o[118];
  assign next_data_o[119] = next_ready_o ? data_reg[119] : data_o[119];
  assign _0514_ = decrypt_i ? outy[11] : outx[11];
  assign next_data_o[11] = next_ready_o ? _0514_ : data_o[11];
  assign next_data_o[120] = next_ready_o ? data_reg[120] : data_o[120];
  assign next_data_o[121] = next_ready_o ? data_reg[121] : data_o[121];
  assign next_data_o[122] = next_ready_o ? data_reg[122] : data_o[122];
  assign next_data_o[123] = next_ready_o ? data_reg[123] : data_o[123];
  assign next_data_o[124] = next_ready_o ? data_reg[124] : data_o[124];
  assign next_data_o[125] = next_ready_o ? data_reg[125] : data_o[125];
  assign next_data_o[126] = next_ready_o ? data_reg[126] : data_o[126];
  assign next_data_o[127] = next_ready_o ? data_reg[127] : data_o[127];
  assign _0515_ = decrypt_i ? outy[12] : outx[12];
  assign next_data_o[12] = next_ready_o ? _0515_ : data_o[12];
  assign _0516_ = decrypt_i ? outy[13] : outx[13];
  assign next_data_o[13] = next_ready_o ? _0516_ : data_o[13];
  assign _0517_ = decrypt_i ? outy[14] : outx[14];
  assign next_data_o[14] = next_ready_o ? _0517_ : data_o[14];
  assign _0518_ = decrypt_i ? outy[15] : outx[15];
  assign next_data_o[15] = next_ready_o ? _0518_ : data_o[15];
  assign _0519_ = decrypt_i ? outy[16] : outx[16];
  assign next_data_o[16] = next_ready_o ? _0519_ : data_o[16];
  assign _0520_ = decrypt_i ? outy[17] : outx[17];
  assign next_data_o[17] = next_ready_o ? _0520_ : data_o[17];
  assign _0521_ = decrypt_i ? outy[18] : outx[18];
  assign next_data_o[18] = next_ready_o ? _0521_ : data_o[18];
  assign _0522_ = decrypt_i ? outy[19] : outx[19];
  assign next_data_o[19] = next_ready_o ? _0522_ : data_o[19];
  assign _0523_ = decrypt_i ? outy[1] : outx[1];
  assign next_data_o[1] = next_ready_o ? _0523_ : data_o[1];
  assign _0524_ = decrypt_i ? outy[20] : outx[20];
  assign next_data_o[20] = next_ready_o ? _0524_ : data_o[20];
  assign _0525_ = decrypt_i ? outy[21] : outx[21];
  assign next_data_o[21] = next_ready_o ? _0525_ : data_o[21];
  assign _0526_ = decrypt_i ? outy[22] : outx[22];
  assign next_data_o[22] = next_ready_o ? _0526_ : data_o[22];
  assign _0527_ = decrypt_i ? outy[23] : outx[23];
  assign next_data_o[23] = next_ready_o ? _0527_ : data_o[23];
  assign _0528_ = decrypt_i ? outy[24] : outx[24];
  assign next_data_o[24] = next_ready_o ? _0528_ : data_o[24];
  assign _0529_ = decrypt_i ? outy[25] : outx[25];
  assign next_data_o[25] = next_ready_o ? _0529_ : data_o[25];
  assign _0530_ = decrypt_i ? outy[26] : outx[26];
  assign next_data_o[26] = next_ready_o ? _0530_ : data_o[26];
  assign _0531_ = decrypt_i ? outy[27] : outx[27];
  assign next_data_o[27] = next_ready_o ? _0531_ : data_o[27];
  assign _0532_ = decrypt_i ? outy[28] : outx[28];
  assign next_data_o[28] = next_ready_o ? _0532_ : data_o[28];
  assign _0533_ = decrypt_i ? outy[29] : outx[29];
  assign next_data_o[29] = next_ready_o ? _0533_ : data_o[29];
  assign _0534_ = decrypt_i ? outy[2] : outx[2];
  assign next_data_o[2] = next_ready_o ? _0534_ : data_o[2];
  assign _0535_ = decrypt_i ? outy[30] : outx[30];
  assign next_data_o[30] = next_ready_o ? _0535_ : data_o[30];
  assign _0536_ = decrypt_i ? outy[31] : outx[31];
  assign next_data_o[31] = next_ready_o ? _0536_ : data_o[31];
  assign next_data_o[32] = next_ready_o ? data_reg[32] : data_o[32];
  assign next_data_o[33] = next_ready_o ? data_reg[33] : data_o[33];
  assign next_data_o[34] = next_ready_o ? data_reg[34] : data_o[34];
  assign next_data_o[35] = next_ready_o ? data_reg[35] : data_o[35];
  assign next_data_o[36] = next_ready_o ? data_reg[36] : data_o[36];
  assign next_data_o[37] = next_ready_o ? data_reg[37] : data_o[37];
  assign next_data_o[38] = next_ready_o ? data_reg[38] : data_o[38];
  assign next_data_o[39] = next_ready_o ? data_reg[39] : data_o[39];
  assign _0537_ = decrypt_i ? outy[3] : outx[3];
  assign next_data_o[3] = next_ready_o ? _0537_ : data_o[3];
  assign next_data_o[40] = next_ready_o ? data_reg[40] : data_o[40];
  assign next_data_o[41] = next_ready_o ? data_reg[41] : data_o[41];
  assign next_data_o[42] = next_ready_o ? data_reg[42] : data_o[42];
  assign next_data_o[43] = next_ready_o ? data_reg[43] : data_o[43];
  assign next_data_o[44] = next_ready_o ? data_reg[44] : data_o[44];
  assign next_data_o[45] = next_ready_o ? data_reg[45] : data_o[45];
  assign next_data_o[46] = next_ready_o ? data_reg[46] : data_o[46];
  assign next_data_o[47] = next_ready_o ? data_reg[47] : data_o[47];
  assign next_data_o[48] = next_ready_o ? data_reg[48] : data_o[48];
  assign next_data_o[49] = next_ready_o ? data_reg[49] : data_o[49];
  assign _0538_ = decrypt_i ? outy[4] : outx[4];
  assign next_data_o[4] = next_ready_o ? _0538_ : data_o[4];
  assign next_data_o[50] = next_ready_o ? data_reg[50] : data_o[50];
  assign next_data_o[51] = next_ready_o ? data_reg[51] : data_o[51];
  assign next_data_o[52] = next_ready_o ? data_reg[52] : data_o[52];
  assign next_data_o[53] = next_ready_o ? data_reg[53] : data_o[53];
  assign next_data_o[54] = next_ready_o ? data_reg[54] : data_o[54];
  assign next_data_o[55] = next_ready_o ? data_reg[55] : data_o[55];
  assign next_data_o[56] = next_ready_o ? data_reg[56] : data_o[56];
  assign next_data_o[57] = next_ready_o ? data_reg[57] : data_o[57];
  assign next_data_o[58] = next_ready_o ? data_reg[58] : data_o[58];
  assign next_data_o[59] = next_ready_o ? data_reg[59] : data_o[59];
  assign _0539_ = decrypt_i ? outy[5] : outx[5];
  assign next_data_o[5] = next_ready_o ? _0539_ : data_o[5];
  assign next_data_o[60] = next_ready_o ? data_reg[60] : data_o[60];
  assign next_data_o[61] = next_ready_o ? data_reg[61] : data_o[61];
  assign next_data_o[62] = next_ready_o ? data_reg[62] : data_o[62];
  assign next_data_o[63] = next_ready_o ? data_reg[63] : data_o[63];
  assign next_data_o[64] = next_ready_o ? data_reg[64] : data_o[64];
  assign next_data_o[65] = next_ready_o ? data_reg[65] : data_o[65];
  assign next_data_o[66] = next_ready_o ? data_reg[66] : data_o[66];
  assign next_data_o[67] = next_ready_o ? data_reg[67] : data_o[67];
  assign next_data_o[68] = next_ready_o ? data_reg[68] : data_o[68];
  assign next_data_o[69] = next_ready_o ? data_reg[69] : data_o[69];
  assign _0540_ = decrypt_i ? outy[6] : outx[6];
  assign next_data_o[6] = next_ready_o ? _0540_ : data_o[6];
  assign next_data_o[70] = next_ready_o ? data_reg[70] : data_o[70];
  assign next_data_o[71] = next_ready_o ? data_reg[71] : data_o[71];
  assign next_data_o[72] = next_ready_o ? data_reg[72] : data_o[72];
  assign next_data_o[73] = next_ready_o ? data_reg[73] : data_o[73];
  assign next_data_o[74] = next_ready_o ? data_reg[74] : data_o[74];
  assign next_data_o[75] = next_ready_o ? data_reg[75] : data_o[75];
  assign next_data_o[76] = next_ready_o ? data_reg[76] : data_o[76];
  assign next_data_o[77] = next_ready_o ? data_reg[77] : data_o[77];
  assign next_data_o[78] = next_ready_o ? data_reg[78] : data_o[78];
  assign next_data_o[79] = next_ready_o ? data_reg[79] : data_o[79];
  assign _0541_ = decrypt_i ? outy[7] : outx[7];
  assign next_data_o[7] = next_ready_o ? _0541_ : data_o[7];
  assign next_data_o[80] = next_ready_o ? data_reg[80] : data_o[80];
  assign next_data_o[81] = next_ready_o ? data_reg[81] : data_o[81];
  assign next_data_o[82] = next_ready_o ? data_reg[82] : data_o[82];
  assign next_data_o[83] = next_ready_o ? data_reg[83] : data_o[83];
  assign next_data_o[84] = next_ready_o ? data_reg[84] : data_o[84];
  assign next_data_o[85] = next_ready_o ? data_reg[85] : data_o[85];
  assign next_data_o[86] = next_ready_o ? data_reg[86] : data_o[86];
  assign next_data_o[87] = next_ready_o ? data_reg[87] : data_o[87];
  assign next_data_o[88] = next_ready_o ? data_reg[88] : data_o[88];
  assign next_data_o[89] = next_ready_o ? data_reg[89] : data_o[89];
  assign _0542_ = decrypt_i ? outy[8] : outx[8];
  assign next_data_o[8] = next_ready_o ? _0542_ : data_o[8];
  assign next_data_o[90] = next_ready_o ? data_reg[90] : data_o[90];
  assign next_data_o[91] = next_ready_o ? data_reg[91] : data_o[91];
  assign next_data_o[92] = next_ready_o ? data_reg[92] : data_o[92];
  assign next_data_o[93] = next_ready_o ? data_reg[93] : data_o[93];
  assign next_data_o[94] = next_ready_o ? data_reg[94] : data_o[94];
  assign next_data_o[95] = next_ready_o ? data_reg[95] : data_o[95];
  assign next_data_o[96] = next_ready_o ? data_reg[96] : data_o[96];
  assign next_data_o[97] = next_ready_o ? data_reg[97] : data_o[97];
  assign next_data_o[98] = next_ready_o ? data_reg[98] : data_o[98];
  assign next_data_o[99] = next_ready_o ? data_reg[99] : data_o[99];
  assign _0543_ = decrypt_i ? outy[9] : outx[9];
  assign next_data_o[9] = next_ready_o ? _0543_ : data_o[9];
  assign _0544_ = ~state[0];
  assign _0545_ = state[1] & _0544_;
  assign _0546_ = _0545_ & data_i[32];
  assign _0547_ = ~state[1];
  assign _0548_ = _0547_ & _0544_;
  assign _0549_ = data_i[96] & start_i;
  assign _0550_ = _0549_ & _0548_;
  assign _0551_ = _0547_ & state[0];
  assign _0552_ = _0551_ & data_i[64];
  assign _0553_ = _0552_ | _0550_;
  assign _0554_ = _0553_ | _0546_;
  assign mix_word[0] = next_ready_o ? data_i[0] : _0554_;
  assign _0555_ = _0545_ & data_i[42];
  assign _0556_ = data_i[106] & start_i;
  assign _0557_ = _0556_ & _0548_;
  assign _0558_ = _0551_ & data_i[74];
  assign _0559_ = _0558_ | _0557_;
  assign _0560_ = _0559_ | _0555_;
  assign mix_word[10] = next_ready_o ? data_i[10] : _0560_;
  assign _0561_ = _0545_ & data_i[43];
  assign _0562_ = data_i[107] & start_i;
  assign _0563_ = _0562_ & _0548_;
  assign _0564_ = _0551_ & data_i[75];
  assign _0565_ = _0564_ | _0563_;
  assign _0566_ = _0565_ | _0561_;
  assign mix_word[11] = next_ready_o ? data_i[11] : _0566_;
  assign _0567_ = _0545_ & data_i[44];
  assign _0568_ = data_i[108] & start_i;
  assign _0569_ = _0568_ & _0548_;
  assign _0570_ = _0551_ & data_i[76];
  assign _0571_ = _0570_ | _0569_;
  assign _0572_ = _0571_ | _0567_;
  assign mix_word[12] = next_ready_o ? data_i[12] : _0572_;
  assign _0573_ = _0545_ & data_i[45];
  assign _0574_ = data_i[109] & start_i;
  assign _0575_ = _0574_ & _0548_;
  assign _0576_ = _0551_ & data_i[77];
  assign _0577_ = _0576_ | _0575_;
  assign _0578_ = _0577_ | _0573_;
  assign mix_word[13] = next_ready_o ? data_i[13] : _0578_;
  assign _0579_ = _0545_ & data_i[46];
  assign _0580_ = data_i[110] & start_i;
  assign _0581_ = _0580_ & _0548_;
  assign _0582_ = _0551_ & data_i[78];
  assign _0583_ = _0582_ | _0581_;
  assign _0584_ = _0583_ | _0579_;
  assign mix_word[14] = next_ready_o ? data_i[14] : _0584_;
  assign _0585_ = _0545_ & data_i[47];
  assign _0586_ = data_i[111] & start_i;
  assign _0587_ = _0586_ & _0548_;
  assign _0588_ = _0551_ & data_i[79];
  assign _0589_ = _0588_ | _0587_;
  assign _0590_ = _0589_ | _0585_;
  assign mix_word[15] = next_ready_o ? data_i[15] : _0590_;
  assign _0591_ = _0545_ & data_i[48];
  assign _0592_ = data_i[112] & start_i;
  assign _0593_ = _0592_ & _0548_;
  assign _0594_ = _0551_ & data_i[80];
  assign _0595_ = _0594_ | _0593_;
  assign _0596_ = _0595_ | _0591_;
  assign mix_word[16] = next_ready_o ? data_i[16] : _0596_;
  assign _0597_ = _0545_ & data_i[49];
  assign _0598_ = data_i[113] & start_i;
  assign _0599_ = _0598_ & _0548_;
  assign _0600_ = _0551_ & data_i[81];
  assign _0601_ = _0600_ | _0599_;
  assign _0602_ = _0601_ | _0597_;
  assign mix_word[17] = next_ready_o ? data_i[17] : _0602_;
  assign _0603_ = _0545_ & data_i[50];
  assign _0604_ = data_i[114] & start_i;
  assign _0605_ = _0604_ & _0548_;
  assign _0606_ = _0551_ & data_i[82];
  assign _0607_ = _0606_ | _0605_;
  assign _0608_ = _0607_ | _0603_;
  assign mix_word[18] = next_ready_o ? data_i[18] : _0608_;
  assign _0609_ = _0545_ & data_i[51];
  assign _0610_ = data_i[115] & start_i;
  assign _0611_ = _0610_ & _0548_;
  assign _0612_ = _0551_ & data_i[83];
  assign _0613_ = _0612_ | _0611_;
  assign _0614_ = _0613_ | _0609_;
  assign mix_word[19] = next_ready_o ? data_i[19] : _0614_;
  assign _0615_ = _0545_ & data_i[33];
  assign _0616_ = data_i[97] & start_i;
  assign _0617_ = _0616_ & _0548_;
  assign _0618_ = _0551_ & data_i[65];
  assign _0619_ = _0618_ | _0617_;
  assign _0620_ = _0619_ | _0615_;
  assign mix_word[1] = next_ready_o ? data_i[1] : _0620_;
  assign _0621_ = _0545_ & data_i[52];
  assign _0622_ = data_i[116] & start_i;
  assign _0623_ = _0622_ & _0548_;
  assign _0624_ = _0551_ & data_i[84];
  assign _0625_ = _0624_ | _0623_;
  assign _0626_ = _0625_ | _0621_;
  assign mix_word[20] = next_ready_o ? data_i[20] : _0626_;
  assign _0627_ = _0545_ & data_i[53];
  assign _0628_ = data_i[117] & start_i;
  assign _0629_ = _0628_ & _0548_;
  assign _0630_ = _0551_ & data_i[85];
  assign _0631_ = _0630_ | _0629_;
  assign _0632_ = _0631_ | _0627_;
  assign mix_word[21] = next_ready_o ? data_i[21] : _0632_;
  assign _0633_ = _0545_ & data_i[54];
  assign _0634_ = data_i[118] & start_i;
  assign _0635_ = _0634_ & _0548_;
  assign _0636_ = _0551_ & data_i[86];
  assign _0637_ = _0636_ | _0635_;
  assign _0638_ = _0637_ | _0633_;
  assign mix_word[22] = next_ready_o ? data_i[22] : _0638_;
  assign _0639_ = _0545_ & data_i[55];
  assign _0640_ = data_i[119] & start_i;
  assign _0641_ = _0640_ & _0548_;
  assign _0642_ = _0551_ & data_i[87];
  assign _0643_ = _0642_ | _0641_;
  assign _0644_ = _0643_ | _0639_;
  assign mix_word[23] = next_ready_o ? data_i[23] : _0644_;
  assign _0645_ = _0545_ & data_i[56];
  assign _0646_ = data_i[120] & start_i;
  assign _0647_ = _0646_ & _0548_;
  assign _0648_ = _0551_ & data_i[88];
  assign _0649_ = _0648_ | _0647_;
  assign _0650_ = _0649_ | _0645_;
  assign mix_word[24] = next_ready_o ? data_i[24] : _0650_;
  assign _0651_ = _0545_ & data_i[57];
  assign _0652_ = data_i[121] & start_i;
  assign _0653_ = _0652_ & _0548_;
  assign _0654_ = _0551_ & data_i[89];
  assign _0655_ = _0654_ | _0653_;
  assign _0656_ = _0655_ | _0651_;
  assign mix_word[25] = next_ready_o ? data_i[25] : _0656_;
  assign _0657_ = _0545_ & data_i[58];
  assign _0658_ = data_i[122] & start_i;
  assign _0659_ = _0658_ & _0548_;
  assign _0660_ = _0551_ & data_i[90];
  assign _0661_ = _0660_ | _0659_;
  assign _0662_ = _0661_ | _0657_;
  assign mix_word[26] = next_ready_o ? data_i[26] : _0662_;
  assign _0663_ = _0545_ & data_i[59];
  assign _0664_ = data_i[123] & start_i;
  assign _0665_ = _0664_ & _0548_;
  assign _0666_ = _0551_ & data_i[91];
  assign _0667_ = _0666_ | _0665_;
  assign _0668_ = _0667_ | _0663_;
  assign mix_word[27] = next_ready_o ? data_i[27] : _0668_;
  assign _0669_ = _0545_ & data_i[60];
  assign _0670_ = data_i[124] & start_i;
  assign _0671_ = _0670_ & _0548_;
  assign _0672_ = _0551_ & data_i[92];
  assign _0673_ = _0672_ | _0671_;
  assign _0674_ = _0673_ | _0669_;
  assign mix_word[28] = next_ready_o ? data_i[28] : _0674_;
  assign _0675_ = _0545_ & data_i[61];
  assign _0676_ = data_i[125] & start_i;
  assign _0677_ = _0676_ & _0548_;
  assign _0678_ = _0551_ & data_i[93];
  assign _0679_ = _0678_ | _0677_;
  assign _0680_ = _0679_ | _0675_;
  assign mix_word[29] = next_ready_o ? data_i[29] : _0680_;
  assign _0681_ = _0545_ & data_i[34];
  assign _0000_ = data_i[98] & start_i;
  assign _0001_ = _0000_ & _0548_;
  assign _0002_ = _0551_ & data_i[66];
  assign _0003_ = _0002_ | _0001_;
  assign _0004_ = _0003_ | _0681_;
  assign mix_word[2] = next_ready_o ? data_i[2] : _0004_;
  assign _0005_ = _0545_ & data_i[62];
  assign _0006_ = data_i[126] & start_i;
  assign _0007_ = _0006_ & _0548_;
  assign _0008_ = _0551_ & data_i[94];
  assign _0009_ = _0008_ | _0007_;
  assign _0010_ = _0009_ | _0005_;
  assign mix_word[30] = next_ready_o ? data_i[30] : _0010_;
  assign _0011_ = _0545_ & data_i[63];
  assign _0012_ = data_i[127] & start_i;
  assign _0013_ = _0012_ & _0548_;
  assign _0014_ = _0551_ & data_i[95];
  assign _0015_ = _0014_ | _0013_;
  assign _0016_ = _0015_ | _0011_;
  assign mix_word[31] = next_ready_o ? data_i[31] : _0016_;
  assign _0017_ = _0545_ & data_i[35];
  assign _0018_ = data_i[99] & start_i;
  assign _0019_ = _0018_ & _0548_;
  assign _0020_ = _0551_ & data_i[67];
  assign _0021_ = _0020_ | _0019_;
  assign _0022_ = _0021_ | _0017_;
  assign mix_word[3] = next_ready_o ? data_i[3] : _0022_;
  assign _0023_ = _0545_ & data_i[36];
  assign _0024_ = data_i[100] & start_i;
  assign _0025_ = _0024_ & _0548_;
  assign _0026_ = _0551_ & data_i[68];
  assign _0027_ = _0026_ | _0025_;
  assign _0028_ = _0027_ | _0023_;
  assign mix_word[4] = next_ready_o ? data_i[4] : _0028_;
  assign _0029_ = _0545_ & data_i[37];
  assign _0030_ = data_i[101] & start_i;
  assign _0031_ = _0030_ & _0548_;
  assign _0032_ = _0551_ & data_i[69];
  assign _0033_ = _0032_ | _0031_;
  assign _0034_ = _0033_ | _0029_;
  assign mix_word[5] = next_ready_o ? data_i[5] : _0034_;
  assign _0035_ = _0545_ & data_i[38];
  assign _0036_ = data_i[102] & start_i;
  assign _0037_ = _0036_ & _0548_;
  assign _0038_ = _0551_ & data_i[70];
  assign _0039_ = _0038_ | _0037_;
  assign _0040_ = _0039_ | _0035_;
  assign mix_word[6] = next_ready_o ? data_i[6] : _0040_;
  assign _0041_ = _0545_ & data_i[39];
  assign _0042_ = data_i[103] & start_i;
  assign _0043_ = _0042_ & _0548_;
  assign _0044_ = _0551_ & data_i[71];
  assign _0045_ = _0044_ | _0043_;
  assign _0046_ = _0045_ | _0041_;
  assign mix_word[7] = next_ready_o ? data_i[7] : _0046_;
  assign _0047_ = _0545_ & data_i[40];
  assign _0048_ = data_i[104] & start_i;
  assign _0049_ = _0048_ & _0548_;
  assign _0050_ = _0551_ & data_i[72];
  assign _0051_ = _0050_ | _0049_;
  assign _0052_ = _0051_ | _0047_;
  assign mix_word[8] = next_ready_o ? data_i[8] : _0052_;
  assign _0053_ = _0545_ & data_i[41];
  assign _0054_ = data_i[105] & start_i;
  assign _0055_ = _0054_ & _0548_;
  assign _0056_ = _0551_ & data_i[73];
  assign _0057_ = _0056_ | _0055_;
  assign _0058_ = _0057_ | _0053_;
  assign mix_word[9] = next_ready_o ? data_i[9] : _0058_;
  assign _0059_ = ~start_i;
  assign _0060_ = _0059_ ? data_reg[100] : _0538_;
  assign _0061_ = _0060_ & _0548_;
  assign _0062_ = _0551_ & data_reg[100];
  assign _0063_ = _0545_ & data_reg[100];
  assign _0064_ = _0063_ | _0062_;
  assign _0065_ = _0064_ | _0061_;
  assign next_data_reg[100] = next_ready_o ? data_reg[100] : _0065_;
  assign _0066_ = _0059_ ? data_reg[101] : _0539_;
  assign _0067_ = _0066_ & _0548_;
  assign _0068_ = _0551_ & data_reg[101];
  assign _0069_ = _0545_ & data_reg[101];
  assign _0070_ = _0069_ | _0068_;
  assign _0071_ = _0070_ | _0067_;
  assign next_data_reg[101] = next_ready_o ? data_reg[101] : _0071_;
  assign _0072_ = _0059_ ? data_reg[102] : _0540_;
  assign _0073_ = _0072_ & _0548_;
  assign _0074_ = _0551_ & data_reg[102];
  assign _0075_ = _0545_ & data_reg[102];
  assign _0076_ = _0075_ | _0074_;
  assign _0077_ = _0076_ | _0073_;
  assign next_data_reg[102] = next_ready_o ? data_reg[102] : _0077_;
  assign _0078_ = _0059_ ? data_reg[103] : _0541_;
  assign _0079_ = _0078_ & _0548_;
  assign _0080_ = _0551_ & data_reg[103];
  assign _0081_ = _0545_ & data_reg[103];
  assign _0082_ = _0081_ | _0080_;
  assign _0083_ = _0082_ | _0079_;
  assign next_data_reg[103] = next_ready_o ? data_reg[103] : _0083_;
  assign _0084_ = _0059_ ? data_reg[104] : _0542_;
  assign _0085_ = _0084_ & _0548_;
  assign _0086_ = _0551_ & data_reg[104];
  assign _0087_ = _0545_ & data_reg[104];
  assign _0088_ = _0087_ | _0086_;
  assign _0089_ = _0088_ | _0085_;
  assign next_data_reg[104] = next_ready_o ? data_reg[104] : _0089_;
  assign _0090_ = _0059_ ? data_reg[105] : _0543_;
  assign _0091_ = _0090_ & _0548_;
  assign _0092_ = _0551_ & data_reg[105];
  assign _0093_ = _0545_ & data_reg[105];
  assign _0094_ = _0093_ | _0092_;
  assign _0095_ = _0094_ | _0091_;
  assign next_data_reg[105] = next_ready_o ? data_reg[105] : _0095_;
  assign _0096_ = _0059_ ? data_reg[106] : _0513_;
  assign _0097_ = _0096_ & _0548_;
  assign _0098_ = _0551_ & data_reg[106];
  assign _0099_ = _0545_ & data_reg[106];
  assign _0100_ = _0099_ | _0098_;
  assign _0101_ = _0100_ | _0097_;
  assign next_data_reg[106] = next_ready_o ? data_reg[106] : _0101_;
  assign _0102_ = _0059_ ? data_reg[107] : _0514_;
  assign _0103_ = _0102_ & _0548_;
  assign _0104_ = _0551_ & data_reg[107];
  assign _0105_ = _0545_ & data_reg[107];
  assign _0106_ = _0105_ | _0104_;
  assign _0107_ = _0106_ | _0103_;
  assign next_data_reg[107] = next_ready_o ? data_reg[107] : _0107_;
  assign _0108_ = _0059_ ? data_reg[108] : _0515_;
  assign _0109_ = _0108_ & _0548_;
  assign _0110_ = _0551_ & data_reg[108];
  assign _0111_ = _0545_ & data_reg[108];
  assign _0112_ = _0111_ | _0110_;
  assign _0113_ = _0112_ | _0109_;
  assign next_data_reg[108] = next_ready_o ? data_reg[108] : _0113_;
  assign _0114_ = _0059_ ? data_reg[109] : _0516_;
  assign _0115_ = _0114_ & _0548_;
  assign _0116_ = _0551_ & data_reg[109];
  assign _0117_ = _0545_ & data_reg[109];
  assign _0118_ = _0117_ | _0116_;
  assign _0119_ = _0118_ | _0115_;
  assign next_data_reg[109] = next_ready_o ? data_reg[109] : _0119_;
  assign _0120_ = _0059_ ? data_reg[110] : _0517_;
  assign _0121_ = _0120_ & _0548_;
  assign _0122_ = _0551_ & data_reg[110];
  assign _0123_ = _0545_ & data_reg[110];
  assign _0124_ = _0123_ | _0122_;
  assign _0125_ = _0124_ | _0121_;
  assign next_data_reg[110] = next_ready_o ? data_reg[110] : _0125_;
  assign _0126_ = _0059_ ? data_reg[111] : _0518_;
  assign _0127_ = _0126_ & _0548_;
  assign _0128_ = _0551_ & data_reg[111];
  assign _0129_ = _0545_ & data_reg[111];
  assign _0130_ = _0129_ | _0128_;
  assign _0131_ = _0130_ | _0127_;
  assign next_data_reg[111] = next_ready_o ? data_reg[111] : _0131_;
  assign _0132_ = _0059_ ? data_reg[112] : _0519_;
  assign _0133_ = _0132_ & _0548_;
  assign _0134_ = _0551_ & data_reg[112];
  assign _0135_ = _0545_ & data_reg[112];
  assign _0136_ = _0135_ | _0134_;
  assign _0137_ = _0136_ | _0133_;
  assign next_data_reg[112] = next_ready_o ? data_reg[112] : _0137_;
  assign _0138_ = _0059_ ? data_reg[113] : _0520_;
  assign _0139_ = _0138_ & _0548_;
  assign _0140_ = _0551_ & data_reg[113];
  assign _0141_ = _0545_ & data_reg[113];
  assign _0142_ = _0141_ | _0140_;
  assign _0143_ = _0142_ | _0139_;
  assign next_data_reg[113] = next_ready_o ? data_reg[113] : _0143_;
  assign _0144_ = _0059_ ? data_reg[114] : _0521_;
  assign _0145_ = _0144_ & _0548_;
  assign _0146_ = _0551_ & data_reg[114];
  assign _0147_ = _0545_ & data_reg[114];
  assign _0148_ = _0147_ | _0146_;
  assign _0149_ = _0148_ | _0145_;
  assign next_data_reg[114] = next_ready_o ? data_reg[114] : _0149_;
  assign _0150_ = _0059_ ? data_reg[115] : _0522_;
  assign _0151_ = _0150_ & _0548_;
  assign _0152_ = _0551_ & data_reg[115];
  assign _0153_ = _0545_ & data_reg[115];
  assign _0154_ = _0153_ | _0152_;
  assign _0155_ = _0154_ | _0151_;
  assign next_data_reg[115] = next_ready_o ? data_reg[115] : _0155_;
  assign _0156_ = _0059_ ? data_reg[116] : _0524_;
  assign _0157_ = _0156_ & _0548_;
  assign _0158_ = _0551_ & data_reg[116];
  assign _0159_ = _0545_ & data_reg[116];
  assign _0160_ = _0159_ | _0158_;
  assign _0161_ = _0160_ | _0157_;
  assign next_data_reg[116] = next_ready_o ? data_reg[116] : _0161_;
  assign _0162_ = _0059_ ? data_reg[117] : _0525_;
  assign _0163_ = _0162_ & _0548_;
  assign _0164_ = _0551_ & data_reg[117];
  assign _0165_ = _0545_ & data_reg[117];
  assign _0166_ = _0165_ | _0164_;
  assign _0167_ = _0166_ | _0163_;
  assign next_data_reg[117] = next_ready_o ? data_reg[117] : _0167_;
  assign _0168_ = _0059_ ? data_reg[118] : _0526_;
  assign _0169_ = _0168_ & _0548_;
  assign _0170_ = _0551_ & data_reg[118];
  assign _0171_ = _0545_ & data_reg[118];
  assign _0172_ = _0171_ | _0170_;
  assign _0173_ = _0172_ | _0169_;
  assign next_data_reg[118] = next_ready_o ? data_reg[118] : _0173_;
  assign _0174_ = _0059_ ? data_reg[119] : _0527_;
  assign _0175_ = _0174_ & _0548_;
  assign _0176_ = _0551_ & data_reg[119];
  assign _0177_ = _0545_ & data_reg[119];
  assign _0178_ = _0177_ | _0176_;
  assign _0179_ = _0178_ | _0175_;
  assign next_data_reg[119] = next_ready_o ? data_reg[119] : _0179_;
  assign _0180_ = _0059_ ? data_reg[120] : _0528_;
  assign _0181_ = _0180_ & _0548_;
  assign _0182_ = _0551_ & data_reg[120];
  assign _0183_ = _0545_ & data_reg[120];
  assign _0184_ = _0183_ | _0182_;
  assign _0185_ = _0184_ | _0181_;
  assign next_data_reg[120] = next_ready_o ? data_reg[120] : _0185_;
  assign _0186_ = _0059_ ? data_reg[121] : _0529_;
  assign _0187_ = _0186_ & _0548_;
  assign _0188_ = _0551_ & data_reg[121];
  assign _0189_ = _0545_ & data_reg[121];
  assign _0190_ = _0189_ | _0188_;
  assign _0191_ = _0190_ | _0187_;
  assign next_data_reg[121] = next_ready_o ? data_reg[121] : _0191_;
  assign _0192_ = _0059_ ? data_reg[122] : _0530_;
  assign _0193_ = _0192_ & _0548_;
  assign _0194_ = _0551_ & data_reg[122];
  assign _0195_ = _0545_ & data_reg[122];
  assign _0196_ = _0195_ | _0194_;
  assign _0197_ = _0196_ | _0193_;
  assign next_data_reg[122] = next_ready_o ? data_reg[122] : _0197_;
  assign _0198_ = _0059_ ? data_reg[123] : _0531_;
  assign _0199_ = _0198_ & _0548_;
  assign _0200_ = _0551_ & data_reg[123];
  assign _0201_ = _0545_ & data_reg[123];
  assign _0202_ = _0201_ | _0200_;
  assign _0203_ = _0202_ | _0199_;
  assign next_data_reg[123] = next_ready_o ? data_reg[123] : _0203_;
  assign _0204_ = _0059_ ? data_reg[124] : _0532_;
  assign _0205_ = _0204_ & _0548_;
  assign _0206_ = _0551_ & data_reg[124];
  assign _0207_ = _0545_ & data_reg[124];
  assign _0208_ = _0207_ | _0206_;
  assign _0209_ = _0208_ | _0205_;
  assign next_data_reg[124] = next_ready_o ? data_reg[124] : _0209_;
  assign _0210_ = _0059_ ? data_reg[125] : _0533_;
  assign _0211_ = _0210_ & _0548_;
  assign _0212_ = _0551_ & data_reg[125];
  assign _0213_ = _0545_ & data_reg[125];
  assign _0214_ = _0213_ | _0212_;
  assign _0215_ = _0214_ | _0211_;
  assign next_data_reg[125] = next_ready_o ? data_reg[125] : _0215_;
  assign _0216_ = _0059_ ? data_reg[126] : _0535_;
  assign _0217_ = _0216_ & _0548_;
  assign _0218_ = _0551_ & data_reg[126];
  assign _0219_ = _0545_ & data_reg[126];
  assign _0220_ = _0219_ | _0218_;
  assign _0221_ = _0220_ | _0217_;
  assign next_data_reg[126] = next_ready_o ? data_reg[126] : _0221_;
  assign _0222_ = _0059_ ? data_reg[127] : _0536_;
  assign _0223_ = _0222_ & _0548_;
  assign _0224_ = _0551_ & data_reg[127];
  assign _0225_ = _0545_ & data_reg[127];
  assign _0226_ = _0225_ | _0224_;
  assign _0227_ = _0226_ | _0223_;
  assign next_data_reg[127] = next_ready_o ? data_reg[127] : _0227_;
  assign _0228_ = _0512_ & _0545_;
  assign _0229_ = _0548_ & data_reg[32];
  assign _0230_ = _0551_ & data_reg[32];
  assign _0231_ = _0230_ | _0229_;
  assign _0232_ = _0231_ | _0228_;
  assign next_data_reg[32] = next_ready_o ? data_reg[32] : _0232_;
  assign _0233_ = _0523_ & _0545_;
  assign _0234_ = _0548_ & data_reg[33];
  assign _0235_ = _0551_ & data_reg[33];
  assign _0236_ = _0235_ | _0234_;
  assign _0237_ = _0236_ | _0233_;
  assign next_data_reg[33] = next_ready_o ? data_reg[33] : _0237_;
  assign _0238_ = _0534_ & _0545_;
  assign _0239_ = _0548_ & data_reg[34];
  assign _0240_ = _0551_ & data_reg[34];
  assign _0241_ = _0240_ | _0239_;
  assign _0242_ = _0241_ | _0238_;
  assign next_data_reg[34] = next_ready_o ? data_reg[34] : _0242_;
  assign _0243_ = _0537_ & _0545_;
  assign _0244_ = _0548_ & data_reg[35];
  assign _0245_ = _0551_ & data_reg[35];
  assign _0246_ = _0245_ | _0244_;
  assign _0247_ = _0246_ | _0243_;
  assign next_data_reg[35] = next_ready_o ? data_reg[35] : _0247_;
  assign _0248_ = _0538_ & _0545_;
  assign _0249_ = _0548_ & data_reg[36];
  assign _0250_ = _0551_ & data_reg[36];
  assign _0251_ = _0250_ | _0249_;
  assign _0252_ = _0251_ | _0248_;
  assign next_data_reg[36] = next_ready_o ? data_reg[36] : _0252_;
  assign _0253_ = _0539_ & _0545_;
  assign _0254_ = _0548_ & data_reg[37];
  assign _0255_ = _0551_ & data_reg[37];
  assign _0256_ = _0255_ | _0254_;
  assign _0257_ = _0256_ | _0253_;
  assign next_data_reg[37] = next_ready_o ? data_reg[37] : _0257_;
  assign _0258_ = _0540_ & _0545_;
  assign _0259_ = _0548_ & data_reg[38];
  assign _0260_ = _0551_ & data_reg[38];
  assign _0261_ = _0260_ | _0259_;
  assign _0262_ = _0261_ | _0258_;
  assign next_data_reg[38] = next_ready_o ? data_reg[38] : _0262_;
  assign _0263_ = _0541_ & _0545_;
  assign _0264_ = _0548_ & data_reg[39];
  assign _0265_ = _0551_ & data_reg[39];
  assign _0266_ = _0265_ | _0264_;
  assign _0267_ = _0266_ | _0263_;
  assign next_data_reg[39] = next_ready_o ? data_reg[39] : _0267_;
  assign _0268_ = _0542_ & _0545_;
  assign _0269_ = _0548_ & data_reg[40];
  assign _0270_ = _0551_ & data_reg[40];
  assign _0271_ = _0270_ | _0269_;
  assign _0272_ = _0271_ | _0268_;
  assign next_data_reg[40] = next_ready_o ? data_reg[40] : _0272_;
  assign _0273_ = _0543_ & _0545_;
  assign _0274_ = _0548_ & data_reg[41];
  assign _0275_ = _0551_ & data_reg[41];
  assign _0276_ = _0275_ | _0274_;
  assign _0277_ = _0276_ | _0273_;
  assign next_data_reg[41] = next_ready_o ? data_reg[41] : _0277_;
  assign _0278_ = _0513_ & _0545_;
  assign _0279_ = _0548_ & data_reg[42];
  assign _0280_ = _0551_ & data_reg[42];
  assign _0281_ = _0280_ | _0279_;
  assign _0282_ = _0281_ | _0278_;
  assign next_data_reg[42] = next_ready_o ? data_reg[42] : _0282_;
  assign _0283_ = _0514_ & _0545_;
  assign _0284_ = _0548_ & data_reg[43];
  assign _0285_ = _0551_ & data_reg[43];
  assign _0286_ = _0285_ | _0284_;
  assign _0287_ = _0286_ | _0283_;
  assign next_data_reg[43] = next_ready_o ? data_reg[43] : _0287_;
  assign _0288_ = _0515_ & _0545_;
  assign _0289_ = _0548_ & data_reg[44];
  assign _0290_ = _0551_ & data_reg[44];
  assign _0291_ = _0290_ | _0289_;
  assign _0292_ = _0291_ | _0288_;
  assign next_data_reg[44] = next_ready_o ? data_reg[44] : _0292_;
  assign _0293_ = _0516_ & _0545_;
  assign _0294_ = _0548_ & data_reg[45];
  assign _0295_ = _0551_ & data_reg[45];
  assign _0296_ = _0295_ | _0294_;
  assign _0297_ = _0296_ | _0293_;
  assign next_data_reg[45] = next_ready_o ? data_reg[45] : _0297_;
  assign _0298_ = _0517_ & _0545_;
  assign _0299_ = _0548_ & data_reg[46];
  assign _0300_ = _0551_ & data_reg[46];
  assign _0301_ = _0300_ | _0299_;
  assign _0302_ = _0301_ | _0298_;
  assign next_data_reg[46] = next_ready_o ? data_reg[46] : _0302_;
  assign _0303_ = _0518_ & _0545_;
  assign _0304_ = _0548_ & data_reg[47];
  assign _0305_ = _0551_ & data_reg[47];
  assign _0306_ = _0305_ | _0304_;
  assign _0307_ = _0306_ | _0303_;
  assign next_data_reg[47] = next_ready_o ? data_reg[47] : _0307_;
  assign _0308_ = _0519_ & _0545_;
  assign _0309_ = _0548_ & data_reg[48];
  assign _0310_ = _0551_ & data_reg[48];
  assign _0311_ = _0310_ | _0309_;
  assign _0312_ = _0311_ | _0308_;
  assign next_data_reg[48] = next_ready_o ? data_reg[48] : _0312_;
  assign _0313_ = _0520_ & _0545_;
  assign _0314_ = _0548_ & data_reg[49];
  assign _0315_ = _0551_ & data_reg[49];
  assign _0316_ = _0315_ | _0314_;
  assign _0317_ = _0316_ | _0313_;
  assign next_data_reg[49] = next_ready_o ? data_reg[49] : _0317_;
  assign _0318_ = _0521_ & _0545_;
  assign _0319_ = _0548_ & data_reg[50];
  assign _0320_ = _0551_ & data_reg[50];
  assign _0321_ = _0320_ | _0319_;
  assign _0322_ = _0321_ | _0318_;
  assign next_data_reg[50] = next_ready_o ? data_reg[50] : _0322_;
  assign _0323_ = _0522_ & _0545_;
  assign _0324_ = _0548_ & data_reg[51];
  assign _0325_ = _0551_ & data_reg[51];
  assign _0326_ = _0325_ | _0324_;
  assign _0327_ = _0326_ | _0323_;
  assign next_data_reg[51] = next_ready_o ? data_reg[51] : _0327_;
  assign _0328_ = _0524_ & _0545_;
  assign _0329_ = _0548_ & data_reg[52];
  assign _0330_ = _0551_ & data_reg[52];
  assign _0331_ = _0330_ | _0329_;
  assign _0332_ = _0331_ | _0328_;
  assign next_data_reg[52] = next_ready_o ? data_reg[52] : _0332_;
  assign _0333_ = _0525_ & _0545_;
  assign _0334_ = _0548_ & data_reg[53];
  assign _0335_ = _0551_ & data_reg[53];
  assign _0336_ = _0335_ | _0334_;
  assign _0337_ = _0336_ | _0333_;
  assign next_data_reg[53] = next_ready_o ? data_reg[53] : _0337_;
  assign _0338_ = _0526_ & _0545_;
  assign _0339_ = _0548_ & data_reg[54];
  assign _0340_ = _0551_ & data_reg[54];
  assign _0341_ = _0340_ | _0339_;
  assign _0342_ = _0341_ | _0338_;
  assign next_data_reg[54] = next_ready_o ? data_reg[54] : _0342_;
  assign _0343_ = _0527_ & _0545_;
  assign _0344_ = _0548_ & data_reg[55];
  assign _0345_ = _0551_ & data_reg[55];
  assign _0346_ = _0345_ | _0344_;
  assign _0347_ = _0346_ | _0343_;
  assign next_data_reg[55] = next_ready_o ? data_reg[55] : _0347_;
  assign _0348_ = _0528_ & _0545_;
  assign _0349_ = _0548_ & data_reg[56];
  assign _0350_ = _0551_ & data_reg[56];
  assign _0351_ = _0350_ | _0349_;
  assign _0352_ = _0351_ | _0348_;
  assign next_data_reg[56] = next_ready_o ? data_reg[56] : _0352_;
  assign _0353_ = _0529_ & _0545_;
  assign _0354_ = _0548_ & data_reg[57];
  assign _0355_ = _0551_ & data_reg[57];
  assign _0356_ = _0355_ | _0354_;
  assign _0357_ = _0356_ | _0353_;
  assign next_data_reg[57] = next_ready_o ? data_reg[57] : _0357_;
  assign _0358_ = _0530_ & _0545_;
  assign _0359_ = _0548_ & data_reg[58];
  assign _0360_ = _0551_ & data_reg[58];
  assign _0361_ = _0360_ | _0359_;
  assign _0362_ = _0361_ | _0358_;
  assign next_data_reg[58] = next_ready_o ? data_reg[58] : _0362_;
  assign _0363_ = _0531_ & _0545_;
  assign _0364_ = _0548_ & data_reg[59];
  assign _0365_ = _0551_ & data_reg[59];
  assign _0366_ = _0365_ | _0364_;
  assign _0367_ = _0366_ | _0363_;
  assign next_data_reg[59] = next_ready_o ? data_reg[59] : _0367_;
  assign _0368_ = _0532_ & _0545_;
  assign _0369_ = _0548_ & data_reg[60];
  assign _0370_ = _0551_ & data_reg[60];
  assign _0371_ = _0370_ | _0369_;
  assign _0372_ = _0371_ | _0368_;
  assign next_data_reg[60] = next_ready_o ? data_reg[60] : _0372_;
  assign _0373_ = _0533_ & _0545_;
  assign _0374_ = _0548_ & data_reg[61];
  assign _0375_ = _0551_ & data_reg[61];
  assign _0376_ = _0375_ | _0374_;
  assign _0377_ = _0376_ | _0373_;
  assign next_data_reg[61] = next_ready_o ? data_reg[61] : _0377_;
  assign _0378_ = _0535_ & _0545_;
  assign _0379_ = _0548_ & data_reg[62];
  assign _0380_ = _0551_ & data_reg[62];
  assign _0381_ = _0380_ | _0379_;
  assign _0382_ = _0381_ | _0378_;
  assign next_data_reg[62] = next_ready_o ? data_reg[62] : _0382_;
  assign _0383_ = _0536_ & _0545_;
  assign _0384_ = _0548_ & data_reg[63];
  assign _0385_ = _0551_ & data_reg[63];
  assign _0386_ = _0385_ | _0384_;
  assign _0387_ = _0386_ | _0383_;
  assign next_data_reg[63] = next_ready_o ? data_reg[63] : _0387_;
  assign _0388_ = _0512_ & _0551_;
  assign _0389_ = _0544_ & data_reg[64];
  assign _0390_ = _0389_ | _0388_;
  assign next_data_reg[64] = next_ready_o ? data_reg[64] : _0390_;
  assign _0391_ = _0523_ & _0551_;
  assign _0392_ = _0544_ & data_reg[65];
  assign _0393_ = _0392_ | _0391_;
  assign next_data_reg[65] = next_ready_o ? data_reg[65] : _0393_;
  assign _0394_ = _0534_ & _0551_;
  assign _0395_ = _0544_ & data_reg[66];
  assign _0396_ = _0395_ | _0394_;
  assign next_data_reg[66] = next_ready_o ? data_reg[66] : _0396_;
  assign _0397_ = _0537_ & _0551_;
  assign _0398_ = _0544_ & data_reg[67];
  assign _0399_ = _0398_ | _0397_;
  assign next_data_reg[67] = next_ready_o ? data_reg[67] : _0399_;
  assign _0400_ = _0538_ & _0551_;
  assign _0401_ = _0544_ & data_reg[68];
  assign _0402_ = _0401_ | _0400_;
  assign next_data_reg[68] = next_ready_o ? data_reg[68] : _0402_;
  assign _0403_ = _0539_ & _0551_;
  assign _0404_ = _0544_ & data_reg[69];
  assign _0405_ = _0404_ | _0403_;
  assign next_data_reg[69] = next_ready_o ? data_reg[69] : _0405_;
  assign _0406_ = _0540_ & _0551_;
  assign _0407_ = _0544_ & data_reg[70];
  assign _0408_ = _0407_ | _0406_;
  assign next_data_reg[70] = next_ready_o ? data_reg[70] : _0408_;
  assign _0409_ = _0541_ & _0551_;
  assign _0410_ = _0544_ & data_reg[71];
  assign _0411_ = _0410_ | _0409_;
  assign next_data_reg[71] = next_ready_o ? data_reg[71] : _0411_;
  assign _0412_ = _0542_ & _0551_;
  assign _0413_ = _0544_ & data_reg[72];
  assign _0414_ = _0413_ | _0412_;
  assign next_data_reg[72] = next_ready_o ? data_reg[72] : _0414_;
  assign _0415_ = _0543_ & _0551_;
  assign _0416_ = _0544_ & data_reg[73];
  assign _0417_ = _0416_ | _0415_;
  assign next_data_reg[73] = next_ready_o ? data_reg[73] : _0417_;
  assign _0418_ = _0513_ & _0551_;
  assign _0419_ = _0544_ & data_reg[74];
  assign _0420_ = _0419_ | _0418_;
  assign next_data_reg[74] = next_ready_o ? data_reg[74] : _0420_;
  assign _0421_ = _0514_ & _0551_;
  assign _0422_ = _0544_ & data_reg[75];
  assign _0423_ = _0422_ | _0421_;
  assign next_data_reg[75] = next_ready_o ? data_reg[75] : _0423_;
  assign _0424_ = _0515_ & _0551_;
  assign _0425_ = _0544_ & data_reg[76];
  assign _0426_ = _0425_ | _0424_;
  assign next_data_reg[76] = next_ready_o ? data_reg[76] : _0426_;
  assign _0427_ = _0516_ & _0551_;
  assign _0428_ = _0544_ & data_reg[77];
  assign _0429_ = _0428_ | _0427_;
  assign next_data_reg[77] = next_ready_o ? data_reg[77] : _0429_;
  assign _0430_ = _0517_ & _0551_;
  assign _0431_ = _0544_ & data_reg[78];
  assign _0432_ = _0431_ | _0430_;
  assign next_data_reg[78] = next_ready_o ? data_reg[78] : _0432_;
  assign _0433_ = _0518_ & _0551_;
  assign _0434_ = _0544_ & data_reg[79];
  assign _0435_ = _0434_ | _0433_;
  assign next_data_reg[79] = next_ready_o ? data_reg[79] : _0435_;
  assign _0436_ = _0519_ & _0551_;
  assign _0437_ = _0544_ & data_reg[80];
  assign _0438_ = _0437_ | _0436_;
  assign next_data_reg[80] = next_ready_o ? data_reg[80] : _0438_;
  assign _0439_ = _0520_ & _0551_;
  assign _0440_ = _0544_ & data_reg[81];
  assign _0441_ = _0440_ | _0439_;
  assign next_data_reg[81] = next_ready_o ? data_reg[81] : _0441_;
  assign _0442_ = _0521_ & _0551_;
  assign _0443_ = _0544_ & data_reg[82];
  assign _0444_ = _0443_ | _0442_;
  assign next_data_reg[82] = next_ready_o ? data_reg[82] : _0444_;
  assign _0445_ = _0522_ & _0551_;
  assign _0446_ = _0544_ & data_reg[83];
  assign _0447_ = _0446_ | _0445_;
  assign next_data_reg[83] = next_ready_o ? data_reg[83] : _0447_;
  assign _0448_ = _0524_ & _0551_;
  assign _0449_ = _0544_ & data_reg[84];
  assign _0450_ = _0449_ | _0448_;
  assign next_data_reg[84] = next_ready_o ? data_reg[84] : _0450_;
  assign _0451_ = _0525_ & _0551_;
  assign _0452_ = _0544_ & data_reg[85];
  assign _0453_ = _0452_ | _0451_;
  assign next_data_reg[85] = next_ready_o ? data_reg[85] : _0453_;
  assign _0454_ = _0526_ & _0551_;
  assign _0455_ = _0544_ & data_reg[86];
  assign _0456_ = _0455_ | _0454_;
  assign next_data_reg[86] = next_ready_o ? data_reg[86] : _0456_;
  assign _0457_ = _0527_ & _0551_;
  assign _0458_ = _0544_ & data_reg[87];
  assign _0459_ = _0458_ | _0457_;
  assign next_data_reg[87] = next_ready_o ? data_reg[87] : _0459_;
  assign _0460_ = _0528_ & _0551_;
  assign _0461_ = _0544_ & data_reg[88];
  assign _0462_ = _0461_ | _0460_;
  assign next_data_reg[88] = next_ready_o ? data_reg[88] : _0462_;
  assign _0463_ = _0529_ & _0551_;
  assign _0464_ = _0544_ & data_reg[89];
  assign _0465_ = _0464_ | _0463_;
  assign next_data_reg[89] = next_ready_o ? data_reg[89] : _0465_;
  assign _0466_ = _0530_ & _0551_;
  assign _0467_ = _0544_ & data_reg[90];
  assign _0468_ = _0467_ | _0466_;
  assign next_data_reg[90] = next_ready_o ? data_reg[90] : _0468_;
  assign _0469_ = _0531_ & _0551_;
  assign _0470_ = _0544_ & data_reg[91];
  assign _0471_ = _0470_ | _0469_;
  assign next_data_reg[91] = next_ready_o ? data_reg[91] : _0471_;
  assign _0472_ = _0532_ & _0551_;
  assign _0473_ = _0544_ & data_reg[92];
  assign _0474_ = _0473_ | _0472_;
  assign next_data_reg[92] = next_ready_o ? data_reg[92] : _0474_;
  assign _0475_ = _0533_ & _0551_;
  assign _0476_ = _0544_ & data_reg[93];
  assign _0477_ = _0476_ | _0475_;
  assign next_data_reg[93] = next_ready_o ? data_reg[93] : _0477_;
  assign _0478_ = _0535_ & _0551_;
  assign _0479_ = _0544_ & data_reg[94];
  assign _0480_ = _0479_ | _0478_;
  assign next_data_reg[94] = next_ready_o ? data_reg[94] : _0480_;
  assign _0481_ = _0536_ & _0551_;
  assign _0482_ = _0544_ & data_reg[95];
  assign _0483_ = _0482_ | _0481_;
  assign next_data_reg[95] = next_ready_o ? data_reg[95] : _0483_;
  assign _0484_ = _0059_ ? data_reg[96] : _0512_;
  assign _0485_ = _0484_ & _0548_;
  assign _0486_ = _0551_ & data_reg[96];
  assign _0487_ = _0545_ & data_reg[96];
  assign _0488_ = _0487_ | _0486_;
  assign _0489_ = _0488_ | _0485_;
  assign next_data_reg[96] = next_ready_o ? data_reg[96] : _0489_;
  assign _0490_ = _0059_ ? data_reg[97] : _0523_;
  assign _0491_ = _0490_ & _0548_;
  assign _0492_ = _0551_ & data_reg[97];
  assign _0493_ = _0545_ & data_reg[97];
  assign _0494_ = _0493_ | _0492_;
  assign _0495_ = _0494_ | _0491_;
  assign next_data_reg[97] = next_ready_o ? data_reg[97] : _0495_;
  assign _0496_ = _0059_ ? data_reg[98] : _0534_;
  assign _0497_ = _0496_ & _0548_;
  assign _0498_ = _0551_ & data_reg[98];
  assign _0499_ = _0545_ & data_reg[98];
  assign _0500_ = _0499_ | _0498_;
  assign _0501_ = _0500_ | _0497_;
  assign next_data_reg[98] = next_ready_o ? data_reg[98] : _0501_;
  assign _0502_ = _0059_ ? data_reg[99] : _0537_;
  assign _0503_ = _0502_ & _0548_;
  assign _0504_ = _0551_ & data_reg[99];
  assign _0505_ = _0545_ & data_reg[99];
  assign _0506_ = _0505_ | _0504_;
  assign _0507_ = _0506_ | _0503_;
  assign next_data_reg[99] = next_ready_o ? data_reg[99] : _0507_;
  assign _0508_ = state[0] | start_i;
  assign _0509_ = _0508_ & _0548_;
  assign next_state[0] = state[1] ? _0544_ : _0509_;
  assign _0510_ = ~next_ready_o;
  assign _0511_ = state[1] ^ state[0];
  assign next_state[1] = _0511_ & _0510_;
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[0] <= 0;
    else
      data_o[0] <= next_data_o[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[100] <= 0;
    else
      data_o[100] <= next_data_o[100];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[101] <= 0;
    else
      data_o[101] <= next_data_o[101];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[102] <= 0;
    else
      data_o[102] <= next_data_o[102];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[103] <= 0;
    else
      data_o[103] <= next_data_o[103];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[104] <= 0;
    else
      data_o[104] <= next_data_o[104];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[105] <= 0;
    else
      data_o[105] <= next_data_o[105];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[106] <= 0;
    else
      data_o[106] <= next_data_o[106];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[107] <= 0;
    else
      data_o[107] <= next_data_o[107];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[108] <= 0;
    else
      data_o[108] <= next_data_o[108];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[109] <= 0;
    else
      data_o[109] <= next_data_o[109];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[10] <= 0;
    else
      data_o[10] <= next_data_o[10];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[110] <= 0;
    else
      data_o[110] <= next_data_o[110];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[111] <= 0;
    else
      data_o[111] <= next_data_o[111];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[112] <= 0;
    else
      data_o[112] <= next_data_o[112];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[113] <= 0;
    else
      data_o[113] <= next_data_o[113];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[114] <= 0;
    else
      data_o[114] <= next_data_o[114];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[115] <= 0;
    else
      data_o[115] <= next_data_o[115];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[116] <= 0;
    else
      data_o[116] <= next_data_o[116];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[117] <= 0;
    else
      data_o[117] <= next_data_o[117];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[118] <= 0;
    else
      data_o[118] <= next_data_o[118];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[119] <= 0;
    else
      data_o[119] <= next_data_o[119];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[11] <= 0;
    else
      data_o[11] <= next_data_o[11];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[120] <= 0;
    else
      data_o[120] <= next_data_o[120];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[121] <= 0;
    else
      data_o[121] <= next_data_o[121];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[122] <= 0;
    else
      data_o[122] <= next_data_o[122];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[123] <= 0;
    else
      data_o[123] <= next_data_o[123];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[124] <= 0;
    else
      data_o[124] <= next_data_o[124];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[125] <= 0;
    else
      data_o[125] <= next_data_o[125];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[126] <= 0;
    else
      data_o[126] <= next_data_o[126];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[127] <= 0;
    else
      data_o[127] <= next_data_o[127];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[12] <= 0;
    else
      data_o[12] <= next_data_o[12];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[13] <= 0;
    else
      data_o[13] <= next_data_o[13];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[14] <= 0;
    else
      data_o[14] <= next_data_o[14];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[15] <= 0;
    else
      data_o[15] <= next_data_o[15];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[16] <= 0;
    else
      data_o[16] <= next_data_o[16];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[17] <= 0;
    else
      data_o[17] <= next_data_o[17];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[18] <= 0;
    else
      data_o[18] <= next_data_o[18];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[19] <= 0;
    else
      data_o[19] <= next_data_o[19];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[1] <= 0;
    else
      data_o[1] <= next_data_o[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[20] <= 0;
    else
      data_o[20] <= next_data_o[20];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[21] <= 0;
    else
      data_o[21] <= next_data_o[21];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[22] <= 0;
    else
      data_o[22] <= next_data_o[22];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[23] <= 0;
    else
      data_o[23] <= next_data_o[23];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[24] <= 0;
    else
      data_o[24] <= next_data_o[24];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[25] <= 0;
    else
      data_o[25] <= next_data_o[25];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[26] <= 0;
    else
      data_o[26] <= next_data_o[26];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[27] <= 0;
    else
      data_o[27] <= next_data_o[27];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[28] <= 0;
    else
      data_o[28] <= next_data_o[28];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[29] <= 0;
    else
      data_o[29] <= next_data_o[29];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[2] <= 0;
    else
      data_o[2] <= next_data_o[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[30] <= 0;
    else
      data_o[30] <= next_data_o[30];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[31] <= 0;
    else
      data_o[31] <= next_data_o[31];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[32] <= 0;
    else
      data_o[32] <= next_data_o[32];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[33] <= 0;
    else
      data_o[33] <= next_data_o[33];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[34] <= 0;
    else
      data_o[34] <= next_data_o[34];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[35] <= 0;
    else
      data_o[35] <= next_data_o[35];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[36] <= 0;
    else
      data_o[36] <= next_data_o[36];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[37] <= 0;
    else
      data_o[37] <= next_data_o[37];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[38] <= 0;
    else
      data_o[38] <= next_data_o[38];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[39] <= 0;
    else
      data_o[39] <= next_data_o[39];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[3] <= 0;
    else
      data_o[3] <= next_data_o[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[40] <= 0;
    else
      data_o[40] <= next_data_o[40];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[41] <= 0;
    else
      data_o[41] <= next_data_o[41];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[42] <= 0;
    else
      data_o[42] <= next_data_o[42];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[43] <= 0;
    else
      data_o[43] <= next_data_o[43];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[44] <= 0;
    else
      data_o[44] <= next_data_o[44];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[45] <= 0;
    else
      data_o[45] <= next_data_o[45];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[46] <= 0;
    else
      data_o[46] <= next_data_o[46];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[47] <= 0;
    else
      data_o[47] <= next_data_o[47];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[48] <= 0;
    else
      data_o[48] <= next_data_o[48];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[49] <= 0;
    else
      data_o[49] <= next_data_o[49];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[4] <= 0;
    else
      data_o[4] <= next_data_o[4];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[50] <= 0;
    else
      data_o[50] <= next_data_o[50];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[51] <= 0;
    else
      data_o[51] <= next_data_o[51];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[52] <= 0;
    else
      data_o[52] <= next_data_o[52];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[53] <= 0;
    else
      data_o[53] <= next_data_o[53];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[54] <= 0;
    else
      data_o[54] <= next_data_o[54];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[55] <= 0;
    else
      data_o[55] <= next_data_o[55];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[56] <= 0;
    else
      data_o[56] <= next_data_o[56];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[57] <= 0;
    else
      data_o[57] <= next_data_o[57];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[58] <= 0;
    else
      data_o[58] <= next_data_o[58];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[59] <= 0;
    else
      data_o[59] <= next_data_o[59];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[5] <= 0;
    else
      data_o[5] <= next_data_o[5];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[60] <= 0;
    else
      data_o[60] <= next_data_o[60];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[61] <= 0;
    else
      data_o[61] <= next_data_o[61];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[62] <= 0;
    else
      data_o[62] <= next_data_o[62];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[63] <= 0;
    else
      data_o[63] <= next_data_o[63];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[64] <= 0;
    else
      data_o[64] <= next_data_o[64];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[65] <= 0;
    else
      data_o[65] <= next_data_o[65];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[66] <= 0;
    else
      data_o[66] <= next_data_o[66];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[67] <= 0;
    else
      data_o[67] <= next_data_o[67];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[68] <= 0;
    else
      data_o[68] <= next_data_o[68];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[69] <= 0;
    else
      data_o[69] <= next_data_o[69];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[6] <= 0;
    else
      data_o[6] <= next_data_o[6];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[70] <= 0;
    else
      data_o[70] <= next_data_o[70];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[71] <= 0;
    else
      data_o[71] <= next_data_o[71];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[72] <= 0;
    else
      data_o[72] <= next_data_o[72];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[73] <= 0;
    else
      data_o[73] <= next_data_o[73];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[74] <= 0;
    else
      data_o[74] <= next_data_o[74];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[75] <= 0;
    else
      data_o[75] <= next_data_o[75];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[76] <= 0;
    else
      data_o[76] <= next_data_o[76];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[77] <= 0;
    else
      data_o[77] <= next_data_o[77];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[78] <= 0;
    else
      data_o[78] <= next_data_o[78];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[79] <= 0;
    else
      data_o[79] <= next_data_o[79];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[7] <= 0;
    else
      data_o[7] <= next_data_o[7];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[80] <= 0;
    else
      data_o[80] <= next_data_o[80];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[81] <= 0;
    else
      data_o[81] <= next_data_o[81];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[82] <= 0;
    else
      data_o[82] <= next_data_o[82];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[83] <= 0;
    else
      data_o[83] <= next_data_o[83];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[84] <= 0;
    else
      data_o[84] <= next_data_o[84];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[85] <= 0;
    else
      data_o[85] <= next_data_o[85];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[86] <= 0;
    else
      data_o[86] <= next_data_o[86];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[87] <= 0;
    else
      data_o[87] <= next_data_o[87];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[88] <= 0;
    else
      data_o[88] <= next_data_o[88];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[89] <= 0;
    else
      data_o[89] <= next_data_o[89];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[8] <= 0;
    else
      data_o[8] <= next_data_o[8];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[90] <= 0;
    else
      data_o[90] <= next_data_o[90];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[91] <= 0;
    else
      data_o[91] <= next_data_o[91];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[92] <= 0;
    else
      data_o[92] <= next_data_o[92];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[93] <= 0;
    else
      data_o[93] <= next_data_o[93];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[94] <= 0;
    else
      data_o[94] <= next_data_o[94];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[95] <= 0;
    else
      data_o[95] <= next_data_o[95];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[96] <= 0;
    else
      data_o[96] <= next_data_o[96];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[97] <= 0;
    else
      data_o[97] <= next_data_o[97];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[98] <= 0;
    else
      data_o[98] <= next_data_o[98];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[99] <= 0;
    else
      data_o[99] <= next_data_o[99];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[9] <= 0;
    else
      data_o[9] <= next_data_o[9];
  reg \data_reg_reg[100] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[100]  <= 0;
    else
      \data_reg_reg[100]  <= next_data_reg[100];
  assign data_reg[100] = \data_reg_reg[100] ;
  reg \data_reg_reg[101] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[101]  <= 0;
    else
      \data_reg_reg[101]  <= next_data_reg[101];
  assign data_reg[101] = \data_reg_reg[101] ;
  reg \data_reg_reg[102] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[102]  <= 0;
    else
      \data_reg_reg[102]  <= next_data_reg[102];
  assign data_reg[102] = \data_reg_reg[102] ;
  reg \data_reg_reg[103] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[103]  <= 0;
    else
      \data_reg_reg[103]  <= next_data_reg[103];
  assign data_reg[103] = \data_reg_reg[103] ;
  reg \data_reg_reg[104] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[104]  <= 0;
    else
      \data_reg_reg[104]  <= next_data_reg[104];
  assign data_reg[104] = \data_reg_reg[104] ;
  reg \data_reg_reg[105] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[105]  <= 0;
    else
      \data_reg_reg[105]  <= next_data_reg[105];
  assign data_reg[105] = \data_reg_reg[105] ;
  reg \data_reg_reg[106] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[106]  <= 0;
    else
      \data_reg_reg[106]  <= next_data_reg[106];
  assign data_reg[106] = \data_reg_reg[106] ;
  reg \data_reg_reg[107] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[107]  <= 0;
    else
      \data_reg_reg[107]  <= next_data_reg[107];
  assign data_reg[107] = \data_reg_reg[107] ;
  reg \data_reg_reg[108] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[108]  <= 0;
    else
      \data_reg_reg[108]  <= next_data_reg[108];
  assign data_reg[108] = \data_reg_reg[108] ;
  reg \data_reg_reg[109] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[109]  <= 0;
    else
      \data_reg_reg[109]  <= next_data_reg[109];
  assign data_reg[109] = \data_reg_reg[109] ;
  reg \data_reg_reg[110] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[110]  <= 0;
    else
      \data_reg_reg[110]  <= next_data_reg[110];
  assign data_reg[110] = \data_reg_reg[110] ;
  reg \data_reg_reg[111] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[111]  <= 0;
    else
      \data_reg_reg[111]  <= next_data_reg[111];
  assign data_reg[111] = \data_reg_reg[111] ;
  reg \data_reg_reg[112] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[112]  <= 0;
    else
      \data_reg_reg[112]  <= next_data_reg[112];
  assign data_reg[112] = \data_reg_reg[112] ;
  reg \data_reg_reg[113] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[113]  <= 0;
    else
      \data_reg_reg[113]  <= next_data_reg[113];
  assign data_reg[113] = \data_reg_reg[113] ;
  reg \data_reg_reg[114] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[114]  <= 0;
    else
      \data_reg_reg[114]  <= next_data_reg[114];
  assign data_reg[114] = \data_reg_reg[114] ;
  reg \data_reg_reg[115] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[115]  <= 0;
    else
      \data_reg_reg[115]  <= next_data_reg[115];
  assign data_reg[115] = \data_reg_reg[115] ;
  reg \data_reg_reg[116] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[116]  <= 0;
    else
      \data_reg_reg[116]  <= next_data_reg[116];
  assign data_reg[116] = \data_reg_reg[116] ;
  reg \data_reg_reg[117] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[117]  <= 0;
    else
      \data_reg_reg[117]  <= next_data_reg[117];
  assign data_reg[117] = \data_reg_reg[117] ;
  reg \data_reg_reg[118] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[118]  <= 0;
    else
      \data_reg_reg[118]  <= next_data_reg[118];
  assign data_reg[118] = \data_reg_reg[118] ;
  reg \data_reg_reg[119] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[119]  <= 0;
    else
      \data_reg_reg[119]  <= next_data_reg[119];
  assign data_reg[119] = \data_reg_reg[119] ;
  reg \data_reg_reg[120] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[120]  <= 0;
    else
      \data_reg_reg[120]  <= next_data_reg[120];
  assign data_reg[120] = \data_reg_reg[120] ;
  reg \data_reg_reg[121] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[121]  <= 0;
    else
      \data_reg_reg[121]  <= next_data_reg[121];
  assign data_reg[121] = \data_reg_reg[121] ;
  reg \data_reg_reg[122] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[122]  <= 0;
    else
      \data_reg_reg[122]  <= next_data_reg[122];
  assign data_reg[122] = \data_reg_reg[122] ;
  reg \data_reg_reg[123] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[123]  <= 0;
    else
      \data_reg_reg[123]  <= next_data_reg[123];
  assign data_reg[123] = \data_reg_reg[123] ;
  reg \data_reg_reg[124] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[124]  <= 0;
    else
      \data_reg_reg[124]  <= next_data_reg[124];
  assign data_reg[124] = \data_reg_reg[124] ;
  reg \data_reg_reg[125] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[125]  <= 0;
    else
      \data_reg_reg[125]  <= next_data_reg[125];
  assign data_reg[125] = \data_reg_reg[125] ;
  reg \data_reg_reg[126] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[126]  <= 0;
    else
      \data_reg_reg[126]  <= next_data_reg[126];
  assign data_reg[126] = \data_reg_reg[126] ;
  reg \data_reg_reg[127] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[127]  <= 0;
    else
      \data_reg_reg[127]  <= next_data_reg[127];
  assign data_reg[127] = \data_reg_reg[127] ;
  reg \data_reg_reg[32] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[32]  <= 0;
    else
      \data_reg_reg[32]  <= next_data_reg[32];
  assign data_reg[32] = \data_reg_reg[32] ;
  reg \data_reg_reg[33] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[33]  <= 0;
    else
      \data_reg_reg[33]  <= next_data_reg[33];
  assign data_reg[33] = \data_reg_reg[33] ;
  reg \data_reg_reg[34] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[34]  <= 0;
    else
      \data_reg_reg[34]  <= next_data_reg[34];
  assign data_reg[34] = \data_reg_reg[34] ;
  reg \data_reg_reg[35] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[35]  <= 0;
    else
      \data_reg_reg[35]  <= next_data_reg[35];
  assign data_reg[35] = \data_reg_reg[35] ;
  reg \data_reg_reg[36] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[36]  <= 0;
    else
      \data_reg_reg[36]  <= next_data_reg[36];
  assign data_reg[36] = \data_reg_reg[36] ;
  reg \data_reg_reg[37] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[37]  <= 0;
    else
      \data_reg_reg[37]  <= next_data_reg[37];
  assign data_reg[37] = \data_reg_reg[37] ;
  reg \data_reg_reg[38] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[38]  <= 0;
    else
      \data_reg_reg[38]  <= next_data_reg[38];
  assign data_reg[38] = \data_reg_reg[38] ;
  reg \data_reg_reg[39] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[39]  <= 0;
    else
      \data_reg_reg[39]  <= next_data_reg[39];
  assign data_reg[39] = \data_reg_reg[39] ;
  reg \data_reg_reg[40] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[40]  <= 0;
    else
      \data_reg_reg[40]  <= next_data_reg[40];
  assign data_reg[40] = \data_reg_reg[40] ;
  reg \data_reg_reg[41] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[41]  <= 0;
    else
      \data_reg_reg[41]  <= next_data_reg[41];
  assign data_reg[41] = \data_reg_reg[41] ;
  reg \data_reg_reg[42] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[42]  <= 0;
    else
      \data_reg_reg[42]  <= next_data_reg[42];
  assign data_reg[42] = \data_reg_reg[42] ;
  reg \data_reg_reg[43] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[43]  <= 0;
    else
      \data_reg_reg[43]  <= next_data_reg[43];
  assign data_reg[43] = \data_reg_reg[43] ;
  reg \data_reg_reg[44] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[44]  <= 0;
    else
      \data_reg_reg[44]  <= next_data_reg[44];
  assign data_reg[44] = \data_reg_reg[44] ;
  reg \data_reg_reg[45] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[45]  <= 0;
    else
      \data_reg_reg[45]  <= next_data_reg[45];
  assign data_reg[45] = \data_reg_reg[45] ;
  reg \data_reg_reg[46] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[46]  <= 0;
    else
      \data_reg_reg[46]  <= next_data_reg[46];
  assign data_reg[46] = \data_reg_reg[46] ;
  reg \data_reg_reg[47] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[47]  <= 0;
    else
      \data_reg_reg[47]  <= next_data_reg[47];
  assign data_reg[47] = \data_reg_reg[47] ;
  reg \data_reg_reg[48] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[48]  <= 0;
    else
      \data_reg_reg[48]  <= next_data_reg[48];
  assign data_reg[48] = \data_reg_reg[48] ;
  reg \data_reg_reg[49] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[49]  <= 0;
    else
      \data_reg_reg[49]  <= next_data_reg[49];
  assign data_reg[49] = \data_reg_reg[49] ;
  reg \data_reg_reg[50] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[50]  <= 0;
    else
      \data_reg_reg[50]  <= next_data_reg[50];
  assign data_reg[50] = \data_reg_reg[50] ;
  reg \data_reg_reg[51] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[51]  <= 0;
    else
      \data_reg_reg[51]  <= next_data_reg[51];
  assign data_reg[51] = \data_reg_reg[51] ;
  reg \data_reg_reg[52] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[52]  <= 0;
    else
      \data_reg_reg[52]  <= next_data_reg[52];
  assign data_reg[52] = \data_reg_reg[52] ;
  reg \data_reg_reg[53] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[53]  <= 0;
    else
      \data_reg_reg[53]  <= next_data_reg[53];
  assign data_reg[53] = \data_reg_reg[53] ;
  reg \data_reg_reg[54] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[54]  <= 0;
    else
      \data_reg_reg[54]  <= next_data_reg[54];
  assign data_reg[54] = \data_reg_reg[54] ;
  reg \data_reg_reg[55] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[55]  <= 0;
    else
      \data_reg_reg[55]  <= next_data_reg[55];
  assign data_reg[55] = \data_reg_reg[55] ;
  reg \data_reg_reg[56] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[56]  <= 0;
    else
      \data_reg_reg[56]  <= next_data_reg[56];
  assign data_reg[56] = \data_reg_reg[56] ;
  reg \data_reg_reg[57] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[57]  <= 0;
    else
      \data_reg_reg[57]  <= next_data_reg[57];
  assign data_reg[57] = \data_reg_reg[57] ;
  reg \data_reg_reg[58] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[58]  <= 0;
    else
      \data_reg_reg[58]  <= next_data_reg[58];
  assign data_reg[58] = \data_reg_reg[58] ;
  reg \data_reg_reg[59] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[59]  <= 0;
    else
      \data_reg_reg[59]  <= next_data_reg[59];
  assign data_reg[59] = \data_reg_reg[59] ;
  reg \data_reg_reg[60] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[60]  <= 0;
    else
      \data_reg_reg[60]  <= next_data_reg[60];
  assign data_reg[60] = \data_reg_reg[60] ;
  reg \data_reg_reg[61] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[61]  <= 0;
    else
      \data_reg_reg[61]  <= next_data_reg[61];
  assign data_reg[61] = \data_reg_reg[61] ;
  reg \data_reg_reg[62] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[62]  <= 0;
    else
      \data_reg_reg[62]  <= next_data_reg[62];
  assign data_reg[62] = \data_reg_reg[62] ;
  reg \data_reg_reg[63] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[63]  <= 0;
    else
      \data_reg_reg[63]  <= next_data_reg[63];
  assign data_reg[63] = \data_reg_reg[63] ;
  reg \data_reg_reg[64] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[64]  <= 0;
    else
      \data_reg_reg[64]  <= next_data_reg[64];
  assign data_reg[64] = \data_reg_reg[64] ;
  reg \data_reg_reg[65] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[65]  <= 0;
    else
      \data_reg_reg[65]  <= next_data_reg[65];
  assign data_reg[65] = \data_reg_reg[65] ;
  reg \data_reg_reg[66] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[66]  <= 0;
    else
      \data_reg_reg[66]  <= next_data_reg[66];
  assign data_reg[66] = \data_reg_reg[66] ;
  reg \data_reg_reg[67] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[67]  <= 0;
    else
      \data_reg_reg[67]  <= next_data_reg[67];
  assign data_reg[67] = \data_reg_reg[67] ;
  reg \data_reg_reg[68] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[68]  <= 0;
    else
      \data_reg_reg[68]  <= next_data_reg[68];
  assign data_reg[68] = \data_reg_reg[68] ;
  reg \data_reg_reg[69] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[69]  <= 0;
    else
      \data_reg_reg[69]  <= next_data_reg[69];
  assign data_reg[69] = \data_reg_reg[69] ;
  reg \data_reg_reg[70] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[70]  <= 0;
    else
      \data_reg_reg[70]  <= next_data_reg[70];
  assign data_reg[70] = \data_reg_reg[70] ;
  reg \data_reg_reg[71] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[71]  <= 0;
    else
      \data_reg_reg[71]  <= next_data_reg[71];
  assign data_reg[71] = \data_reg_reg[71] ;
  reg \data_reg_reg[72] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[72]  <= 0;
    else
      \data_reg_reg[72]  <= next_data_reg[72];
  assign data_reg[72] = \data_reg_reg[72] ;
  reg \data_reg_reg[73] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[73]  <= 0;
    else
      \data_reg_reg[73]  <= next_data_reg[73];
  assign data_reg[73] = \data_reg_reg[73] ;
  reg \data_reg_reg[74] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[74]  <= 0;
    else
      \data_reg_reg[74]  <= next_data_reg[74];
  assign data_reg[74] = \data_reg_reg[74] ;
  reg \data_reg_reg[75] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[75]  <= 0;
    else
      \data_reg_reg[75]  <= next_data_reg[75];
  assign data_reg[75] = \data_reg_reg[75] ;
  reg \data_reg_reg[76] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[76]  <= 0;
    else
      \data_reg_reg[76]  <= next_data_reg[76];
  assign data_reg[76] = \data_reg_reg[76] ;
  reg \data_reg_reg[77] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[77]  <= 0;
    else
      \data_reg_reg[77]  <= next_data_reg[77];
  assign data_reg[77] = \data_reg_reg[77] ;
  reg \data_reg_reg[78] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[78]  <= 0;
    else
      \data_reg_reg[78]  <= next_data_reg[78];
  assign data_reg[78] = \data_reg_reg[78] ;
  reg \data_reg_reg[79] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[79]  <= 0;
    else
      \data_reg_reg[79]  <= next_data_reg[79];
  assign data_reg[79] = \data_reg_reg[79] ;
  reg \data_reg_reg[80] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[80]  <= 0;
    else
      \data_reg_reg[80]  <= next_data_reg[80];
  assign data_reg[80] = \data_reg_reg[80] ;
  reg \data_reg_reg[81] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[81]  <= 0;
    else
      \data_reg_reg[81]  <= next_data_reg[81];
  assign data_reg[81] = \data_reg_reg[81] ;
  reg \data_reg_reg[82] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[82]  <= 0;
    else
      \data_reg_reg[82]  <= next_data_reg[82];
  assign data_reg[82] = \data_reg_reg[82] ;
  reg \data_reg_reg[83] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[83]  <= 0;
    else
      \data_reg_reg[83]  <= next_data_reg[83];
  assign data_reg[83] = \data_reg_reg[83] ;
  reg \data_reg_reg[84] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[84]  <= 0;
    else
      \data_reg_reg[84]  <= next_data_reg[84];
  assign data_reg[84] = \data_reg_reg[84] ;
  reg \data_reg_reg[85] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[85]  <= 0;
    else
      \data_reg_reg[85]  <= next_data_reg[85];
  assign data_reg[85] = \data_reg_reg[85] ;
  reg \data_reg_reg[86] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[86]  <= 0;
    else
      \data_reg_reg[86]  <= next_data_reg[86];
  assign data_reg[86] = \data_reg_reg[86] ;
  reg \data_reg_reg[87] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[87]  <= 0;
    else
      \data_reg_reg[87]  <= next_data_reg[87];
  assign data_reg[87] = \data_reg_reg[87] ;
  reg \data_reg_reg[88] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[88]  <= 0;
    else
      \data_reg_reg[88]  <= next_data_reg[88];
  assign data_reg[88] = \data_reg_reg[88] ;
  reg \data_reg_reg[89] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[89]  <= 0;
    else
      \data_reg_reg[89]  <= next_data_reg[89];
  assign data_reg[89] = \data_reg_reg[89] ;
  reg \data_reg_reg[90] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[90]  <= 0;
    else
      \data_reg_reg[90]  <= next_data_reg[90];
  assign data_reg[90] = \data_reg_reg[90] ;
  reg \data_reg_reg[91] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[91]  <= 0;
    else
      \data_reg_reg[91]  <= next_data_reg[91];
  assign data_reg[91] = \data_reg_reg[91] ;
  reg \data_reg_reg[92] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[92]  <= 0;
    else
      \data_reg_reg[92]  <= next_data_reg[92];
  assign data_reg[92] = \data_reg_reg[92] ;
  reg \data_reg_reg[93] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[93]  <= 0;
    else
      \data_reg_reg[93]  <= next_data_reg[93];
  assign data_reg[93] = \data_reg_reg[93] ;
  reg \data_reg_reg[94] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[94]  <= 0;
    else
      \data_reg_reg[94]  <= next_data_reg[94];
  assign data_reg[94] = \data_reg_reg[94] ;
  reg \data_reg_reg[95] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[95]  <= 0;
    else
      \data_reg_reg[95]  <= next_data_reg[95];
  assign data_reg[95] = \data_reg_reg[95] ;
  reg \data_reg_reg[96] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[96]  <= 0;
    else
      \data_reg_reg[96]  <= next_data_reg[96];
  assign data_reg[96] = \data_reg_reg[96] ;
  reg \data_reg_reg[97] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[97]  <= 0;
    else
      \data_reg_reg[97]  <= next_data_reg[97];
  assign data_reg[97] = \data_reg_reg[97] ;
  reg \data_reg_reg[98] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[98]  <= 0;
    else
      \data_reg_reg[98]  <= next_data_reg[98];
  assign data_reg[98] = \data_reg_reg[98] ;
  reg \data_reg_reg[99] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      \data_reg_reg[99]  <= 0;
    else
      \data_reg_reg[99]  <= next_data_reg[99];
  assign data_reg[99] = \data_reg_reg[99] ;
  always @(posedge clk or negedge reset)
    if (!reset)
      ready_o <= 0;
    else
      ready_o <= next_ready_o;
  always @(posedge clk or negedge reset)
    if (!reset)
      state[0] <= 0;
    else
      state[0] <= next_state[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[1] <= 0;
    else
      state[1] <= next_state[1];
  word_mixcolum w1 (
    .in(mix_word),
    .outx(outx),
    .outy(outy)
  );
  assign data_i_var = data_i;
  assign data_o_reg = data_o;
endmodule

module sbox(clk, reset, data_i, decrypt_i, data_o);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire [3:0] ah;
  wire [3:0] ah2;
  reg [3:0] ah_reg;
  reg [3:0] alph;
  input clk;
  input [7:0] data_i;
  output [7:0] data_o;
  input decrypt_i;
  wire first_mux_aB;
  wire [3:0] first_mux_ah_t;
  wire [7:0] first_mux_data_var;
  wire [3:0] intermediate_to_invert_var;
  reg [3:0] inversion_to_invert_var;
  wire [3:0] next_ah_reg;
  wire [3:0] next_alph;
  wire [3:0] next_to_invert;
  input reset;
  wire [3:0] square1_ah_t;
  wire [3:0] sum1_alph_t;
  wire [3:0] to_invert;
  assign _171_ = ~decrypt_i;
  assign _172_ = ~data_i[4];
  assign _173_ = ~data_i[1];
  assign _174_ = data_i[6] ^ data_i[3];
  assign _175_ = _174_ ^ _173_;
  assign _176_ = _171_ ? _172_ : _175_;
  assign _177_ = ~_176_;
  assign _178_ = ~data_i[6];
  assign _179_ = ~data_i[3];
  assign _180_ = data_i[0] ^ data_i[5];
  assign _181_ = _180_ ^ _179_;
  assign _182_ = _171_ ? _178_ : _181_;
  assign _183_ = _182_ ^ _177_;
  assign _184_ = ~data_i[5];
  assign _185_ = data_i[2] ^ data_i[7];
  assign _186_ = _185_ ^ _172_;
  assign _187_ = _171_ ? _184_ : _186_;
  assign _188_ = ~_187_;
  assign _189_ = _188_ ^ _183_;
  assign ah[0] = ~_189_;
  assign _190_ = ~_183_;
  assign _191_ = ~data_i[0];
  assign _192_ = _174_ ^ _191_;
  assign _193_ = _171_ ? _173_ : _192_;
  assign _194_ = ~_193_;
  assign _195_ = ~data_i[7];
  assign _196_ = data_i[4] ^ data_i[1];
  assign _197_ = _196_ ^ _178_;
  assign _198_ = _171_ ? _195_ : _197_;
  assign _199_ = _198_ ^ _194_;
  assign _200_ = _199_ ^ _190_;
  assign ah[1] = ~_200_;
  assign _201_ = _198_ ^ _188_;
  assign ah[3] = ~_201_;
  assign _202_ = ~data_i[2];
  assign _203_ = _196_ ^ data_i[7];
  assign _204_ = _171_ ? _202_ : _203_;
  assign _205_ = _204_ ^ ah[3];
  assign _206_ = _180_ ^ _202_;
  assign _207_ = _171_ ? _179_ : _206_;
  assign ah[2] = _207_ ^ _205_;
  assign _208_ = ~alph[0];
  assign _209_ = inversion_to_invert_var[1] & inversion_to_invert_var[2];
  assign _210_ = ~inversion_to_invert_var[3];
  assign _211_ = inversion_to_invert_var[1] ^ inversion_to_invert_var[2];
  assign _212_ = _211_ ^ _210_;
  assign _213_ = _209_ & inversion_to_invert_var[3];
  assign _214_ = _213_ ^ _212_;
  assign _215_ = _214_ ^ inversion_to_invert_var[0];
  assign _216_ = inversion_to_invert_var[0] & inversion_to_invert_var[2];
  assign _217_ = _216_ ^ _215_;
  assign _218_ = _217_ ^ _209_;
  assign _219_ = inversion_to_invert_var[0] & inversion_to_invert_var[1];
  assign _220_ = _219_ & inversion_to_invert_var[2];
  assign _221_ = _220_ ^ _218_;
  assign _222_ = _221_ | _208_;
  assign _223_ = inversion_to_invert_var[0] & inversion_to_invert_var[3];
  assign _224_ = _223_ ^ _214_;
  assign _225_ = inversion_to_invert_var[3] & inversion_to_invert_var[1];
  assign _000_ = _225_ ^ _224_;
  assign _001_ = inversion_to_invert_var[3] & inversion_to_invert_var[2];
  assign _002_ = _001_ ^ _000_;
  assign _003_ = ~_002_;
  assign _004_ = _003_ & alph[1];
  assign _005_ = _004_ ^ _222_;
  assign _006_ = inversion_to_invert_var[0] ? inversion_to_invert_var[1] : inversion_to_invert_var[2];
  assign _007_ = _006_ ^ _210_;
  assign _008_ = _007_ ^ _223_;
  assign _009_ = _216_ & inversion_to_invert_var[3];
  assign _010_ = _009_ ^ _008_;
  assign _011_ = ~_010_;
  assign _012_ = _011_ & alph[2];
  assign _013_ = _012_ ^ _005_;
  assign _014_ = ~alph[3];
  assign _015_ = ~_209_;
  assign _016_ = _219_ ^ _216_;
  assign _017_ = _016_ ^ _015_;
  assign _018_ = _017_ ^ inversion_to_invert_var[3];
  assign _019_ = _018_ ^ _225_;
  assign _020_ = _219_ & inversion_to_invert_var[3];
  assign _021_ = _020_ ^ _019_;
  assign _022_ = _021_ | _014_;
  assign _023_ = _022_ ^ _013_;
  assign _024_ = _217_ ^ _015_;
  assign _025_ = _220_ ^ _024_;
  assign _026_ = _025_ & ah_reg[0];
  assign _027_ = ~ah_reg[3];
  assign _028_ = _021_ | _027_;
  assign _029_ = _028_ ^ _026_;
  assign _030_ = _011_ & ah_reg[2];
  assign _031_ = _030_ ^ _029_;
  assign _032_ = _003_ & ah_reg[1];
  assign _033_ = ~_032_;
  assign _034_ = _033_ ^ _031_;
  assign _035_ = _034_ ^ _023_;
  assign _036_ = _021_ | _208_;
  assign _037_ = _002_ ^ _221_;
  assign _038_ = _037_ & alph[1];
  assign _039_ = _038_ ^ _036_;
  assign _040_ = _010_ ^ _002_;
  assign _041_ = _040_ & alph[2];
  assign _042_ = _041_ ^ _039_;
  assign _043_ = _021_ ^ _010_;
  assign _044_ = _043_ & alph[3];
  assign _045_ = _044_ ^ _042_;
  assign _046_ = _221_ | _027_;
  assign _047_ = ~_021_;
  assign _048_ = _047_ & ah_reg[2];
  assign _049_ = _048_ ^ _046_;
  assign _050_ = _011_ & ah_reg[1];
  assign _051_ = _050_ ^ _049_;
  assign _052_ = ah_reg[3] ^ ah_reg[0];
  assign _053_ = _052_ & _003_;
  assign _054_ = _053_ ^ _051_;
  assign _055_ = _054_ ^ _045_;
  assign _056_ = _032_ ^ _031_;
  assign _057_ = ~ah_reg[1];
  assign _058_ = _221_ | _057_;
  assign _059_ = _052_ & _047_;
  assign _060_ = _059_ ^ _058_;
  assign _061_ = ah_reg[2] ^ ah_reg[3];
  assign _062_ = _061_ & _011_;
  assign _063_ = _062_ ^ _060_;
  assign _064_ = ah_reg[1] ^ ah_reg[2];
  assign _065_ = _064_ & _003_;
  assign _066_ = _065_ ^ _063_;
  assign _067_ = _066_ ^ _056_;
  assign _068_ = _067_ ^ _055_;
  assign _069_ = _002_ | _208_;
  assign _070_ = _011_ & alph[1];
  assign _071_ = _070_ ^ _069_;
  assign _072_ = ~alph[2];
  assign _073_ = _021_ | _072_;
  assign _074_ = _073_ ^ _071_;
  assign _075_ = _037_ & alph[3];
  assign _076_ = _075_ ^ _074_;
  assign _077_ = _076_ ^ _068_;
  assign _078_ = _010_ | _208_;
  assign _079_ = _047_ & alph[1];
  assign _080_ = _079_ ^ _078_;
  assign _081_ = _037_ & alph[2];
  assign _082_ = _081_ ^ _080_;
  assign _083_ = _040_ & alph[3];
  assign _084_ = _083_ ^ _082_;
  assign _085_ = _084_ ^ _067_;
  assign _086_ = ~_085_;
  assign _087_ = _086_ ^ _077_;
  assign _088_ = _087_ ^ _035_;
  assign _089_ = _084_ ^ _055_;
  assign _090_ = _089_ ^ _076_;
  assign _091_ = _090_ ^ _034_;
  assign _092_ = _085_ ^ _054_;
  assign _093_ = _092_ ^ _091_;
  assign _094_ = _093_ ^ _088_;
  assign data_o[0] = decrypt_i ? _035_ : _094_;
  assign _095_ = _067_ ^ _054_;
  assign _096_ = ~_095_;
  assign _097_ = _095_ ^ _035_;
  assign _098_ = _097_ ^ _085_;
  assign _099_ = _098_ ^ _093_;
  assign data_o[1] = decrypt_i ? _096_ : _099_;
  assign _100_ = _066_ ^ _034_;
  assign _101_ = _045_ ^ _035_;
  assign _102_ = _101_ ^ _093_;
  assign data_o[2] = decrypt_i ? _068_ : _102_;
  assign _103_ = _100_ ^ _045_;
  assign _104_ = _025_ & ah_reg[2];
  assign _105_ = _021_ | _057_;
  assign _106_ = _105_ ^ _104_;
  assign _107_ = _052_ & _011_;
  assign _108_ = _107_ ^ _106_;
  assign _109_ = _061_ & _003_;
  assign _110_ = _109_ ^ _108_;
  assign _111_ = _110_ ^ _103_;
  assign _112_ = ~_111_;
  assign _113_ = _097_ ^ _092_;
  assign _114_ = _111_ ^ _068_;
  assign _115_ = _114_ ^ _113_;
  assign data_o[3] = decrypt_i ? _112_ : _115_;
  assign _116_ = _097_ ^ _077_;
  assign _117_ = _116_ ^ _114_;
  assign data_o[4] = decrypt_i ? _077_ : _117_;
  assign _118_ = _114_ ^ _095_;
  assign _119_ = _118_ ^ _090_;
  assign data_o[5] = decrypt_i ? _086_ : _119_;
  assign _120_ = ~_091_;
  assign _121_ = _114_ ^ _091_;
  assign _122_ = _121_ ^ _090_;
  assign data_o[6] = decrypt_i ? _120_ : _122_;
  assign _123_ = _111_ ^ _087_;
  assign _124_ = _123_ ^ _093_;
  assign data_o[7] = decrypt_i ? _092_ : _124_;
  assign _125_ = _200_ ^ ah[2];
  assign _126_ = _185_ ^ _184_;
  assign _127_ = _171_ ? data_i[0] : _126_;
  assign _128_ = _127_ ^ _183_;
  assign _129_ = _128_ ^ _188_;
  assign _130_ = _129_ ^ _199_;
  assign _131_ = _130_ ^ _125_;
  assign _132_ = _129_ | _189_;
  assign _133_ = _204_ ^ _177_;
  assign _134_ = ~_133_;
  assign _135_ = _134_ & ah[1];
  assign _136_ = _135_ ^ _132_;
  assign _137_ = ~_199_;
  assign _138_ = ah[2] & _137_;
  assign _139_ = _138_ ^ _136_;
  assign _140_ = _204_ ^ _194_;
  assign _141_ = ~_140_;
  assign _142_ = _141_ & ah[3];
  assign _143_ = _142_ ^ _139_;
  assign intermediate_to_invert_var[0] = _143_ ^ _131_;
  assign _144_ = _189_ ^ _137_;
  assign _145_ = _140_ | _189_;
  assign _146_ = _133_ ^ _129_;
  assign _147_ = _146_ & ah[1];
  assign _148_ = _147_ ^ _145_;
  assign _149_ = _133_ ^ _199_;
  assign _150_ = _149_ & ah[2];
  assign _151_ = _150_ ^ _148_;
  assign _152_ = _140_ ^ _199_;
  assign _153_ = _152_ & ah[3];
  assign _154_ = _153_ ^ _151_;
  assign intermediate_to_invert_var[1] = _154_ ^ _144_;
  assign _155_ = _137_ & ah[0];
  assign _156_ = _140_ | _200_;
  assign _157_ = _156_ ^ _155_;
  assign _158_ = _146_ & ah[2];
  assign _159_ = _158_ ^ _157_;
  assign _160_ = _149_ & ah[3];
  assign _161_ = _160_ ^ _159_;
  assign intermediate_to_invert_var[2] = _161_ ^ _176_;
  assign _162_ = _200_ ^ ah[0];
  assign _163_ = _162_ ^ _134_;
  assign _164_ = _133_ | _189_;
  assign _165_ = _137_ & _183_;
  assign _166_ = _165_ ^ _164_;
  assign _167_ = _141_ & ah[2];
  assign _168_ = _167_ ^ _166_;
  assign _169_ = _146_ & ah[3];
  assign _170_ = _169_ ^ _168_;
  assign intermediate_to_invert_var[3] = _170_ ^ _163_;
  assign next_alph[0] = _129_ ^ _189_;
  assign next_alph[1] = _140_ ^ _200_;
  assign next_alph[2] = ah[2] ^ _137_;
  assign next_alph[3] = _133_ ^ _201_;
  always @(posedge clk or negedge reset)
    if (!reset)
      ah_reg[0] <= 0;
    else
      ah_reg[0] <= ah[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      ah_reg[1] <= 0;
    else
      ah_reg[1] <= ah[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      ah_reg[2] <= 0;
    else
      ah_reg[2] <= ah[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      ah_reg[3] <= 0;
    else
      ah_reg[3] <= ah[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      alph[0] <= 0;
    else
      alph[0] <= next_alph[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      alph[1] <= 0;
    else
      alph[1] <= next_alph[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      alph[2] <= 0;
    else
      alph[2] <= next_alph[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      alph[3] <= 0;
    else
      alph[3] <= next_alph[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      inversion_to_invert_var[0] <= 0;
    else
      inversion_to_invert_var[0] <= intermediate_to_invert_var[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      inversion_to_invert_var[1] <= 0;
    else
      inversion_to_invert_var[1] <= intermediate_to_invert_var[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      inversion_to_invert_var[2] <= 0;
    else
      inversion_to_invert_var[2] <= intermediate_to_invert_var[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      inversion_to_invert_var[3] <= 0;
    else
      inversion_to_invert_var[3] <= intermediate_to_invert_var[3];
  assign { ah2[3], ah2[1] } = ah[3:2];
  assign first_mux_aB = ah[3];
  assign first_mux_ah_t = ah;
  assign first_mux_data_var = data_i;
  assign next_ah_reg = ah;
  assign next_to_invert = intermediate_to_invert_var;
  assign square1_ah_t = { ah[3], ah2[2], ah[2], ah2[0] };
  assign sum1_alph_t = next_alph;
  assign to_invert = inversion_to_invert_var;
endmodule

module subbytes(clk, reset, start_i, decrypt_i, data_i, ready_o, data_o, sbox_data_o, sbox_data_i, sbox_decrypt_o);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  input clk;
  wire [7:0] \data_array[0] ;
  wire [7:0] \data_array[10] ;
  wire [7:0] \data_array[11] ;
  wire [7:0] \data_array[12] ;
  wire [7:0] \data_array[13] ;
  wire [7:0] \data_array[14] ;
  wire [7:0] \data_array[15] ;
  wire [7:0] \data_array[1] ;
  wire [7:0] \data_array[2] ;
  wire [7:0] \data_array[3] ;
  wire [7:0] \data_array[4] ;
  wire [7:0] \data_array[5] ;
  wire [7:0] \data_array[6] ;
  wire [7:0] \data_array[7] ;
  wire [7:0] \data_array[8] ;
  wire [7:0] \data_array[9] ;
  input [127:0] data_i;
  wire [127:0] data_i_var;
  output [127:0] data_o;
  reg [127:0] data_o;
  wire [127:0] data_reg;
  input decrypt_i;
  wire [127:0] next_data_reg;
  wire next_ready_o;
  wire [4:0] next_state;
  output ready_o;
  reg ready_o;
  input reset;
  input [7:0] sbox_data_i;
  output [7:0] sbox_data_o;
  output sbox_decrypt_o;
  input start_i;
  reg [4:0] state;
  assign _0447_ = ~state[3];
  assign _0448_ = ~state[2];
  assign _0449_ = ~state[0];
  assign _0450_ = ~state[1];
  assign _0451_ = _0450_ & _0449_;
  assign _0452_ = _0451_ & _0448_;
  assign _0453_ = _0452_ & _0447_;
  assign next_ready_o = _0453_ & state[4];
  assign _0454_ = state[1] | state[0];
  assign _0455_ = _0454_ | state[2];
  assign _0456_ = _0455_ | state[3];
  assign _0457_ = _0456_ | state[4];
  assign _0458_ = ~_0457_;
  assign _0459_ = _0458_ & data_o[0];
  assign _0460_ = decrypt_i ? data_o[96] : data_o[32];
  assign _0461_ = _0460_ & next_ready_o;
  assign _0462_ = _0461_ | _0459_;
  assign _0463_ = _0455_ ^ _0447_;
  assign _0464_ = _0454_ ^ _0448_;
  assign _0465_ = state[1] | _0449_;
  assign _0466_ = _0465_ | _0464_;
  assign _0467_ = _0466_ | _0463_;
  assign _0468_ = _0450_ | state[0];
  assign _0469_ = _0468_ | _0464_;
  assign _0470_ = _0469_ | _0463_;
  assign _0471_ = _0450_ | _0449_;
  assign _0472_ = _0471_ | _0464_;
  assign _0473_ = _0472_ | _0463_;
  assign _0474_ = _0455_ ^ state[3];
  assign _0475_ = _0454_ ^ state[2];
  assign _0476_ = _0471_ | _0475_;
  assign _0477_ = _0476_ | _0474_;
  assign _0478_ = _0468_ | _0475_;
  assign _0479_ = _0478_ | _0474_;
  assign _0480_ = _0465_ | _0475_;
  assign _0481_ = _0480_ | _0474_;
  assign _0482_ = _0472_ | _0474_;
  assign _0483_ = _0466_ | _0474_;
  assign _0484_ = _0469_ | _0474_;
  assign _0485_ = _0480_ | _0463_;
  assign _0486_ = _0478_ | _0463_;
  assign _0487_ = _0476_ | _0463_;
  assign _0488_ = _0453_ ? sbox_data_i[0] : data_o[0];
  assign next_data_reg[0] = _0453_ ? _0462_ : _0488_;
  assign _0489_ = _0458_ & data_o[100];
  assign _0490_ = decrypt_i ? data_o[68] : sbox_data_i[4];
  assign _0491_ = _0490_ & next_ready_o;
  assign _0492_ = _0491_ | _0489_;
  assign _0493_ = _0170_ ? data_o[100] : sbox_data_i[4];
  assign next_data_reg[100] = _0456_ ? _0493_ : _0492_;
  assign _0494_ = _0458_ & data_o[101];
  assign _0495_ = decrypt_i ? data_o[69] : sbox_data_i[5];
  assign _0496_ = _0495_ & next_ready_o;
  assign _0497_ = _0496_ | _0494_;
  assign _0498_ = _0170_ ? data_o[101] : sbox_data_i[5];
  assign next_data_reg[101] = _0456_ ? _0498_ : _0497_;
  assign _0499_ = _0458_ & data_o[102];
  assign _0500_ = decrypt_i ? data_o[70] : sbox_data_i[6];
  assign _0501_ = _0500_ & next_ready_o;
  assign _0502_ = _0501_ | _0499_;
  assign _0503_ = _0170_ ? data_o[102] : sbox_data_i[6];
  assign next_data_reg[102] = _0456_ ? _0503_ : _0502_;
  assign _0504_ = _0458_ & data_o[103];
  assign _0505_ = decrypt_i ? data_o[71] : sbox_data_i[7];
  assign _0506_ = _0505_ & next_ready_o;
  assign _0507_ = _0506_ | _0504_;
  assign _0508_ = _0170_ ? data_o[103] : sbox_data_i[7];
  assign next_data_reg[103] = _0456_ ? _0508_ : _0507_;
  assign _0509_ = _0458_ & data_o[104];
  assign _0510_ = next_ready_o & data_o[40];
  assign _0511_ = _0510_ | _0509_;
  assign _0512_ = _0473_ ? data_o[104] : sbox_data_i[0];
  assign next_data_reg[104] = _0456_ ? _0512_ : _0511_;
  assign _0513_ = _0458_ & data_o[105];
  assign _0514_ = next_ready_o & data_o[41];
  assign _0515_ = _0514_ | _0513_;
  assign _0516_ = _0473_ ? data_o[105] : sbox_data_i[1];
  assign next_data_reg[105] = _0456_ ? _0516_ : _0515_;
  assign _0517_ = _0458_ & data_o[106];
  assign _0518_ = next_ready_o & data_o[42];
  assign _0519_ = _0518_ | _0517_;
  assign _0520_ = _0473_ ? data_o[106] : sbox_data_i[2];
  assign next_data_reg[106] = _0456_ ? _0520_ : _0519_;
  assign _0521_ = _0458_ & data_o[107];
  assign _0522_ = next_ready_o & data_o[43];
  assign _0523_ = _0522_ | _0521_;
  assign _0524_ = _0473_ ? data_o[107] : sbox_data_i[3];
  assign next_data_reg[107] = _0456_ ? _0524_ : _0523_;
  assign _0525_ = _0458_ & data_o[108];
  assign _0526_ = next_ready_o & data_o[44];
  assign _0527_ = _0526_ | _0525_;
  assign _0528_ = _0473_ ? data_o[108] : sbox_data_i[4];
  assign next_data_reg[108] = _0456_ ? _0528_ : _0527_;
  assign _0529_ = _0458_ & data_o[109];
  assign _0530_ = next_ready_o & data_o[45];
  assign _0531_ = _0530_ | _0529_;
  assign _0532_ = _0473_ ? data_o[109] : sbox_data_i[5];
  assign next_data_reg[109] = _0456_ ? _0532_ : _0531_;
  assign _0533_ = _0458_ & data_o[10];
  assign _0534_ = next_ready_o & data_o[74];
  assign _0535_ = _0534_ | _0533_;
  assign _0536_ = _0477_ ? data_o[10] : sbox_data_i[2];
  assign next_data_reg[10] = _0456_ ? _0536_ : _0535_;
  assign _0537_ = _0458_ & data_o[110];
  assign _0538_ = next_ready_o & data_o[46];
  assign _0539_ = _0538_ | _0537_;
  assign _0540_ = _0473_ ? data_o[110] : sbox_data_i[6];
  assign next_data_reg[110] = _0456_ ? _0540_ : _0539_;
  assign _0541_ = _0458_ & data_o[111];
  assign _0542_ = next_ready_o & data_o[47];
  assign _0543_ = _0542_ | _0541_;
  assign _0544_ = _0473_ ? data_o[111] : sbox_data_i[7];
  assign next_data_reg[111] = _0456_ ? _0544_ : _0543_;
  assign _0545_ = _0458_ & data_o[112];
  assign _0546_ = decrypt_i ? data_o[16] : data_o[80];
  assign _0547_ = _0546_ & next_ready_o;
  assign _0548_ = _0547_ | _0545_;
  assign _0549_ = _0470_ ? data_o[112] : sbox_data_i[0];
  assign next_data_reg[112] = _0456_ ? _0549_ : _0548_;
  assign _0550_ = _0458_ & data_o[113];
  assign _0551_ = decrypt_i ? data_o[17] : data_o[81];
  assign _0552_ = _0551_ & next_ready_o;
  assign _0553_ = _0552_ | _0550_;
  assign _0554_ = _0470_ ? data_o[113] : sbox_data_i[1];
  assign next_data_reg[113] = _0456_ ? _0554_ : _0553_;
  assign _0555_ = _0458_ & data_o[114];
  assign _0556_ = decrypt_i ? data_o[18] : data_o[82];
  assign _0557_ = _0556_ & next_ready_o;
  assign _0558_ = _0557_ | _0555_;
  assign _0559_ = _0470_ ? data_o[114] : sbox_data_i[2];
  assign next_data_reg[114] = _0456_ ? _0559_ : _0558_;
  assign _0560_ = _0458_ & data_o[115];
  assign _0561_ = decrypt_i ? data_o[19] : data_o[83];
  assign _0562_ = _0561_ & next_ready_o;
  assign _0563_ = _0562_ | _0560_;
  assign _0564_ = _0470_ ? data_o[115] : sbox_data_i[3];
  assign next_data_reg[115] = _0456_ ? _0564_ : _0563_;
  assign _0565_ = _0458_ & data_o[116];
  assign _0566_ = decrypt_i ? data_o[20] : data_o[84];
  assign _0567_ = _0566_ & next_ready_o;
  assign _0568_ = _0567_ | _0565_;
  assign _0569_ = _0470_ ? data_o[116] : sbox_data_i[4];
  assign next_data_reg[116] = _0456_ ? _0569_ : _0568_;
  assign _0570_ = _0458_ & data_o[117];
  assign _0571_ = decrypt_i ? data_o[21] : data_o[85];
  assign _0572_ = _0571_ & next_ready_o;
  assign _0573_ = _0572_ | _0570_;
  assign _0574_ = _0470_ ? data_o[117] : sbox_data_i[5];
  assign next_data_reg[117] = _0456_ ? _0574_ : _0573_;
  assign _0575_ = _0458_ & data_o[118];
  assign _0576_ = decrypt_i ? data_o[22] : data_o[86];
  assign _0577_ = _0576_ & next_ready_o;
  assign _0578_ = _0577_ | _0575_;
  assign _0579_ = _0470_ ? data_o[118] : sbox_data_i[6];
  assign next_data_reg[118] = _0456_ ? _0579_ : _0578_;
  assign _0580_ = _0458_ & data_o[119];
  assign _0581_ = decrypt_i ? data_o[23] : data_o[87];
  assign _0582_ = _0581_ & next_ready_o;
  assign _0583_ = _0582_ | _0580_;
  assign _0584_ = _0470_ ? data_o[119] : sbox_data_i[7];
  assign next_data_reg[119] = _0456_ ? _0584_ : _0583_;
  assign _0585_ = _0458_ & data_o[11];
  assign _0586_ = next_ready_o & data_o[75];
  assign _0587_ = _0586_ | _0585_;
  assign _0588_ = _0477_ ? data_o[11] : sbox_data_i[3];
  assign next_data_reg[11] = _0456_ ? _0588_ : _0587_;
  assign _0589_ = _0458_ & data_o[120];
  assign _0590_ = next_ready_o & data_o[120];
  assign _0591_ = _0590_ | _0589_;
  assign _0592_ = _0467_ ? data_o[120] : sbox_data_i[0];
  assign next_data_reg[120] = _0456_ ? _0592_ : _0591_;
  assign _0593_ = _0458_ & data_o[121];
  assign _0594_ = next_ready_o & data_o[121];
  assign _0595_ = _0594_ | _0593_;
  assign _0596_ = _0467_ ? data_o[121] : sbox_data_i[1];
  assign next_data_reg[121] = _0456_ ? _0596_ : _0595_;
  assign _0597_ = _0458_ & data_o[122];
  assign _0598_ = next_ready_o & data_o[122];
  assign _0599_ = _0598_ | _0597_;
  assign _0600_ = _0467_ ? data_o[122] : sbox_data_i[2];
  assign next_data_reg[122] = _0456_ ? _0600_ : _0599_;
  assign _0601_ = _0458_ & data_o[123];
  assign _0602_ = next_ready_o & data_o[123];
  assign _0603_ = _0602_ | _0601_;
  assign _0604_ = _0467_ ? data_o[123] : sbox_data_i[3];
  assign next_data_reg[123] = _0456_ ? _0604_ : _0603_;
  assign _0605_ = _0458_ & data_o[124];
  assign _0606_ = next_ready_o & data_o[124];
  assign _0607_ = _0606_ | _0605_;
  assign _0608_ = _0467_ ? data_o[124] : sbox_data_i[4];
  assign next_data_reg[124] = _0456_ ? _0608_ : _0607_;
  assign _0609_ = _0458_ & data_o[125];
  assign _0610_ = next_ready_o & data_o[125];
  assign _0611_ = _0610_ | _0609_;
  assign _0612_ = _0467_ ? data_o[125] : sbox_data_i[5];
  assign next_data_reg[125] = _0456_ ? _0612_ : _0611_;
  assign _0613_ = _0458_ & data_o[126];
  assign _0614_ = next_ready_o & data_o[126];
  assign _0615_ = _0614_ | _0613_;
  assign _0616_ = _0467_ ? data_o[126] : sbox_data_i[6];
  assign next_data_reg[126] = _0456_ ? _0616_ : _0615_;
  assign _0617_ = _0458_ & data_o[127];
  assign _0618_ = next_ready_o & data_o[127];
  assign _0619_ = _0618_ | _0617_;
  assign _0620_ = _0467_ ? data_o[127] : sbox_data_i[7];
  assign next_data_reg[127] = _0456_ ? _0620_ : _0619_;
  assign _0621_ = _0458_ & data_o[12];
  assign _0622_ = next_ready_o & data_o[76];
  assign _0623_ = _0622_ | _0621_;
  assign _0624_ = _0477_ ? data_o[12] : sbox_data_i[4];
  assign next_data_reg[12] = _0456_ ? _0624_ : _0623_;
  assign _0625_ = _0458_ & data_o[13];
  assign _0626_ = next_ready_o & data_o[77];
  assign _0627_ = _0626_ | _0625_;
  assign _0628_ = _0477_ ? data_o[13] : sbox_data_i[5];
  assign next_data_reg[13] = _0456_ ? _0628_ : _0627_;
  assign _0629_ = _0458_ & data_o[14];
  assign _0630_ = next_ready_o & data_o[78];
  assign _0631_ = _0630_ | _0629_;
  assign _0632_ = _0477_ ? data_o[14] : sbox_data_i[6];
  assign next_data_reg[14] = _0456_ ? _0632_ : _0631_;
  assign _0633_ = _0458_ & data_o[15];
  assign _0634_ = next_ready_o & data_o[79];
  assign _0635_ = _0634_ | _0633_;
  assign _0636_ = _0477_ ? data_o[15] : sbox_data_i[7];
  assign next_data_reg[15] = _0456_ ? _0636_ : _0635_;
  assign _0637_ = _0458_ & data_o[16];
  assign _0638_ = decrypt_i ? data_o[48] : data_o[112];
  assign _0639_ = _0638_ & next_ready_o;
  assign _0640_ = _0639_ | _0637_;
  assign _0641_ = _0479_ ? data_o[16] : sbox_data_i[0];
  assign next_data_reg[16] = _0456_ ? _0641_ : _0640_;
  assign _0642_ = _0458_ & data_o[17];
  assign _0643_ = decrypt_i ? data_o[49] : data_o[113];
  assign _0644_ = _0643_ & next_ready_o;
  assign _0645_ = _0644_ | _0642_;
  assign _0646_ = _0479_ ? data_o[17] : sbox_data_i[1];
  assign next_data_reg[17] = _0456_ ? _0646_ : _0645_;
  assign _0647_ = _0458_ & data_o[18];
  assign _0648_ = decrypt_i ? data_o[50] : data_o[114];
  assign _0649_ = _0648_ & next_ready_o;
  assign _0650_ = _0649_ | _0647_;
  assign _0651_ = _0479_ ? data_o[18] : sbox_data_i[2];
  assign next_data_reg[18] = _0456_ ? _0651_ : _0650_;
  assign _0652_ = _0458_ & data_o[19];
  assign _0653_ = decrypt_i ? data_o[51] : data_o[115];
  assign _0654_ = _0653_ & next_ready_o;
  assign _0655_ = _0654_ | _0652_;
  assign _0656_ = _0479_ ? data_o[19] : sbox_data_i[3];
  assign next_data_reg[19] = _0456_ ? _0656_ : _0655_;
  assign _0657_ = _0458_ & data_o[1];
  assign _0658_ = decrypt_i ? data_o[97] : data_o[33];
  assign _0659_ = _0658_ & next_ready_o;
  assign _0660_ = _0659_ | _0657_;
  assign _0661_ = _0453_ ? sbox_data_i[1] : data_o[1];
  assign next_data_reg[1] = _0453_ ? _0660_ : _0661_;
  assign _0662_ = _0458_ & data_o[20];
  assign _0663_ = decrypt_i ? data_o[52] : data_o[116];
  assign _0664_ = _0663_ & next_ready_o;
  assign _0665_ = _0664_ | _0662_;
  assign _0666_ = _0479_ ? data_o[20] : sbox_data_i[4];
  assign next_data_reg[20] = _0456_ ? _0666_ : _0665_;
  assign _0667_ = _0458_ & data_o[21];
  assign _0668_ = decrypt_i ? data_o[53] : data_o[117];
  assign _0669_ = _0668_ & next_ready_o;
  assign _0670_ = _0669_ | _0667_;
  assign _0671_ = _0479_ ? data_o[21] : sbox_data_i[5];
  assign next_data_reg[21] = _0456_ ? _0671_ : _0670_;
  assign _0672_ = _0458_ & data_o[22];
  assign _0673_ = decrypt_i ? data_o[54] : data_o[118];
  assign _0674_ = _0673_ & next_ready_o;
  assign _0675_ = _0674_ | _0672_;
  assign _0676_ = _0479_ ? data_o[22] : sbox_data_i[6];
  assign next_data_reg[22] = _0456_ ? _0676_ : _0675_;
  assign _0677_ = _0458_ & data_o[23];
  assign _0678_ = decrypt_i ? data_o[55] : data_o[119];
  assign _0679_ = _0678_ & next_ready_o;
  assign _0680_ = _0679_ | _0677_;
  assign _0681_ = _0479_ ? data_o[23] : sbox_data_i[7];
  assign next_data_reg[23] = _0456_ ? _0681_ : _0680_;
  assign _0682_ = _0458_ & data_o[24];
  assign _0683_ = next_ready_o & data_o[24];
  assign _0684_ = _0683_ | _0682_;
  assign _0685_ = _0481_ ? data_o[24] : sbox_data_i[0];
  assign next_data_reg[24] = _0456_ ? _0685_ : _0684_;
  assign _0686_ = _0458_ & data_o[25];
  assign _0687_ = next_ready_o & data_o[25];
  assign _0688_ = _0687_ | _0686_;
  assign _0689_ = _0481_ ? data_o[25] : sbox_data_i[1];
  assign next_data_reg[25] = _0456_ ? _0689_ : _0688_;
  assign _0690_ = _0458_ & data_o[26];
  assign _0691_ = next_ready_o & data_o[26];
  assign _0692_ = _0691_ | _0690_;
  assign _0693_ = _0481_ ? data_o[26] : sbox_data_i[2];
  assign next_data_reg[26] = _0456_ ? _0693_ : _0692_;
  assign _0694_ = _0458_ & data_o[27];
  assign _0695_ = next_ready_o & data_o[27];
  assign _0696_ = _0695_ | _0694_;
  assign _0697_ = _0481_ ? data_o[27] : sbox_data_i[3];
  assign next_data_reg[27] = _0456_ ? _0697_ : _0696_;
  assign _0698_ = _0458_ & data_o[28];
  assign _0699_ = next_ready_o & data_o[28];
  assign _0700_ = _0699_ | _0698_;
  assign _0701_ = _0481_ ? data_o[28] : sbox_data_i[4];
  assign next_data_reg[28] = _0456_ ? _0701_ : _0700_;
  assign _0702_ = _0458_ & data_o[29];
  assign _0703_ = next_ready_o & data_o[29];
  assign _0704_ = _0703_ | _0702_;
  assign _0705_ = _0481_ ? data_o[29] : sbox_data_i[5];
  assign next_data_reg[29] = _0456_ ? _0705_ : _0704_;
  assign _0706_ = _0458_ & data_o[2];
  assign _0707_ = decrypt_i ? data_o[98] : data_o[34];
  assign _0708_ = _0707_ & next_ready_o;
  assign _0709_ = _0708_ | _0706_;
  assign _0710_ = _0453_ ? sbox_data_i[2] : data_o[2];
  assign next_data_reg[2] = _0453_ ? _0709_ : _0710_;
  assign _0711_ = _0458_ & data_o[30];
  assign _0712_ = next_ready_o & data_o[30];
  assign _0713_ = _0712_ | _0711_;
  assign _0714_ = _0481_ ? data_o[30] : sbox_data_i[6];
  assign next_data_reg[30] = _0456_ ? _0714_ : _0713_;
  assign _0715_ = _0458_ & data_o[31];
  assign _0716_ = next_ready_o & data_o[31];
  assign _0717_ = _0716_ | _0715_;
  assign _0718_ = _0481_ ? data_o[31] : sbox_data_i[7];
  assign next_data_reg[31] = _0456_ ? _0718_ : _0717_;
  assign _0719_ = _0458_ & data_o[32];
  assign _0720_ = decrypt_i ? sbox_data_i[0] : data_o[64];
  assign _0721_ = _0720_ & next_ready_o;
  assign _0722_ = _0721_ | _0719_;
  assign _0723_ = _0175_ ? data_o[32] : sbox_data_i[0];
  assign next_data_reg[32] = _0456_ ? _0723_ : _0722_;
  assign _0724_ = _0458_ & data_o[33];
  assign _0725_ = decrypt_i ? sbox_data_i[1] : data_o[65];
  assign _0726_ = _0725_ & next_ready_o;
  assign _0727_ = _0726_ | _0724_;
  assign _0728_ = _0175_ ? data_o[33] : sbox_data_i[1];
  assign next_data_reg[33] = _0456_ ? _0728_ : _0727_;
  assign _0729_ = _0458_ & data_o[34];
  assign _0730_ = decrypt_i ? sbox_data_i[2] : data_o[66];
  assign _0731_ = _0730_ & next_ready_o;
  assign _0732_ = _0731_ | _0729_;
  assign _0733_ = _0175_ ? data_o[34] : sbox_data_i[2];
  assign next_data_reg[34] = _0456_ ? _0733_ : _0732_;
  assign _0734_ = _0458_ & data_o[35];
  assign _0735_ = decrypt_i ? sbox_data_i[3] : data_o[67];
  assign _0736_ = _0735_ & next_ready_o;
  assign _0737_ = _0736_ | _0734_;
  assign _0738_ = _0175_ ? data_o[35] : sbox_data_i[3];
  assign next_data_reg[35] = _0456_ ? _0738_ : _0737_;
  assign _0739_ = _0458_ & data_o[36];
  assign _0740_ = decrypt_i ? sbox_data_i[4] : data_o[68];
  assign _0741_ = _0740_ & next_ready_o;
  assign _0742_ = _0741_ | _0739_;
  assign _0743_ = _0175_ ? data_o[36] : sbox_data_i[4];
  assign next_data_reg[36] = _0456_ ? _0743_ : _0742_;
  assign _0744_ = _0458_ & data_o[37];
  assign _0745_ = decrypt_i ? sbox_data_i[5] : data_o[69];
  assign _0746_ = _0745_ & next_ready_o;
  assign _0747_ = _0746_ | _0744_;
  assign _0748_ = _0175_ ? data_o[37] : sbox_data_i[5];
  assign next_data_reg[37] = _0456_ ? _0748_ : _0747_;
  assign _0749_ = _0458_ & data_o[38];
  assign _0750_ = decrypt_i ? sbox_data_i[6] : data_o[70];
  assign _0751_ = _0750_ & next_ready_o;
  assign _0752_ = _0751_ | _0749_;
  assign _0753_ = _0175_ ? data_o[38] : sbox_data_i[6];
  assign next_data_reg[38] = _0456_ ? _0753_ : _0752_;
  assign _0754_ = _0458_ & data_o[39];
  assign _0755_ = decrypt_i ? sbox_data_i[7] : data_o[71];
  assign _0756_ = _0755_ & next_ready_o;
  assign _0757_ = _0756_ | _0754_;
  assign _0758_ = _0175_ ? data_o[39] : sbox_data_i[7];
  assign next_data_reg[39] = _0456_ ? _0758_ : _0757_;
  assign _0759_ = _0458_ & data_o[3];
  assign _0760_ = decrypt_i ? data_o[99] : data_o[35];
  assign _0761_ = _0760_ & next_ready_o;
  assign _0762_ = _0761_ | _0759_;
  assign _0763_ = _0453_ ? sbox_data_i[3] : data_o[3];
  assign next_data_reg[3] = _0453_ ? _0762_ : _0763_;
  assign _0764_ = _0458_ & data_o[40];
  assign _0765_ = next_ready_o & data_o[104];
  assign _0766_ = _0765_ | _0764_;
  assign _0767_ = _0482_ ? data_o[40] : sbox_data_i[0];
  assign next_data_reg[40] = _0456_ ? _0767_ : _0766_;
  assign _0768_ = _0458_ & data_o[41];
  assign _0769_ = next_ready_o & data_o[105];
  assign _0770_ = _0769_ | _0768_;
  assign _0771_ = _0482_ ? data_o[41] : sbox_data_i[1];
  assign next_data_reg[41] = _0456_ ? _0771_ : _0770_;
  assign _0772_ = _0458_ & data_o[42];
  assign _0773_ = next_ready_o & data_o[106];
  assign _0774_ = _0773_ | _0772_;
  assign _0775_ = _0482_ ? data_o[42] : sbox_data_i[2];
  assign next_data_reg[42] = _0456_ ? _0775_ : _0774_;
  assign _0776_ = _0458_ & data_o[43];
  assign _0777_ = next_ready_o & data_o[107];
  assign _0778_ = _0777_ | _0776_;
  assign _0779_ = _0482_ ? data_o[43] : sbox_data_i[3];
  assign next_data_reg[43] = _0456_ ? _0779_ : _0778_;
  assign _0780_ = _0458_ & data_o[44];
  assign _0781_ = next_ready_o & data_o[108];
  assign _0782_ = _0781_ | _0780_;
  assign _0783_ = _0482_ ? data_o[44] : sbox_data_i[4];
  assign next_data_reg[44] = _0456_ ? _0783_ : _0782_;
  assign _0784_ = _0458_ & data_o[45];
  assign _0785_ = next_ready_o & data_o[109];
  assign _0786_ = _0785_ | _0784_;
  assign _0787_ = _0482_ ? data_o[45] : sbox_data_i[5];
  assign next_data_reg[45] = _0456_ ? _0787_ : _0786_;
  assign _0788_ = _0458_ & data_o[46];
  assign _0789_ = next_ready_o & data_o[110];
  assign _0790_ = _0789_ | _0788_;
  assign _0791_ = _0482_ ? data_o[46] : sbox_data_i[6];
  assign next_data_reg[46] = _0456_ ? _0791_ : _0790_;
  assign _0792_ = _0458_ & data_o[47];
  assign _0793_ = next_ready_o & data_o[111];
  assign _0794_ = _0793_ | _0792_;
  assign _0795_ = _0482_ ? data_o[47] : sbox_data_i[7];
  assign next_data_reg[47] = _0456_ ? _0795_ : _0794_;
  assign _0796_ = _0458_ & data_o[48];
  assign _0797_ = decrypt_i ? data_o[80] : data_o[16];
  assign _0798_ = _0797_ & next_ready_o;
  assign _0799_ = _0798_ | _0796_;
  assign _0800_ = _0484_ ? data_o[48] : sbox_data_i[0];
  assign next_data_reg[48] = _0456_ ? _0800_ : _0799_;
  assign _0801_ = _0458_ & data_o[49];
  assign _0802_ = decrypt_i ? data_o[81] : data_o[17];
  assign _0803_ = _0802_ & next_ready_o;
  assign _0804_ = _0803_ | _0801_;
  assign _0805_ = _0484_ ? data_o[49] : sbox_data_i[1];
  assign next_data_reg[49] = _0456_ ? _0805_ : _0804_;
  assign _0806_ = _0458_ & data_o[4];
  assign _0807_ = decrypt_i ? data_o[100] : data_o[36];
  assign _0808_ = _0807_ & next_ready_o;
  assign _0809_ = _0808_ | _0806_;
  assign _0810_ = _0453_ ? sbox_data_i[4] : data_o[4];
  assign next_data_reg[4] = _0453_ ? _0809_ : _0810_;
  assign _0811_ = _0458_ & data_o[50];
  assign _0812_ = decrypt_i ? data_o[82] : data_o[18];
  assign _0813_ = _0812_ & next_ready_o;
  assign _0814_ = _0813_ | _0811_;
  assign _0815_ = _0484_ ? data_o[50] : sbox_data_i[2];
  assign next_data_reg[50] = _0456_ ? _0815_ : _0814_;
  assign _0816_ = _0458_ & data_o[51];
  assign _0817_ = decrypt_i ? data_o[83] : data_o[19];
  assign _0818_ = _0817_ & next_ready_o;
  assign _0819_ = _0818_ | _0816_;
  assign _0820_ = _0484_ ? data_o[51] : sbox_data_i[3];
  assign next_data_reg[51] = _0456_ ? _0820_ : _0819_;
  assign _0821_ = _0458_ & data_o[52];
  assign _0822_ = decrypt_i ? data_o[84] : data_o[20];
  assign _0823_ = _0822_ & next_ready_o;
  assign _0824_ = _0823_ | _0821_;
  assign _0825_ = _0484_ ? data_o[52] : sbox_data_i[4];
  assign next_data_reg[52] = _0456_ ? _0825_ : _0824_;
  assign _0826_ = _0458_ & data_o[53];
  assign _0827_ = decrypt_i ? data_o[85] : data_o[21];
  assign _0828_ = _0827_ & next_ready_o;
  assign _0829_ = _0828_ | _0826_;
  assign _0830_ = _0484_ ? data_o[53] : sbox_data_i[5];
  assign next_data_reg[53] = _0456_ ? _0830_ : _0829_;
  assign _0831_ = _0458_ & data_o[54];
  assign _0832_ = decrypt_i ? data_o[86] : data_o[22];
  assign _0833_ = _0832_ & next_ready_o;
  assign _0834_ = _0833_ | _0831_;
  assign _0835_ = _0484_ ? data_o[54] : sbox_data_i[6];
  assign next_data_reg[54] = _0456_ ? _0835_ : _0834_;
  assign _0836_ = _0458_ & data_o[55];
  assign _0837_ = decrypt_i ? data_o[87] : data_o[23];
  assign _0838_ = _0837_ & next_ready_o;
  assign _0839_ = _0838_ | _0836_;
  assign _0840_ = _0484_ ? data_o[55] : sbox_data_i[7];
  assign next_data_reg[55] = _0456_ ? _0840_ : _0839_;
  assign _0841_ = _0458_ & data_o[56];
  assign _0842_ = next_ready_o & data_o[56];
  assign _0843_ = _0842_ | _0841_;
  assign _0844_ = _0483_ ? data_o[56] : sbox_data_i[0];
  assign next_data_reg[56] = _0456_ ? _0844_ : _0843_;
  assign _0845_ = _0458_ & data_o[57];
  assign _0846_ = next_ready_o & data_o[57];
  assign _0847_ = _0846_ | _0845_;
  assign _0848_ = _0483_ ? data_o[57] : sbox_data_i[1];
  assign next_data_reg[57] = _0456_ ? _0848_ : _0847_;
  assign _0849_ = _0458_ & data_o[58];
  assign _0850_ = next_ready_o & data_o[58];
  assign _0851_ = _0850_ | _0849_;
  assign _0852_ = _0483_ ? data_o[58] : sbox_data_i[2];
  assign next_data_reg[58] = _0456_ ? _0852_ : _0851_;
  assign _0853_ = _0458_ & data_o[59];
  assign _0854_ = next_ready_o & data_o[59];
  assign _0855_ = _0854_ | _0853_;
  assign _0856_ = _0483_ ? data_o[59] : sbox_data_i[3];
  assign next_data_reg[59] = _0456_ ? _0856_ : _0855_;
  assign _0857_ = _0458_ & data_o[5];
  assign _0858_ = decrypt_i ? data_o[101] : data_o[37];
  assign _0859_ = _0858_ & next_ready_o;
  assign _0860_ = _0859_ | _0857_;
  assign _0861_ = _0453_ ? sbox_data_i[5] : data_o[5];
  assign next_data_reg[5] = _0453_ ? _0860_ : _0861_;
  assign _0862_ = _0458_ & data_o[60];
  assign _0863_ = next_ready_o & data_o[60];
  assign _0864_ = _0863_ | _0862_;
  assign _0865_ = _0483_ ? data_o[60] : sbox_data_i[4];
  assign next_data_reg[60] = _0456_ ? _0865_ : _0864_;
  assign _0866_ = _0458_ & data_o[61];
  assign _0867_ = next_ready_o & data_o[61];
  assign _0868_ = _0867_ | _0866_;
  assign _0869_ = _0483_ ? data_o[61] : sbox_data_i[5];
  assign next_data_reg[61] = _0456_ ? _0869_ : _0868_;
  assign _0870_ = _0458_ & data_o[62];
  assign _0871_ = next_ready_o & data_o[62];
  assign _0872_ = _0871_ | _0870_;
  assign _0873_ = _0483_ ? data_o[62] : sbox_data_i[6];
  assign next_data_reg[62] = _0456_ ? _0873_ : _0872_;
  assign _0874_ = _0458_ & data_o[63];
  assign _0875_ = next_ready_o & data_o[63];
  assign _0876_ = _0875_ | _0874_;
  assign _0877_ = _0483_ ? data_o[63] : sbox_data_i[7];
  assign next_data_reg[63] = _0456_ ? _0877_ : _0876_;
  assign _0878_ = _0458_ & data_o[64];
  assign _0879_ = decrypt_i ? data_o[32] : data_o[96];
  assign _0880_ = _0879_ & next_ready_o;
  assign _0881_ = _0880_ | _0878_;
  assign _0882_ = _0176_ ? data_o[64] : sbox_data_i[0];
  assign next_data_reg[64] = _0456_ ? _0882_ : _0881_;
  assign _0883_ = _0458_ & data_o[65];
  assign _0884_ = decrypt_i ? data_o[33] : data_o[97];
  assign _0885_ = _0884_ & next_ready_o;
  assign _0886_ = _0885_ | _0883_;
  assign _0887_ = _0176_ ? data_o[65] : sbox_data_i[1];
  assign next_data_reg[65] = _0456_ ? _0887_ : _0886_;
  assign _0888_ = _0458_ & data_o[66];
  assign _0889_ = decrypt_i ? data_o[34] : data_o[98];
  assign _0890_ = _0889_ & next_ready_o;
  assign _0891_ = _0890_ | _0888_;
  assign _0892_ = _0176_ ? data_o[66] : sbox_data_i[2];
  assign next_data_reg[66] = _0456_ ? _0892_ : _0891_;
  assign _0893_ = _0458_ & data_o[67];
  assign _0894_ = decrypt_i ? data_o[35] : data_o[99];
  assign _0895_ = _0894_ & next_ready_o;
  assign _0896_ = _0895_ | _0893_;
  assign _0897_ = _0176_ ? data_o[67] : sbox_data_i[3];
  assign next_data_reg[67] = _0456_ ? _0897_ : _0896_;
  assign _0898_ = _0458_ & data_o[68];
  assign _0899_ = decrypt_i ? data_o[36] : data_o[100];
  assign _0900_ = _0899_ & next_ready_o;
  assign _0901_ = _0900_ | _0898_;
  assign _0902_ = _0176_ ? data_o[68] : sbox_data_i[4];
  assign next_data_reg[68] = _0456_ ? _0902_ : _0901_;
  assign _0903_ = _0458_ & data_o[69];
  assign _0904_ = decrypt_i ? data_o[37] : data_o[101];
  assign _0905_ = _0904_ & next_ready_o;
  assign _0906_ = _0905_ | _0903_;
  assign _0907_ = _0176_ ? data_o[69] : sbox_data_i[5];
  assign next_data_reg[69] = _0456_ ? _0907_ : _0906_;
  assign _0908_ = _0458_ & data_o[6];
  assign _0909_ = decrypt_i ? data_o[102] : data_o[38];
  assign _0910_ = _0909_ & next_ready_o;
  assign _0911_ = _0910_ | _0908_;
  assign _0912_ = _0453_ ? sbox_data_i[6] : data_o[6];
  assign next_data_reg[6] = _0453_ ? _0911_ : _0912_;
  assign _0000_ = _0458_ & data_o[70];
  assign _0001_ = decrypt_i ? data_o[38] : data_o[102];
  assign _0002_ = _0001_ & next_ready_o;
  assign _0003_ = _0002_ | _0000_;
  assign _0004_ = _0176_ ? data_o[70] : sbox_data_i[6];
  assign next_data_reg[70] = _0456_ ? _0004_ : _0003_;
  assign _0005_ = _0458_ & data_o[71];
  assign _0006_ = decrypt_i ? data_o[39] : data_o[103];
  assign _0007_ = _0006_ & next_ready_o;
  assign _0008_ = _0007_ | _0005_;
  assign _0009_ = _0176_ ? data_o[71] : sbox_data_i[7];
  assign next_data_reg[71] = _0456_ ? _0009_ : _0008_;
  assign _0010_ = _0458_ & data_o[72];
  assign _0011_ = next_ready_o & data_o[8];
  assign _0012_ = _0011_ | _0010_;
  assign _0013_ = _0487_ ? data_o[72] : sbox_data_i[0];
  assign next_data_reg[72] = _0456_ ? _0013_ : _0012_;
  assign _0014_ = _0458_ & data_o[73];
  assign _0015_ = next_ready_o & data_o[9];
  assign _0016_ = _0015_ | _0014_;
  assign _0017_ = _0487_ ? data_o[73] : sbox_data_i[1];
  assign next_data_reg[73] = _0456_ ? _0017_ : _0016_;
  assign _0018_ = _0458_ & data_o[74];
  assign _0019_ = next_ready_o & data_o[10];
  assign _0020_ = _0019_ | _0018_;
  assign _0021_ = _0487_ ? data_o[74] : sbox_data_i[2];
  assign next_data_reg[74] = _0456_ ? _0021_ : _0020_;
  assign _0022_ = _0458_ & data_o[75];
  assign _0023_ = next_ready_o & data_o[11];
  assign _0024_ = _0023_ | _0022_;
  assign _0025_ = _0487_ ? data_o[75] : sbox_data_i[3];
  assign next_data_reg[75] = _0456_ ? _0025_ : _0024_;
  assign _0026_ = _0458_ & data_o[76];
  assign _0027_ = next_ready_o & data_o[12];
  assign _0028_ = _0027_ | _0026_;
  assign _0029_ = _0487_ ? data_o[76] : sbox_data_i[4];
  assign next_data_reg[76] = _0456_ ? _0029_ : _0028_;
  assign _0030_ = _0458_ & data_o[77];
  assign _0031_ = next_ready_o & data_o[13];
  assign _0032_ = _0031_ | _0030_;
  assign _0033_ = _0487_ ? data_o[77] : sbox_data_i[5];
  assign next_data_reg[77] = _0456_ ? _0033_ : _0032_;
  assign _0034_ = _0458_ & data_o[78];
  assign _0035_ = next_ready_o & data_o[14];
  assign _0036_ = _0035_ | _0034_;
  assign _0037_ = _0487_ ? data_o[78] : sbox_data_i[6];
  assign next_data_reg[78] = _0456_ ? _0037_ : _0036_;
  assign _0038_ = _0458_ & data_o[79];
  assign _0039_ = next_ready_o & data_o[15];
  assign _0040_ = _0039_ | _0038_;
  assign _0041_ = _0487_ ? data_o[79] : sbox_data_i[7];
  assign next_data_reg[79] = _0456_ ? _0041_ : _0040_;
  assign _0042_ = _0458_ & data_o[7];
  assign _0043_ = decrypt_i ? data_o[103] : data_o[39];
  assign _0044_ = _0043_ & next_ready_o;
  assign _0045_ = _0044_ | _0042_;
  assign _0046_ = _0453_ ? sbox_data_i[7] : data_o[7];
  assign next_data_reg[7] = _0453_ ? _0045_ : _0046_;
  assign _0047_ = _0458_ & data_o[80];
  assign _0048_ = decrypt_i ? data_o[112] : data_o[48];
  assign _0049_ = _0048_ & next_ready_o;
  assign _0050_ = _0049_ | _0047_;
  assign _0051_ = _0486_ ? data_o[80] : sbox_data_i[0];
  assign next_data_reg[80] = _0456_ ? _0051_ : _0050_;
  assign _0052_ = _0458_ & data_o[81];
  assign _0053_ = decrypt_i ? data_o[113] : data_o[49];
  assign _0054_ = _0053_ & next_ready_o;
  assign _0055_ = _0054_ | _0052_;
  assign _0056_ = _0486_ ? data_o[81] : sbox_data_i[1];
  assign next_data_reg[81] = _0456_ ? _0056_ : _0055_;
  assign _0057_ = _0458_ & data_o[82];
  assign _0058_ = decrypt_i ? data_o[114] : data_o[50];
  assign _0059_ = _0058_ & next_ready_o;
  assign _0060_ = _0059_ | _0057_;
  assign _0061_ = _0486_ ? data_o[82] : sbox_data_i[2];
  assign next_data_reg[82] = _0456_ ? _0061_ : _0060_;
  assign _0062_ = _0458_ & data_o[83];
  assign _0063_ = decrypt_i ? data_o[115] : data_o[51];
  assign _0064_ = _0063_ & next_ready_o;
  assign _0065_ = _0064_ | _0062_;
  assign _0066_ = _0486_ ? data_o[83] : sbox_data_i[3];
  assign next_data_reg[83] = _0456_ ? _0066_ : _0065_;
  assign _0067_ = _0458_ & data_o[84];
  assign _0068_ = decrypt_i ? data_o[116] : data_o[52];
  assign _0069_ = _0068_ & next_ready_o;
  assign _0070_ = _0069_ | _0067_;
  assign _0071_ = _0486_ ? data_o[84] : sbox_data_i[4];
  assign next_data_reg[84] = _0456_ ? _0071_ : _0070_;
  assign _0072_ = _0458_ & data_o[85];
  assign _0073_ = decrypt_i ? data_o[117] : data_o[53];
  assign _0074_ = _0073_ & next_ready_o;
  assign _0075_ = _0074_ | _0072_;
  assign _0076_ = _0486_ ? data_o[85] : sbox_data_i[5];
  assign next_data_reg[85] = _0456_ ? _0076_ : _0075_;
  assign _0077_ = _0458_ & data_o[86];
  assign _0078_ = decrypt_i ? data_o[118] : data_o[54];
  assign _0079_ = _0078_ & next_ready_o;
  assign _0080_ = _0079_ | _0077_;
  assign _0081_ = _0486_ ? data_o[86] : sbox_data_i[6];
  assign next_data_reg[86] = _0456_ ? _0081_ : _0080_;
  assign _0082_ = _0458_ & data_o[87];
  assign _0083_ = decrypt_i ? data_o[119] : data_o[55];
  assign _0084_ = _0083_ & next_ready_o;
  assign _0085_ = _0084_ | _0082_;
  assign _0086_ = _0486_ ? data_o[87] : sbox_data_i[7];
  assign next_data_reg[87] = _0456_ ? _0086_ : _0085_;
  assign _0087_ = _0458_ & data_o[88];
  assign _0088_ = next_ready_o & data_o[88];
  assign _0089_ = _0088_ | _0087_;
  assign _0090_ = _0485_ ? data_o[88] : sbox_data_i[0];
  assign next_data_reg[88] = _0456_ ? _0090_ : _0089_;
  assign _0091_ = _0458_ & data_o[89];
  assign _0092_ = next_ready_o & data_o[89];
  assign _0093_ = _0092_ | _0091_;
  assign _0094_ = _0485_ ? data_o[89] : sbox_data_i[1];
  assign next_data_reg[89] = _0456_ ? _0094_ : _0093_;
  assign _0095_ = _0458_ & data_o[8];
  assign _0096_ = next_ready_o & data_o[72];
  assign _0097_ = _0096_ | _0095_;
  assign _0098_ = _0477_ ? data_o[8] : sbox_data_i[0];
  assign next_data_reg[8] = _0456_ ? _0098_ : _0097_;
  assign _0099_ = _0458_ & data_o[90];
  assign _0100_ = next_ready_o & data_o[90];
  assign _0101_ = _0100_ | _0099_;
  assign _0102_ = _0485_ ? data_o[90] : sbox_data_i[2];
  assign next_data_reg[90] = _0456_ ? _0102_ : _0101_;
  assign _0103_ = _0458_ & data_o[91];
  assign _0104_ = next_ready_o & data_o[91];
  assign _0105_ = _0104_ | _0103_;
  assign _0106_ = _0485_ ? data_o[91] : sbox_data_i[3];
  assign next_data_reg[91] = _0456_ ? _0106_ : _0105_;
  assign _0107_ = _0458_ & data_o[92];
  assign _0108_ = next_ready_o & data_o[92];
  assign _0109_ = _0108_ | _0107_;
  assign _0110_ = _0485_ ? data_o[92] : sbox_data_i[4];
  assign next_data_reg[92] = _0456_ ? _0110_ : _0109_;
  assign _0111_ = _0458_ & data_o[93];
  assign _0112_ = next_ready_o & data_o[93];
  assign _0113_ = _0112_ | _0111_;
  assign _0114_ = _0485_ ? data_o[93] : sbox_data_i[5];
  assign next_data_reg[93] = _0456_ ? _0114_ : _0113_;
  assign _0115_ = _0458_ & data_o[94];
  assign _0116_ = next_ready_o & data_o[94];
  assign _0117_ = _0116_ | _0115_;
  assign _0118_ = _0485_ ? data_o[94] : sbox_data_i[6];
  assign next_data_reg[94] = _0456_ ? _0118_ : _0117_;
  assign _0119_ = _0458_ & data_o[95];
  assign _0120_ = next_ready_o & data_o[95];
  assign _0121_ = _0120_ | _0119_;
  assign _0122_ = _0485_ ? data_o[95] : sbox_data_i[7];
  assign next_data_reg[95] = _0456_ ? _0122_ : _0121_;
  assign _0123_ = _0458_ & data_o[96];
  assign _0124_ = decrypt_i ? data_o[64] : sbox_data_i[0];
  assign _0125_ = _0124_ & next_ready_o;
  assign _0126_ = _0125_ | _0123_;
  assign _0127_ = _0170_ ? data_o[96] : sbox_data_i[0];
  assign next_data_reg[96] = _0456_ ? _0127_ : _0126_;
  assign _0128_ = _0458_ & data_o[97];
  assign _0129_ = decrypt_i ? data_o[65] : sbox_data_i[1];
  assign _0130_ = _0129_ & next_ready_o;
  assign _0131_ = _0130_ | _0128_;
  assign _0132_ = _0170_ ? data_o[97] : sbox_data_i[1];
  assign next_data_reg[97] = _0456_ ? _0132_ : _0131_;
  assign _0133_ = _0458_ & data_o[98];
  assign _0134_ = decrypt_i ? data_o[66] : sbox_data_i[2];
  assign _0135_ = _0134_ & next_ready_o;
  assign _0136_ = _0135_ | _0133_;
  assign _0137_ = _0170_ ? data_o[98] : sbox_data_i[2];
  assign next_data_reg[98] = _0456_ ? _0137_ : _0136_;
  assign _0138_ = _0458_ & data_o[99];
  assign _0139_ = decrypt_i ? data_o[67] : sbox_data_i[3];
  assign _0140_ = _0139_ & next_ready_o;
  assign _0141_ = _0140_ | _0138_;
  assign _0142_ = _0170_ ? data_o[99] : sbox_data_i[3];
  assign next_data_reg[99] = _0456_ ? _0142_ : _0141_;
  assign _0143_ = _0458_ & data_o[9];
  assign _0144_ = next_ready_o & data_o[73];
  assign _0145_ = _0144_ | _0143_;
  assign _0146_ = _0477_ ? data_o[9] : sbox_data_i[1];
  assign next_data_reg[9] = _0456_ ? _0146_ : _0145_;
  assign _0147_ = start_i | state[0];
  assign _0148_ = _0147_ & _0458_;
  assign next_state[0] = _0456_ ? _0449_ : _0148_;
  assign _0149_ = ~start_i;
  assign _0150_ = _0149_ & state[1];
  assign _0151_ = _0150_ & _0458_;
  assign _0152_ = state[1] ^ state[0];
  assign next_state[1] = _0456_ ? _0152_ : _0151_;
  assign _0153_ = _0149_ & state[2];
  assign _0154_ = _0153_ & _0458_;
  assign _0155_ = state[1] & state[0];
  assign _0156_ = _0155_ ^ state[2];
  assign next_state[2] = _0456_ ? _0156_ : _0154_;
  assign _0157_ = _0149_ & state[3];
  assign _0158_ = _0157_ & _0458_;
  assign _0159_ = _0155_ & state[2];
  assign _0160_ = _0159_ ^ state[3];
  assign next_state[3] = _0456_ ? _0160_ : _0158_;
  assign _0161_ = _0149_ & state[4];
  assign _0162_ = _0161_ & _0458_;
  assign _0163_ = _0159_ & state[3];
  assign _0164_ = _0163_ ^ state[4];
  assign next_state[4] = _0456_ ? _0164_ : _0162_;
  assign _0165_ = data_i[120] & start_i;
  assign _0166_ = _0165_ & _0458_;
  assign _0167_ = _0155_ & _0448_;
  assign _0168_ = _0167_ & _0447_;
  assign _0169_ = _0454_ | _0448_;
  assign _0170_ = _0169_ | state[3];
  assign _0171_ = _0159_ & _0447_;
  assign _0172_ = state[1] & _0449_;
  assign _0173_ = _0172_ & state[2];
  assign _0174_ = _0173_ & state[3];
  assign _0175_ = _0169_ | _0447_;
  assign _0176_ = _0455_ | _0447_;
  assign _0177_ = _0167_ & state[3];
  assign _0178_ = _0451_ & state[2];
  assign _0179_ = _0178_ & _0447_;
  assign _0180_ = _0179_ & data_i[88];
  assign _0181_ = _0450_ & state[0];
  assign _0182_ = _0181_ & state[2];
  assign _0183_ = _0182_ & _0447_;
  assign _0184_ = _0183_ & data_i[80];
  assign _0185_ = _0184_ | _0180_;
  assign _0186_ = _0173_ & _0447_;
  assign _0187_ = _0186_ & data_i[72];
  assign _0188_ = _0171_ & data_i[64];
  assign _0189_ = _0188_ | _0187_;
  assign _0190_ = _0189_ | _0185_;
  assign _0191_ = _0453_ & data_i[120];
  assign _0192_ = _0181_ & _0448_;
  assign _0193_ = _0192_ & _0447_;
  assign _0194_ = _0193_ & data_i[112];
  assign _0195_ = _0194_ | _0191_;
  assign _0196_ = _0172_ & _0448_;
  assign _0197_ = _0196_ & _0447_;
  assign _0198_ = _0197_ & data_i[104];
  assign _0199_ = _0168_ & data_i[96];
  assign _0200_ = _0199_ | _0198_;
  assign _0201_ = _0200_ | _0195_;
  assign _0202_ = _0201_ | _0190_;
  assign _0203_ = _0174_ & data_i[8];
  assign _0204_ = _0178_ & state[3];
  assign _0205_ = _0204_ & data_i[24];
  assign _0206_ = _0182_ & state[3];
  assign _0207_ = _0206_ & data_i[16];
  assign _0208_ = _0207_ | _0205_;
  assign _0209_ = _0208_ | _0203_;
  assign _0210_ = _0452_ & state[3];
  assign _0211_ = _0210_ & data_i[56];
  assign _0212_ = _0192_ & state[3];
  assign _0213_ = _0212_ & data_i[48];
  assign _0214_ = _0213_ | _0211_;
  assign _0215_ = _0196_ & state[3];
  assign _0216_ = _0215_ & data_i[40];
  assign _0217_ = _0177_ & data_i[32];
  assign _0218_ = _0217_ | _0216_;
  assign _0219_ = _0218_ | _0214_;
  assign _0220_ = _0219_ | _0209_;
  assign _0221_ = _0220_ | _0202_;
  assign _0222_ = _0163_ ? data_i[0] : _0221_;
  assign sbox_data_o[0] = _0453_ ? _0166_ : _0222_;
  assign _0223_ = data_i[121] & start_i;
  assign _0224_ = _0223_ & _0458_;
  assign _0225_ = _0179_ & data_i[89];
  assign _0226_ = _0183_ & data_i[81];
  assign _0227_ = _0226_ | _0225_;
  assign _0228_ = _0186_ & data_i[73];
  assign _0229_ = _0171_ & data_i[65];
  assign _0230_ = _0229_ | _0228_;
  assign _0231_ = _0230_ | _0227_;
  assign _0232_ = _0453_ & data_i[121];
  assign _0233_ = _0193_ & data_i[113];
  assign _0234_ = _0233_ | _0232_;
  assign _0235_ = _0197_ & data_i[105];
  assign _0236_ = _0168_ & data_i[97];
  assign _0237_ = _0236_ | _0235_;
  assign _0238_ = _0237_ | _0234_;
  assign _0239_ = _0238_ | _0231_;
  assign _0240_ = _0174_ & data_i[9];
  assign _0241_ = _0204_ & data_i[25];
  assign _0242_ = _0206_ & data_i[17];
  assign _0243_ = _0242_ | _0241_;
  assign _0244_ = _0243_ | _0240_;
  assign _0245_ = _0210_ & data_i[57];
  assign _0246_ = _0212_ & data_i[49];
  assign _0247_ = _0246_ | _0245_;
  assign _0248_ = _0215_ & data_i[41];
  assign _0249_ = _0177_ & data_i[33];
  assign _0250_ = _0249_ | _0248_;
  assign _0251_ = _0250_ | _0247_;
  assign _0252_ = _0251_ | _0244_;
  assign _0253_ = _0252_ | _0239_;
  assign _0254_ = _0163_ ? data_i[1] : _0253_;
  assign sbox_data_o[1] = _0453_ ? _0224_ : _0254_;
  assign _0255_ = data_i[122] & start_i;
  assign _0256_ = _0255_ & _0458_;
  assign _0257_ = _0179_ & data_i[90];
  assign _0258_ = _0183_ & data_i[82];
  assign _0259_ = _0258_ | _0257_;
  assign _0260_ = _0186_ & data_i[74];
  assign _0261_ = _0171_ & data_i[66];
  assign _0262_ = _0261_ | _0260_;
  assign _0263_ = _0262_ | _0259_;
  assign _0264_ = _0453_ & data_i[122];
  assign _0265_ = _0193_ & data_i[114];
  assign _0266_ = _0265_ | _0264_;
  assign _0267_ = _0197_ & data_i[106];
  assign _0268_ = _0168_ & data_i[98];
  assign _0269_ = _0268_ | _0267_;
  assign _0270_ = _0269_ | _0266_;
  assign _0271_ = _0270_ | _0263_;
  assign _0272_ = _0174_ & data_i[10];
  assign _0273_ = _0204_ & data_i[26];
  assign _0274_ = _0206_ & data_i[18];
  assign _0275_ = _0274_ | _0273_;
  assign _0276_ = _0275_ | _0272_;
  assign _0277_ = _0210_ & data_i[58];
  assign _0278_ = _0212_ & data_i[50];
  assign _0279_ = _0278_ | _0277_;
  assign _0280_ = _0215_ & data_i[42];
  assign _0281_ = _0177_ & data_i[34];
  assign _0282_ = _0281_ | _0280_;
  assign _0283_ = _0282_ | _0279_;
  assign _0284_ = _0283_ | _0276_;
  assign _0285_ = _0284_ | _0271_;
  assign _0286_ = _0163_ ? data_i[2] : _0285_;
  assign sbox_data_o[2] = _0453_ ? _0256_ : _0286_;
  assign _0287_ = data_i[123] & start_i;
  assign _0288_ = _0287_ & _0458_;
  assign _0289_ = _0179_ & data_i[91];
  assign _0290_ = _0183_ & data_i[83];
  assign _0291_ = _0290_ | _0289_;
  assign _0292_ = _0186_ & data_i[75];
  assign _0293_ = _0171_ & data_i[67];
  assign _0294_ = _0293_ | _0292_;
  assign _0295_ = _0294_ | _0291_;
  assign _0296_ = _0453_ & data_i[123];
  assign _0297_ = _0193_ & data_i[115];
  assign _0298_ = _0297_ | _0296_;
  assign _0299_ = _0197_ & data_i[107];
  assign _0300_ = _0168_ & data_i[99];
  assign _0301_ = _0300_ | _0299_;
  assign _0302_ = _0301_ | _0298_;
  assign _0303_ = _0302_ | _0295_;
  assign _0304_ = _0174_ & data_i[11];
  assign _0305_ = _0204_ & data_i[27];
  assign _0306_ = _0206_ & data_i[19];
  assign _0307_ = _0306_ | _0305_;
  assign _0308_ = _0307_ | _0304_;
  assign _0309_ = _0210_ & data_i[59];
  assign _0310_ = _0212_ & data_i[51];
  assign _0311_ = _0310_ | _0309_;
  assign _0312_ = _0215_ & data_i[43];
  assign _0313_ = _0177_ & data_i[35];
  assign _0314_ = _0313_ | _0312_;
  assign _0315_ = _0314_ | _0311_;
  assign _0316_ = _0315_ | _0308_;
  assign _0317_ = _0316_ | _0303_;
  assign _0318_ = _0163_ ? data_i[3] : _0317_;
  assign sbox_data_o[3] = _0453_ ? _0288_ : _0318_;
  assign _0319_ = data_i[124] & start_i;
  assign _0320_ = _0319_ & _0458_;
  assign _0321_ = _0179_ & data_i[92];
  assign _0322_ = _0183_ & data_i[84];
  assign _0323_ = _0322_ | _0321_;
  assign _0324_ = _0186_ & data_i[76];
  assign _0325_ = _0171_ & data_i[68];
  assign _0326_ = _0325_ | _0324_;
  assign _0327_ = _0326_ | _0323_;
  assign _0328_ = _0453_ & data_i[124];
  assign _0329_ = _0193_ & data_i[116];
  assign _0330_ = _0329_ | _0328_;
  assign _0331_ = _0197_ & data_i[108];
  assign _0332_ = _0168_ & data_i[100];
  assign _0333_ = _0332_ | _0331_;
  assign _0334_ = _0333_ | _0330_;
  assign _0335_ = _0334_ | _0327_;
  assign _0336_ = _0174_ & data_i[12];
  assign _0337_ = _0204_ & data_i[28];
  assign _0338_ = _0206_ & data_i[20];
  assign _0339_ = _0338_ | _0337_;
  assign _0340_ = _0339_ | _0336_;
  assign _0341_ = _0210_ & data_i[60];
  assign _0342_ = _0212_ & data_i[52];
  assign _0343_ = _0342_ | _0341_;
  assign _0344_ = _0215_ & data_i[44];
  assign _0345_ = _0177_ & data_i[36];
  assign _0346_ = _0345_ | _0344_;
  assign _0347_ = _0346_ | _0343_;
  assign _0348_ = _0347_ | _0340_;
  assign _0349_ = _0348_ | _0335_;
  assign _0350_ = _0163_ ? data_i[4] : _0349_;
  assign sbox_data_o[4] = _0453_ ? _0320_ : _0350_;
  assign _0351_ = data_i[125] & start_i;
  assign _0352_ = _0351_ & _0458_;
  assign _0353_ = _0179_ & data_i[93];
  assign _0354_ = _0183_ & data_i[85];
  assign _0355_ = _0354_ | _0353_;
  assign _0356_ = _0186_ & data_i[77];
  assign _0357_ = _0171_ & data_i[69];
  assign _0358_ = _0357_ | _0356_;
  assign _0359_ = _0358_ | _0355_;
  assign _0360_ = _0453_ & data_i[125];
  assign _0361_ = _0193_ & data_i[117];
  assign _0362_ = _0361_ | _0360_;
  assign _0363_ = _0197_ & data_i[109];
  assign _0364_ = _0168_ & data_i[101];
  assign _0365_ = _0364_ | _0363_;
  assign _0366_ = _0365_ | _0362_;
  assign _0367_ = _0366_ | _0359_;
  assign _0368_ = _0174_ & data_i[13];
  assign _0369_ = _0204_ & data_i[29];
  assign _0370_ = _0206_ & data_i[21];
  assign _0371_ = _0370_ | _0369_;
  assign _0372_ = _0371_ | _0368_;
  assign _0373_ = _0210_ & data_i[61];
  assign _0374_ = _0212_ & data_i[53];
  assign _0375_ = _0374_ | _0373_;
  assign _0376_ = _0215_ & data_i[45];
  assign _0377_ = _0177_ & data_i[37];
  assign _0378_ = _0377_ | _0376_;
  assign _0379_ = _0378_ | _0375_;
  assign _0380_ = _0379_ | _0372_;
  assign _0381_ = _0380_ | _0367_;
  assign _0382_ = _0163_ ? data_i[5] : _0381_;
  assign sbox_data_o[5] = _0453_ ? _0352_ : _0382_;
  assign _0383_ = data_i[126] & start_i;
  assign _0384_ = _0383_ & _0458_;
  assign _0385_ = _0179_ & data_i[94];
  assign _0386_ = _0183_ & data_i[86];
  assign _0387_ = _0386_ | _0385_;
  assign _0388_ = _0186_ & data_i[78];
  assign _0389_ = _0171_ & data_i[70];
  assign _0390_ = _0389_ | _0388_;
  assign _0391_ = _0390_ | _0387_;
  assign _0392_ = _0453_ & data_i[126];
  assign _0393_ = _0193_ & data_i[118];
  assign _0394_ = _0393_ | _0392_;
  assign _0395_ = _0197_ & data_i[110];
  assign _0396_ = _0168_ & data_i[102];
  assign _0397_ = _0396_ | _0395_;
  assign _0398_ = _0397_ | _0394_;
  assign _0399_ = _0398_ | _0391_;
  assign _0400_ = _0174_ & data_i[14];
  assign _0401_ = _0204_ & data_i[30];
  assign _0402_ = _0206_ & data_i[22];
  assign _0403_ = _0402_ | _0401_;
  assign _0404_ = _0403_ | _0400_;
  assign _0405_ = _0210_ & data_i[62];
  assign _0406_ = _0212_ & data_i[54];
  assign _0407_ = _0406_ | _0405_;
  assign _0408_ = _0215_ & data_i[46];
  assign _0409_ = _0177_ & data_i[38];
  assign _0410_ = _0409_ | _0408_;
  assign _0411_ = _0410_ | _0407_;
  assign _0412_ = _0411_ | _0404_;
  assign _0413_ = _0412_ | _0399_;
  assign _0414_ = _0163_ ? data_i[6] : _0413_;
  assign sbox_data_o[6] = _0453_ ? _0384_ : _0414_;
  assign _0415_ = data_i[127] & start_i;
  assign _0416_ = _0415_ & _0458_;
  assign _0417_ = _0179_ & data_i[95];
  assign _0418_ = _0183_ & data_i[87];
  assign _0419_ = _0418_ | _0417_;
  assign _0420_ = _0186_ & data_i[79];
  assign _0421_ = _0171_ & data_i[71];
  assign _0422_ = _0421_ | _0420_;
  assign _0423_ = _0422_ | _0419_;
  assign _0424_ = _0453_ & data_i[127];
  assign _0425_ = _0193_ & data_i[119];
  assign _0426_ = _0425_ | _0424_;
  assign _0427_ = _0197_ & data_i[111];
  assign _0428_ = _0168_ & data_i[103];
  assign _0429_ = _0428_ | _0427_;
  assign _0430_ = _0429_ | _0426_;
  assign _0431_ = _0430_ | _0423_;
  assign _0432_ = _0174_ & data_i[15];
  assign _0433_ = _0204_ & data_i[31];
  assign _0434_ = _0206_ & data_i[23];
  assign _0435_ = _0434_ | _0433_;
  assign _0436_ = _0435_ | _0432_;
  assign _0437_ = _0210_ & data_i[63];
  assign _0438_ = _0212_ & data_i[55];
  assign _0439_ = _0438_ | _0437_;
  assign _0440_ = _0215_ & data_i[47];
  assign _0441_ = _0177_ & data_i[39];
  assign _0442_ = _0441_ | _0440_;
  assign _0443_ = _0442_ | _0439_;
  assign _0444_ = _0443_ | _0436_;
  assign _0445_ = _0444_ | _0431_;
  assign _0446_ = _0163_ ? data_i[7] : _0445_;
  assign sbox_data_o[7] = _0453_ ? _0416_ : _0446_;
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[0] <= 0;
    else
      data_o[0] <= next_data_reg[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[100] <= 0;
    else
      data_o[100] <= next_data_reg[100];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[101] <= 0;
    else
      data_o[101] <= next_data_reg[101];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[102] <= 0;
    else
      data_o[102] <= next_data_reg[102];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[103] <= 0;
    else
      data_o[103] <= next_data_reg[103];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[104] <= 0;
    else
      data_o[104] <= next_data_reg[104];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[105] <= 0;
    else
      data_o[105] <= next_data_reg[105];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[106] <= 0;
    else
      data_o[106] <= next_data_reg[106];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[107] <= 0;
    else
      data_o[107] <= next_data_reg[107];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[108] <= 0;
    else
      data_o[108] <= next_data_reg[108];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[109] <= 0;
    else
      data_o[109] <= next_data_reg[109];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[10] <= 0;
    else
      data_o[10] <= next_data_reg[10];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[110] <= 0;
    else
      data_o[110] <= next_data_reg[110];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[111] <= 0;
    else
      data_o[111] <= next_data_reg[111];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[112] <= 0;
    else
      data_o[112] <= next_data_reg[112];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[113] <= 0;
    else
      data_o[113] <= next_data_reg[113];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[114] <= 0;
    else
      data_o[114] <= next_data_reg[114];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[115] <= 0;
    else
      data_o[115] <= next_data_reg[115];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[116] <= 0;
    else
      data_o[116] <= next_data_reg[116];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[117] <= 0;
    else
      data_o[117] <= next_data_reg[117];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[118] <= 0;
    else
      data_o[118] <= next_data_reg[118];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[119] <= 0;
    else
      data_o[119] <= next_data_reg[119];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[11] <= 0;
    else
      data_o[11] <= next_data_reg[11];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[120] <= 0;
    else
      data_o[120] <= next_data_reg[120];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[121] <= 0;
    else
      data_o[121] <= next_data_reg[121];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[122] <= 0;
    else
      data_o[122] <= next_data_reg[122];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[123] <= 0;
    else
      data_o[123] <= next_data_reg[123];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[124] <= 0;
    else
      data_o[124] <= next_data_reg[124];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[125] <= 0;
    else
      data_o[125] <= next_data_reg[125];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[126] <= 0;
    else
      data_o[126] <= next_data_reg[126];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[127] <= 0;
    else
      data_o[127] <= next_data_reg[127];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[12] <= 0;
    else
      data_o[12] <= next_data_reg[12];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[13] <= 0;
    else
      data_o[13] <= next_data_reg[13];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[14] <= 0;
    else
      data_o[14] <= next_data_reg[14];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[15] <= 0;
    else
      data_o[15] <= next_data_reg[15];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[16] <= 0;
    else
      data_o[16] <= next_data_reg[16];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[17] <= 0;
    else
      data_o[17] <= next_data_reg[17];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[18] <= 0;
    else
      data_o[18] <= next_data_reg[18];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[19] <= 0;
    else
      data_o[19] <= next_data_reg[19];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[1] <= 0;
    else
      data_o[1] <= next_data_reg[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[20] <= 0;
    else
      data_o[20] <= next_data_reg[20];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[21] <= 0;
    else
      data_o[21] <= next_data_reg[21];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[22] <= 0;
    else
      data_o[22] <= next_data_reg[22];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[23] <= 0;
    else
      data_o[23] <= next_data_reg[23];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[24] <= 0;
    else
      data_o[24] <= next_data_reg[24];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[25] <= 0;
    else
      data_o[25] <= next_data_reg[25];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[26] <= 0;
    else
      data_o[26] <= next_data_reg[26];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[27] <= 0;
    else
      data_o[27] <= next_data_reg[27];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[28] <= 0;
    else
      data_o[28] <= next_data_reg[28];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[29] <= 0;
    else
      data_o[29] <= next_data_reg[29];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[2] <= 0;
    else
      data_o[2] <= next_data_reg[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[30] <= 0;
    else
      data_o[30] <= next_data_reg[30];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[31] <= 0;
    else
      data_o[31] <= next_data_reg[31];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[32] <= 0;
    else
      data_o[32] <= next_data_reg[32];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[33] <= 0;
    else
      data_o[33] <= next_data_reg[33];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[34] <= 0;
    else
      data_o[34] <= next_data_reg[34];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[35] <= 0;
    else
      data_o[35] <= next_data_reg[35];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[36] <= 0;
    else
      data_o[36] <= next_data_reg[36];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[37] <= 0;
    else
      data_o[37] <= next_data_reg[37];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[38] <= 0;
    else
      data_o[38] <= next_data_reg[38];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[39] <= 0;
    else
      data_o[39] <= next_data_reg[39];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[3] <= 0;
    else
      data_o[3] <= next_data_reg[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[40] <= 0;
    else
      data_o[40] <= next_data_reg[40];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[41] <= 0;
    else
      data_o[41] <= next_data_reg[41];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[42] <= 0;
    else
      data_o[42] <= next_data_reg[42];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[43] <= 0;
    else
      data_o[43] <= next_data_reg[43];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[44] <= 0;
    else
      data_o[44] <= next_data_reg[44];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[45] <= 0;
    else
      data_o[45] <= next_data_reg[45];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[46] <= 0;
    else
      data_o[46] <= next_data_reg[46];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[47] <= 0;
    else
      data_o[47] <= next_data_reg[47];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[48] <= 0;
    else
      data_o[48] <= next_data_reg[48];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[49] <= 0;
    else
      data_o[49] <= next_data_reg[49];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[4] <= 0;
    else
      data_o[4] <= next_data_reg[4];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[50] <= 0;
    else
      data_o[50] <= next_data_reg[50];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[51] <= 0;
    else
      data_o[51] <= next_data_reg[51];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[52] <= 0;
    else
      data_o[52] <= next_data_reg[52];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[53] <= 0;
    else
      data_o[53] <= next_data_reg[53];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[54] <= 0;
    else
      data_o[54] <= next_data_reg[54];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[55] <= 0;
    else
      data_o[55] <= next_data_reg[55];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[56] <= 0;
    else
      data_o[56] <= next_data_reg[56];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[57] <= 0;
    else
      data_o[57] <= next_data_reg[57];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[58] <= 0;
    else
      data_o[58] <= next_data_reg[58];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[59] <= 0;
    else
      data_o[59] <= next_data_reg[59];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[5] <= 0;
    else
      data_o[5] <= next_data_reg[5];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[60] <= 0;
    else
      data_o[60] <= next_data_reg[60];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[61] <= 0;
    else
      data_o[61] <= next_data_reg[61];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[62] <= 0;
    else
      data_o[62] <= next_data_reg[62];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[63] <= 0;
    else
      data_o[63] <= next_data_reg[63];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[64] <= 0;
    else
      data_o[64] <= next_data_reg[64];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[65] <= 0;
    else
      data_o[65] <= next_data_reg[65];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[66] <= 0;
    else
      data_o[66] <= next_data_reg[66];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[67] <= 0;
    else
      data_o[67] <= next_data_reg[67];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[68] <= 0;
    else
      data_o[68] <= next_data_reg[68];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[69] <= 0;
    else
      data_o[69] <= next_data_reg[69];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[6] <= 0;
    else
      data_o[6] <= next_data_reg[6];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[70] <= 0;
    else
      data_o[70] <= next_data_reg[70];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[71] <= 0;
    else
      data_o[71] <= next_data_reg[71];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[72] <= 0;
    else
      data_o[72] <= next_data_reg[72];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[73] <= 0;
    else
      data_o[73] <= next_data_reg[73];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[74] <= 0;
    else
      data_o[74] <= next_data_reg[74];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[75] <= 0;
    else
      data_o[75] <= next_data_reg[75];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[76] <= 0;
    else
      data_o[76] <= next_data_reg[76];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[77] <= 0;
    else
      data_o[77] <= next_data_reg[77];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[78] <= 0;
    else
      data_o[78] <= next_data_reg[78];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[79] <= 0;
    else
      data_o[79] <= next_data_reg[79];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[7] <= 0;
    else
      data_o[7] <= next_data_reg[7];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[80] <= 0;
    else
      data_o[80] <= next_data_reg[80];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[81] <= 0;
    else
      data_o[81] <= next_data_reg[81];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[82] <= 0;
    else
      data_o[82] <= next_data_reg[82];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[83] <= 0;
    else
      data_o[83] <= next_data_reg[83];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[84] <= 0;
    else
      data_o[84] <= next_data_reg[84];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[85] <= 0;
    else
      data_o[85] <= next_data_reg[85];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[86] <= 0;
    else
      data_o[86] <= next_data_reg[86];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[87] <= 0;
    else
      data_o[87] <= next_data_reg[87];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[88] <= 0;
    else
      data_o[88] <= next_data_reg[88];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[89] <= 0;
    else
      data_o[89] <= next_data_reg[89];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[8] <= 0;
    else
      data_o[8] <= next_data_reg[8];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[90] <= 0;
    else
      data_o[90] <= next_data_reg[90];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[91] <= 0;
    else
      data_o[91] <= next_data_reg[91];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[92] <= 0;
    else
      data_o[92] <= next_data_reg[92];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[93] <= 0;
    else
      data_o[93] <= next_data_reg[93];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[94] <= 0;
    else
      data_o[94] <= next_data_reg[94];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[95] <= 0;
    else
      data_o[95] <= next_data_reg[95];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[96] <= 0;
    else
      data_o[96] <= next_data_reg[96];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[97] <= 0;
    else
      data_o[97] <= next_data_reg[97];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[98] <= 0;
    else
      data_o[98] <= next_data_reg[98];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[99] <= 0;
    else
      data_o[99] <= next_data_reg[99];
  always @(posedge clk or negedge reset)
    if (!reset)
      data_o[9] <= 0;
    else
      data_o[9] <= next_data_reg[9];
  always @(posedge clk or negedge reset)
    if (!reset)
      ready_o <= 0;
    else
      ready_o <= next_ready_o;
  always @(posedge clk or negedge reset)
    if (!reset)
      state[0] <= 0;
    else
      state[0] <= next_state[0];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[1] <= 0;
    else
      state[1] <= next_state[1];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[2] <= 0;
    else
      state[2] <= next_state[2];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[3] <= 0;
    else
      state[3] <= next_state[3];
  always @(posedge clk or negedge reset)
    if (!reset)
      state[4] <= 0;
    else
      state[4] <= next_state[4];
  assign \data_array[0]  = data_i[127:120];
  assign \data_array[10]  = data_i[47:40];
  assign \data_array[11]  = data_i[39:32];
  assign \data_array[12]  = data_i[31:24];
  assign \data_array[13]  = data_i[23:16];
  assign \data_array[14]  = data_i[15:8];
  assign \data_array[15]  = data_i[7:0];
  assign \data_array[1]  = data_i[119:112];
  assign \data_array[2]  = data_i[111:104];
  assign \data_array[3]  = data_i[103:96];
  assign \data_array[4]  = data_i[95:88];
  assign \data_array[5]  = data_i[87:80];
  assign \data_array[6]  = data_i[79:72];
  assign \data_array[7]  = data_i[71:64];
  assign \data_array[8]  = data_i[63:56];
  assign \data_array[9]  = data_i[55:48];
  assign data_i_var = data_i;
  assign data_reg = data_o;
  assign sbox_decrypt_o = decrypt_i;
endmodule

module word_mixcolum(in, outx, outy);
  wire [7:0] a;
  wire [7:0] b;
  wire [7:0] c;
  wire [7:0] d;
  input [31:0] in;
  wire [31:0] in_var;
  output [31:0] outx;
  wire [31:0] outx_var;
  output [31:0] outy;
  wire [31:0] outy_var;
  wire [7:0] x1;
  wire [7:0] x2;
  wire [7:0] x3;
  wire [7:0] x4;
  wire [7:0] y1;
  wire [7:0] y2;
  wire [7:0] y3;
  wire [7:0] y4;
  byte_mixcolum bm1 (
    .a(in[31:24]),
    .b(in[23:16]),
    .c(in[15:8]),
    .d(in[7:0]),
    .outx(outx[31:24]),
    .outy(outy[31:24])
  );
  byte_mixcolum bm2 (
    .a(in[23:16]),
    .b(in[15:8]),
    .c(in[7:0]),
    .d(in[31:24]),
    .outx(outx[23:16]),
    .outy(outy[23:16])
  );
  byte_mixcolum bm3 (
    .a(in[15:8]),
    .b(in[7:0]),
    .c(in[31:24]),
    .d(in[23:16]),
    .outx(outx[15:8]),
    .outy(outy[15:8])
  );
  byte_mixcolum bm4 (
    .a(in[7:0]),
    .b(in[31:24]),
    .c(in[23:16]),
    .d(in[15:8]),
    .outx(outx[7:0]),
    .outy(outy[7:0])
  );
  assign a = in[31:24];
  assign b = in[23:16];
  assign c = in[15:8];
  assign d = in[7:0];
  assign in_var = in;
  assign outx_var = outx;
  assign outy_var = outy;
  assign x1 = outx[31:24];
  assign x2 = outx[23:16];
  assign x3 = outx[15:8];
  assign x4 = outx[7:0];
  assign y1 = outy[31:24];
  assign y2 = outy[23:16];
  assign y3 = outy[15:8];
  assign y4 = outy[7:0];
endmodule
