/*
:name: 22.7--timescale-basic-4
:description: Test
:should_fail: 1
:tags: 22.7
:type: preprocessing
*/
`timescale 1 ns / 1000 ps
