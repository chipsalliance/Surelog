/*
:name: 22.9--unconnected_drive-basic
:description: Test
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull1
`nounconnected_drive
