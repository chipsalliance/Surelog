// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: timescale-directive
:description: Set timescale
:tags: 5.6.4
*/

`timescale 1 ns / 1 ps

module ts();
endmodule
