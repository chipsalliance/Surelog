module top();
   
endmodule
