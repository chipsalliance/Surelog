/*
:name: typedef_test_9
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef data_t my_array_t [k:0][j:0];