/*
:name: class_member_test_44
:description: Test
:tags: 8.3
*/
class constructible;
extern function new;
endclass