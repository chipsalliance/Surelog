/*
:name: class_member_test_50
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
virtual hinterface.some_mod_port winterface;
virtual interface foo_if #(J,K) bar_if, baz_if;
virtual disinterface#(.N(N)).some_mod_port blinterface;
endclass