// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: non_blocking_assignment
:description: non-blocking assignment test
:tags: 10.4.2
*/
module top();

logic a;

initial begin
	a <= 2;
end

endmodule
