// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: iface_class_test_2
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic #(int N = 8, type T = string);
endclass

module test;
endmodule
