// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: class_member_test_26
:description: Test
:tags: 8.3
*/
virtual class myclass;
pure virtual function integer subroutine;
pure virtual function integer compute(int a, bit b);
endclass

module test;
endmodule
