/*
:name: class_member_test_17
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function yourpkg::classy::xtype #(p,q) subr;
endclass