/*
:name: class_member_test_0
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
task subtask;
endtask
endclass