/*
:name: class_test_66
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
  int num_packets;
`ifdef DEBUGGER
  string source_name;
  string dest_name;
`elsif LAZY
`endif
  int router_size;
endclass