module aes_cipher_top(clk, rst, ld, done, key, text_in, text_out);
  wire [3:0] _0000_;
  wire _0001_;
  wire [7:0] _0002_;
  wire [7:0] _0003_;
  wire [7:0] _0004_;
  wire [7:0] _0005_;
  wire [7:0] _0006_;
  wire [7:0] _0007_;
  wire [7:0] _0008_;
  wire [7:0] _0009_;
  wire [7:0] _0010_;
  wire [7:0] _0011_;
  wire [7:0] _0012_;
  wire [7:0] _0013_;
  wire [7:0] _0014_;
  wire [7:0] _0015_;
  wire [7:0] _0016_;
  wire [7:0] _0017_;
  wire [127:0] _0018_;
  wire [7:0] _0019_;
  wire [7:0] _0020_;
  wire [7:0] _0021_;
  wire [7:0] _0022_;
  wire [7:0] _0023_;
  wire [7:0] _0024_;
  wire [7:0] _0025_;
  wire [7:0] _0026_;
  wire [7:0] _0027_;
  wire [7:0] _0028_;
  wire [7:0] _0029_;
  wire [7:0] _0030_;
  wire [7:0] _0031_;
  wire [7:0] _0032_;
  wire [7:0] _0033_;
  wire [7:0] _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  input clk;
  reg [3:0] dcnt;
  output done;
  reg done;
  input [127:0] key;
  input ld;
  reg ld_r;
  input rst;
  reg [7:0] sa00;
  wire [7:0] sa00_sr;
  wire [7:0] sa00_sub;
  reg [7:0] sa01;
  wire [7:0] sa01_sr;
  wire [7:0] sa01_sub;
  reg [7:0] sa02;
  wire [7:0] sa02_sr;
  wire [7:0] sa02_sub;
  reg [7:0] sa03;
  wire [7:0] sa03_sr;
  wire [7:0] sa03_sub;
  reg [7:0] sa10;
  wire [7:0] sa10_sr;
  wire [7:0] sa10_sub;
  reg [7:0] sa11;
  wire [7:0] sa11_sr;
  wire [7:0] sa11_sub;
  reg [7:0] sa12;
  wire [7:0] sa12_sr;
  wire [7:0] sa12_sub;
  reg [7:0] sa13;
  wire [7:0] sa13_sr;
  wire [7:0] sa13_sub;
  reg [7:0] sa20;
  wire [7:0] sa20_sr;
  wire [7:0] sa20_sub;
  reg [7:0] sa21;
  wire [7:0] sa21_sr;
  wire [7:0] sa21_sub;
  reg [7:0] sa22;
  wire [7:0] sa22_sr;
  wire [7:0] sa22_sub;
  reg [7:0] sa23;
  wire [7:0] sa23_sr;
  wire [7:0] sa23_sub;
  reg [7:0] sa30;
  wire [7:0] sa30_sr;
  wire [7:0] sa30_sub;
  reg [7:0] sa31;
  wire [7:0] sa31_sr;
  wire [7:0] sa31_sub;
  reg [7:0] sa32;
  wire [7:0] sa32_sr;
  wire [7:0] sa32_sub;
  reg [7:0] sa33;
  wire [7:0] sa33_sr;
  wire [7:0] sa33_sub;
  input [127:0] text_in;
  reg [127:0] text_in_r;
  output [127:0] text_out;
  reg [127:0] text_out;
  wire [31:0] w0;
  wire [31:0] w1;
  wire [31:0] w2;
  wire [31:0] w3;
  assign _0979_ = ~ld;
  assign _0980_ = _0979_ & dcnt[0];
  assign _0981_ = ~dcnt[3];
  assign _0982_ = ~dcnt[1];
  assign _0983_ = ~dcnt[2];
  assign _0984_ = _0983_ & _0982_;
  assign _0985_ = _0984_ & _0981_;
  assign _0001_ = _0985_ & _0980_;
  assign _0986_ = dcnt[1] | dcnt[0];
  assign _0987_ = dcnt[3] | dcnt[2];
  assign _0988_ = _0987_ | _0986_;
  assign _0989_ = _0988_ ^ dcnt[0];
  assign _0990_ = _0989_ | ld;
  assign _0000_[0] = _0990_ & rst;
  assign _0991_ = _0982_ ^ dcnt[0];
  assign _0992_ = _0988_ ? _0991_ : dcnt[1];
  assign _0993_ = _0992_ | ld;
  assign _0000_[1] = _0993_ & rst;
  assign _0994_ = _0986_ ^ _0983_;
  assign _0995_ = _0988_ ? _0994_ : dcnt[2];
  assign _0996_ = _0979_ & rst;
  assign _0000_[2] = _0996_ & _0995_;
  assign _0997_ = _0986_ | dcnt[2];
  assign _0998_ = _0997_ ^ _0981_;
  assign _0999_ = _0988_ ? _0998_ : dcnt[3];
  assign _1000_ = _0999_ | ld;
  assign _0000_[3] = _1000_ & rst;
  assign _0018_[0] = ld ? text_in[0] : text_in_r[0];
  assign _0018_[100] = ld ? text_in[100] : text_in_r[100];
  assign _0018_[101] = ld ? text_in[101] : text_in_r[101];
  assign _0018_[102] = ld ? text_in[102] : text_in_r[102];
  assign _0018_[103] = ld ? text_in[103] : text_in_r[103];
  assign _0018_[104] = ld ? text_in[104] : text_in_r[104];
  assign _0018_[105] = ld ? text_in[105] : text_in_r[105];
  assign _0018_[106] = ld ? text_in[106] : text_in_r[106];
  assign _0018_[107] = ld ? text_in[107] : text_in_r[107];
  assign _0018_[108] = ld ? text_in[108] : text_in_r[108];
  assign _0018_[109] = ld ? text_in[109] : text_in_r[109];
  assign _0018_[10] = ld ? text_in[10] : text_in_r[10];
  assign _0018_[110] = ld ? text_in[110] : text_in_r[110];
  assign _0018_[111] = ld ? text_in[111] : text_in_r[111];
  assign _0018_[112] = ld ? text_in[112] : text_in_r[112];
  assign _0018_[113] = ld ? text_in[113] : text_in_r[113];
  assign _0018_[114] = ld ? text_in[114] : text_in_r[114];
  assign _0018_[115] = ld ? text_in[115] : text_in_r[115];
  assign _0018_[116] = ld ? text_in[116] : text_in_r[116];
  assign _0018_[117] = ld ? text_in[117] : text_in_r[117];
  assign _0018_[118] = ld ? text_in[118] : text_in_r[118];
  assign _0018_[119] = ld ? text_in[119] : text_in_r[119];
  assign _0018_[11] = ld ? text_in[11] : text_in_r[11];
  assign _0018_[120] = ld ? text_in[120] : text_in_r[120];
  assign _0018_[121] = ld ? text_in[121] : text_in_r[121];
  assign _0018_[122] = ld ? text_in[122] : text_in_r[122];
  assign _0018_[123] = ld ? text_in[123] : text_in_r[123];
  assign _0018_[124] = ld ? text_in[124] : text_in_r[124];
  assign _0018_[125] = ld ? text_in[125] : text_in_r[125];
  assign _0018_[126] = ld ? text_in[126] : text_in_r[126];
  assign _0018_[127] = ld ? text_in[127] : text_in_r[127];
  assign _0018_[12] = ld ? text_in[12] : text_in_r[12];
  assign _0018_[13] = ld ? text_in[13] : text_in_r[13];
  assign _0018_[14] = ld ? text_in[14] : text_in_r[14];
  assign _0018_[15] = ld ? text_in[15] : text_in_r[15];
  assign _0018_[16] = ld ? text_in[16] : text_in_r[16];
  assign _0018_[17] = ld ? text_in[17] : text_in_r[17];
  assign _0018_[18] = ld ? text_in[18] : text_in_r[18];
  assign _0018_[19] = ld ? text_in[19] : text_in_r[19];
  assign _0018_[1] = ld ? text_in[1] : text_in_r[1];
  assign _0018_[20] = ld ? text_in[20] : text_in_r[20];
  assign _0018_[21] = ld ? text_in[21] : text_in_r[21];
  assign _0018_[22] = ld ? text_in[22] : text_in_r[22];
  assign _0018_[23] = ld ? text_in[23] : text_in_r[23];
  assign _0018_[24] = ld ? text_in[24] : text_in_r[24];
  assign _0018_[25] = ld ? text_in[25] : text_in_r[25];
  assign _0018_[26] = ld ? text_in[26] : text_in_r[26];
  assign _0018_[27] = ld ? text_in[27] : text_in_r[27];
  assign _0018_[28] = ld ? text_in[28] : text_in_r[28];
  assign _0018_[29] = ld ? text_in[29] : text_in_r[29];
  assign _0018_[2] = ld ? text_in[2] : text_in_r[2];
  assign _0018_[30] = ld ? text_in[30] : text_in_r[30];
  assign _0018_[31] = ld ? text_in[31] : text_in_r[31];
  assign _0018_[32] = ld ? text_in[32] : text_in_r[32];
  assign _0018_[33] = ld ? text_in[33] : text_in_r[33];
  assign _0018_[34] = ld ? text_in[34] : text_in_r[34];
  assign _0018_[35] = ld ? text_in[35] : text_in_r[35];
  assign _0018_[36] = ld ? text_in[36] : text_in_r[36];
  assign _0018_[37] = ld ? text_in[37] : text_in_r[37];
  assign _0018_[38] = ld ? text_in[38] : text_in_r[38];
  assign _0018_[39] = ld ? text_in[39] : text_in_r[39];
  assign _0018_[3] = ld ? text_in[3] : text_in_r[3];
  assign _0018_[40] = ld ? text_in[40] : text_in_r[40];
  assign _0018_[41] = ld ? text_in[41] : text_in_r[41];
  assign _0018_[42] = ld ? text_in[42] : text_in_r[42];
  assign _0018_[43] = ld ? text_in[43] : text_in_r[43];
  assign _0018_[44] = ld ? text_in[44] : text_in_r[44];
  assign _0018_[45] = ld ? text_in[45] : text_in_r[45];
  assign _0018_[46] = ld ? text_in[46] : text_in_r[46];
  assign _0018_[47] = ld ? text_in[47] : text_in_r[47];
  assign _0018_[48] = ld ? text_in[48] : text_in_r[48];
  assign _0018_[49] = ld ? text_in[49] : text_in_r[49];
  assign _0018_[4] = ld ? text_in[4] : text_in_r[4];
  assign _0018_[50] = ld ? text_in[50] : text_in_r[50];
  assign _0018_[51] = ld ? text_in[51] : text_in_r[51];
  assign _0018_[52] = ld ? text_in[52] : text_in_r[52];
  assign _0018_[53] = ld ? text_in[53] : text_in_r[53];
  assign _0018_[54] = ld ? text_in[54] : text_in_r[54];
  assign _0018_[55] = ld ? text_in[55] : text_in_r[55];
  assign _0018_[56] = ld ? text_in[56] : text_in_r[56];
  assign _0018_[57] = ld ? text_in[57] : text_in_r[57];
  assign _0018_[58] = ld ? text_in[58] : text_in_r[58];
  assign _0018_[59] = ld ? text_in[59] : text_in_r[59];
  assign _0018_[5] = ld ? text_in[5] : text_in_r[5];
  assign _0018_[60] = ld ? text_in[60] : text_in_r[60];
  assign _0018_[61] = ld ? text_in[61] : text_in_r[61];
  assign _0018_[62] = ld ? text_in[62] : text_in_r[62];
  assign _0018_[63] = ld ? text_in[63] : text_in_r[63];
  assign _0018_[64] = ld ? text_in[64] : text_in_r[64];
  assign _0018_[65] = ld ? text_in[65] : text_in_r[65];
  assign _0018_[66] = ld ? text_in[66] : text_in_r[66];
  assign _0018_[67] = ld ? text_in[67] : text_in_r[67];
  assign _0018_[68] = ld ? text_in[68] : text_in_r[68];
  assign _0018_[69] = ld ? text_in[69] : text_in_r[69];
  assign _0018_[6] = ld ? text_in[6] : text_in_r[6];
  assign _0018_[70] = ld ? text_in[70] : text_in_r[70];
  assign _0018_[71] = ld ? text_in[71] : text_in_r[71];
  assign _0018_[72] = ld ? text_in[72] : text_in_r[72];
  assign _0018_[73] = ld ? text_in[73] : text_in_r[73];
  assign _0018_[74] = ld ? text_in[74] : text_in_r[74];
  assign _0018_[75] = ld ? text_in[75] : text_in_r[75];
  assign _0018_[76] = ld ? text_in[76] : text_in_r[76];
  assign _0018_[77] = ld ? text_in[77] : text_in_r[77];
  assign _0018_[78] = ld ? text_in[78] : text_in_r[78];
  assign _0018_[79] = ld ? text_in[79] : text_in_r[79];
  assign _0018_[7] = ld ? text_in[7] : text_in_r[7];
  assign _0018_[80] = ld ? text_in[80] : text_in_r[80];
  assign _0018_[81] = ld ? text_in[81] : text_in_r[81];
  assign _0018_[82] = ld ? text_in[82] : text_in_r[82];
  assign _0018_[83] = ld ? text_in[83] : text_in_r[83];
  assign _0018_[84] = ld ? text_in[84] : text_in_r[84];
  assign _0018_[85] = ld ? text_in[85] : text_in_r[85];
  assign _0018_[86] = ld ? text_in[86] : text_in_r[86];
  assign _0018_[87] = ld ? text_in[87] : text_in_r[87];
  assign _0018_[88] = ld ? text_in[88] : text_in_r[88];
  assign _0018_[89] = ld ? text_in[89] : text_in_r[89];
  assign _0018_[8] = ld ? text_in[8] : text_in_r[8];
  assign _0018_[90] = ld ? text_in[90] : text_in_r[90];
  assign _0018_[91] = ld ? text_in[91] : text_in_r[91];
  assign _0018_[92] = ld ? text_in[92] : text_in_r[92];
  assign _0018_[93] = ld ? text_in[93] : text_in_r[93];
  assign _0018_[94] = ld ? text_in[94] : text_in_r[94];
  assign _0018_[95] = ld ? text_in[95] : text_in_r[95];
  assign _0018_[96] = ld ? text_in[96] : text_in_r[96];
  assign _0018_[97] = ld ? text_in[97] : text_in_r[97];
  assign _0018_[98] = ld ? text_in[98] : text_in_r[98];
  assign _0018_[99] = ld ? text_in[99] : text_in_r[99];
  assign _0018_[9] = ld ? text_in[9] : text_in_r[9];
  assign _0035_ = w3[0] ^ text_in_r[0];
  assign _0036_ = ~w3[0];
  assign _0037_ = ~sa10_sub[0];
  assign _0038_ = sa03_sr[7] ^ sa03_sr[0];
  assign _0039_ = _0038_ ^ _0037_;
  assign _0040_ = _0039_ ^ sa21_sub[0];
  assign _0041_ = _0040_ ^ sa32_sub[7];
  assign _0042_ = _0041_ ^ _0036_;
  assign _0017_[0] = ld_r ? _0035_ : _0042_;
  assign _0043_ = w3[1] ^ text_in_r[1];
  assign _0044_ = ~sa03_sr[1];
  assign _0045_ = _0038_ ^ _0044_;
  assign _0046_ = _0045_ ^ sa10_sub[1];
  assign _0047_ = _0046_ ^ sa21_sub[1];
  assign _0048_ = ~sa32_sub[0];
  assign _0049_ = sa32_sub[7] ^ _0048_;
  assign _0050_ = _0049_ ^ _0047_;
  assign _0051_ = _0050_ ^ w3[1];
  assign _0017_[1] = ld_r ? _0043_ : _0051_;
  assign _0052_ = w3[2] ^ text_in_r[2];
  assign _0053_ = ~w3[2];
  assign _0054_ = ~sa10_sub[2];
  assign _0055_ = sa03_sr[2] ^ sa03_sr[1];
  assign _0056_ = _0055_ ^ _0054_;
  assign _0057_ = _0056_ ^ sa21_sub[2];
  assign _0058_ = _0057_ ^ sa32_sub[1];
  assign _0059_ = _0058_ ^ _0053_;
  assign _0017_[2] = ld_r ? _0052_ : _0059_;
  assign _0060_ = w3[3] ^ text_in_r[3];
  assign _0061_ = ~w3[3];
  assign _0062_ = ~sa10_sub[3];
  assign _0063_ = ~sa03_sr[3];
  assign _0064_ = sa03_sr[7] ^ sa03_sr[2];
  assign _0065_ = _0064_ ^ _0063_;
  assign _0066_ = _0065_ ^ _0062_;
  assign _0067_ = _0066_ ^ sa21_sub[3];
  assign _0068_ = ~sa32_sub[2];
  assign _0069_ = sa32_sub[7] ^ _0068_;
  assign _0070_ = _0069_ ^ _0067_;
  assign _0071_ = _0070_ ^ _0061_;
  assign _0017_[3] = ld_r ? _0060_ : _0071_;
  assign _0072_ = w3[4] ^ text_in_r[4];
  assign _0073_ = ~sa03_sr[4];
  assign _0074_ = sa03_sr[7] ^ sa03_sr[3];
  assign _0075_ = _0074_ ^ _0073_;
  assign _0076_ = _0075_ ^ sa10_sub[4];
  assign _0077_ = _0076_ ^ sa21_sub[4];
  assign _0078_ = ~sa32_sub[3];
  assign _0079_ = sa32_sub[7] ^ _0078_;
  assign _0080_ = _0079_ ^ _0077_;
  assign _0081_ = _0080_ ^ w3[4];
  assign _0017_[4] = ld_r ? _0072_ : _0081_;
  assign _0082_ = w3[5] ^ text_in_r[5];
  assign _0083_ = ~w3[5];
  assign _0084_ = ~sa10_sub[5];
  assign _0085_ = sa03_sr[5] ^ sa03_sr[4];
  assign _0086_ = _0085_ ^ _0084_;
  assign _0087_ = _0086_ ^ sa21_sub[5];
  assign _0088_ = _0087_ ^ sa32_sub[4];
  assign _0089_ = _0088_ ^ _0083_;
  assign _0017_[5] = ld_r ? _0082_ : _0089_;
  assign _0090_ = w3[6] ^ text_in_r[6];
  assign _0091_ = ~w3[6];
  assign _0092_ = ~sa10_sub[6];
  assign _0093_ = sa03_sr[6] ^ sa03_sr[5];
  assign _0094_ = _0093_ ^ _0092_;
  assign _0095_ = _0094_ ^ sa21_sub[6];
  assign _0096_ = _0095_ ^ sa32_sub[5];
  assign _0097_ = _0096_ ^ _0091_;
  assign _0017_[6] = ld_r ? _0090_ : _0097_;
  assign _0098_ = w3[7] ^ text_in_r[7];
  assign _0099_ = ~w3[7];
  assign _0100_ = ~sa10_sub[7];
  assign _0101_ = sa03_sr[7] ^ sa03_sr[6];
  assign _0102_ = _0101_ ^ _0100_;
  assign _0103_ = _0102_ ^ sa21_sub[7];
  assign _0104_ = _0103_ ^ sa32_sub[6];
  assign _0105_ = _0104_ ^ _0099_;
  assign _0017_[7] = ld_r ? _0098_ : _0105_;
  assign _0106_ = w3[8] ^ text_in_r[8];
  assign _0107_ = ~sa21_sub[7];
  assign _0108_ = sa10_sub[0] ^ sa03_sr[0];
  assign _0109_ = _0108_ ^ _0107_;
  assign _0110_ = _0109_ ^ sa32_sub[7];
  assign _0111_ = _0110_ ^ _0048_;
  assign _0112_ = _0111_ ^ w3[8];
  assign _0013_[0] = ld_r ? _0106_ : _0112_;
  assign _0113_ = w3[9] ^ text_in_r[9];
  assign _0114_ = ~w3[9];
  assign _0115_ = sa10_sub[1] ^ sa03_sr[1];
  assign _0116_ = sa21_sub[7] ^ sa21_sub[0];
  assign _0117_ = _0116_ ^ _0115_;
  assign _0118_ = _0117_ ^ _0049_;
  assign _0119_ = _0118_ ^ sa32_sub[1];
  assign _0120_ = _0119_ ^ _0114_;
  assign _0013_[1] = ld_r ? _0113_ : _0120_;
  assign _0121_ = w3[10] ^ text_in_r[10];
  assign _0122_ = ~sa21_sub[1];
  assign _0123_ = sa10_sub[2] ^ sa03_sr[2];
  assign _0124_ = _0123_ ^ _0122_;
  assign _0125_ = _0124_ ^ sa32_sub[1];
  assign _0126_ = _0125_ ^ _0068_;
  assign _0127_ = _0126_ ^ w3[10];
  assign _0013_[2] = ld_r ? _0121_ : _0127_;
  assign _0128_ = w3[11] ^ text_in_r[11];
  assign _0129_ = sa10_sub[3] ^ sa03_sr[3];
  assign _0130_ = sa21_sub[7] ^ sa21_sub[2];
  assign _0131_ = _0130_ ^ _0129_;
  assign _0132_ = _0131_ ^ _0069_;
  assign _0133_ = _0132_ ^ _0078_;
  assign _0134_ = _0133_ ^ w3[11];
  assign _0013_[3] = ld_r ? _0128_ : _0134_;
  assign _0135_ = w3[12] ^ text_in_r[12];
  assign _0136_ = ~w3[12];
  assign _0137_ = sa10_sub[4] ^ sa03_sr[4];
  assign _0138_ = sa21_sub[7] ^ sa21_sub[3];
  assign _0139_ = _0138_ ^ _0137_;
  assign _0140_ = _0139_ ^ _0079_;
  assign _0141_ = _0140_ ^ sa32_sub[4];
  assign _0142_ = _0141_ ^ _0136_;
  assign _0013_[4] = ld_r ? _0135_ : _0142_;
  assign _0143_ = w3[13] ^ text_in_r[13];
  assign _0144_ = ~w3[13];
  assign _0145_ = ~sa21_sub[4];
  assign _0146_ = sa10_sub[5] ^ sa03_sr[5];
  assign _0147_ = _0146_ ^ _0145_;
  assign _0148_ = _0147_ ^ sa32_sub[4];
  assign _0149_ = _0148_ ^ sa32_sub[5];
  assign _0150_ = _0149_ ^ _0144_;
  assign _0013_[5] = ld_r ? _0143_ : _0150_;
  assign _0151_ = w3[14] ^ text_in_r[14];
  assign _0152_ = ~w3[14];
  assign _0153_ = ~sa21_sub[5];
  assign _0154_ = sa10_sub[6] ^ sa03_sr[6];
  assign _0155_ = _0154_ ^ _0153_;
  assign _0156_ = _0155_ ^ sa32_sub[5];
  assign _0157_ = _0156_ ^ sa32_sub[6];
  assign _0158_ = _0157_ ^ _0152_;
  assign _0013_[6] = ld_r ? _0151_ : _0158_;
  assign _0159_ = w3[15] ^ text_in_r[15];
  assign _0160_ = ~w3[15];
  assign _0161_ = ~sa21_sub[6];
  assign _0162_ = sa10_sub[7] ^ sa03_sr[7];
  assign _0163_ = _0162_ ^ _0161_;
  assign _0164_ = _0163_ ^ sa32_sub[6];
  assign _0165_ = _0164_ ^ sa32_sub[7];
  assign _0166_ = _0165_ ^ _0160_;
  assign _0013_[7] = ld_r ? _0159_ : _0166_;
  assign _0167_ = w3[16] ^ text_in_r[16];
  assign _0168_ = sa10_sub[7] ^ sa03_sr[0];
  assign _0169_ = _0168_ ^ _0107_;
  assign _0170_ = _0169_ ^ sa21_sub[0];
  assign _0171_ = _0170_ ^ _0048_;
  assign _0172_ = _0171_ ^ w3[16];
  assign _0009_[0] = ld_r ? _0167_ : _0172_;
  assign _0173_ = w3[17] ^ text_in_r[17];
  assign _0174_ = ~w3[17];
  assign _0175_ = sa10_sub[7] ^ sa10_sub[0];
  assign _0176_ = _0175_ ^ _0044_;
  assign _0177_ = _0176_ ^ _0116_;
  assign _0178_ = _0177_ ^ sa21_sub[1];
  assign _0179_ = _0178_ ^ sa32_sub[1];
  assign _0180_ = _0179_ ^ _0174_;
  assign _0009_[1] = ld_r ? _0173_ : _0180_;
  assign _0181_ = w3[18] ^ text_in_r[18];
  assign _0182_ = sa10_sub[1] ^ sa03_sr[2];
  assign _0183_ = _0182_ ^ _0122_;
  assign _0184_ = _0183_ ^ sa21_sub[2];
  assign _0185_ = _0184_ ^ _0068_;
  assign _0186_ = _0185_ ^ w3[18];
  assign _0009_[2] = ld_r ? _0181_ : _0186_;
  assign _0187_ = w3[19] ^ text_in_r[19];
  assign _0188_ = sa10_sub[7] ^ sa10_sub[2];
  assign _0189_ = _0188_ ^ _0063_;
  assign _0190_ = _0189_ ^ _0130_;
  assign _0191_ = _0190_ ^ sa21_sub[3];
  assign _0192_ = _0191_ ^ _0078_;
  assign _0193_ = _0192_ ^ w3[19];
  assign _0009_[3] = ld_r ? _0187_ : _0193_;
  assign _0194_ = w3[20] ^ text_in_r[20];
  assign _0195_ = ~w3[20];
  assign _0196_ = sa10_sub[7] ^ sa10_sub[3];
  assign _0197_ = _0196_ ^ _0073_;
  assign _0198_ = _0197_ ^ _0138_;
  assign _0199_ = _0198_ ^ sa21_sub[4];
  assign _0200_ = _0199_ ^ sa32_sub[4];
  assign _0201_ = _0200_ ^ _0195_;
  assign _0009_[4] = ld_r ? _0194_ : _0201_;
  assign _0202_ = w3[21] ^ text_in_r[21];
  assign _0203_ = ~w3[21];
  assign _0204_ = sa10_sub[4] ^ sa03_sr[5];
  assign _0205_ = _0204_ ^ _0145_;
  assign _0206_ = _0205_ ^ sa21_sub[5];
  assign _0207_ = _0206_ ^ sa32_sub[5];
  assign _0208_ = _0207_ ^ _0203_;
  assign _0009_[5] = ld_r ? _0202_ : _0208_;
  assign _0209_ = w3[22] ^ text_in_r[22];
  assign _0210_ = ~w3[22];
  assign _0211_ = sa10_sub[5] ^ sa03_sr[6];
  assign _0212_ = _0211_ ^ _0153_;
  assign _0213_ = _0212_ ^ sa21_sub[6];
  assign _0214_ = _0213_ ^ sa32_sub[6];
  assign _0215_ = _0214_ ^ _0210_;
  assign _0009_[6] = ld_r ? _0209_ : _0215_;
  assign _0216_ = w3[23] ^ text_in_r[23];
  assign _0217_ = ~w3[23];
  assign _0218_ = sa10_sub[6] ^ sa03_sr[7];
  assign _0219_ = _0218_ ^ _0161_;
  assign _0220_ = _0219_ ^ sa21_sub[7];
  assign _0221_ = _0220_ ^ sa32_sub[7];
  assign _0222_ = _0221_ ^ _0217_;
  assign _0009_[7] = ld_r ? _0216_ : _0222_;
  assign _0223_ = w3[24] ^ text_in_r[24];
  assign _0224_ = _0162_ ^ _0037_;
  assign _0225_ = _0224_ ^ sa21_sub[0];
  assign _0226_ = _0225_ ^ _0048_;
  assign _0227_ = _0226_ ^ w3[24];
  assign _0005_[0] = ld_r ? _0223_ : _0227_;
  assign _0228_ = w3[25] ^ text_in_r[25];
  assign _0229_ = ~w3[25];
  assign _0230_ = _0175_ ^ _0038_;
  assign _0231_ = _0230_ ^ sa10_sub[1];
  assign _0232_ = _0231_ ^ _0122_;
  assign _0233_ = _0232_ ^ sa32_sub[1];
  assign _0234_ = _0233_ ^ _0229_;
  assign _0005_[1] = ld_r ? _0228_ : _0234_;
  assign _0235_ = w3[26] ^ text_in_r[26];
  assign _0236_ = _0115_ ^ _0054_;
  assign _0237_ = _0236_ ^ sa21_sub[2];
  assign _0238_ = _0237_ ^ _0068_;
  assign _0239_ = _0238_ ^ w3[26];
  assign _0005_[2] = ld_r ? _0235_ : _0239_;
  assign _0240_ = w3[27] ^ text_in_r[27];
  assign _0241_ = _0188_ ^ _0064_;
  assign _0242_ = _0241_ ^ _0062_;
  assign _0243_ = _0242_ ^ sa21_sub[3];
  assign _0244_ = _0243_ ^ _0078_;
  assign _0245_ = _0244_ ^ w3[27];
  assign _0005_[3] = ld_r ? _0240_ : _0245_;
  assign _0246_ = w3[28] ^ text_in_r[28];
  assign _0247_ = ~w3[28];
  assign _0248_ = _0196_ ^ _0074_;
  assign _0249_ = _0248_ ^ sa10_sub[4];
  assign _0250_ = _0249_ ^ _0145_;
  assign _0251_ = _0250_ ^ sa32_sub[4];
  assign _0252_ = _0251_ ^ _0247_;
  assign _0005_[4] = ld_r ? _0246_ : _0252_;
  assign _0253_ = w3[29] ^ text_in_r[29];
  assign _0254_ = ~w3[29];
  assign _0255_ = _0137_ ^ _0084_;
  assign _0256_ = _0255_ ^ sa21_sub[5];
  assign _0257_ = _0256_ ^ sa32_sub[5];
  assign _0258_ = _0257_ ^ _0254_;
  assign _0005_[5] = ld_r ? _0253_ : _0258_;
  assign _0259_ = w3[30] ^ text_in_r[30];
  assign _0260_ = ~w3[30];
  assign _0261_ = _0146_ ^ _0092_;
  assign _0262_ = _0261_ ^ sa21_sub[6];
  assign _0263_ = _0262_ ^ sa32_sub[6];
  assign _0264_ = _0263_ ^ _0260_;
  assign _0005_[6] = ld_r ? _0259_ : _0264_;
  assign _0265_ = w3[31] ^ text_in_r[31];
  assign _0266_ = ~w3[31];
  assign _0267_ = _0154_ ^ _0100_;
  assign _0268_ = _0267_ ^ sa21_sub[7];
  assign _0269_ = _0268_ ^ sa32_sub[7];
  assign _0270_ = _0269_ ^ _0266_;
  assign _0005_[7] = ld_r ? _0265_ : _0270_;
  assign _0271_ = w2[0] ^ text_in_r[32];
  assign _0272_ = ~w2[0];
  assign _0273_ = ~sa12_sr[0];
  assign _0274_ = sa02_sr[7] ^ sa02_sr[0];
  assign _0275_ = _0274_ ^ _0273_;
  assign _0276_ = _0275_ ^ sa20_sub[0];
  assign _0277_ = _0276_ ^ sa31_sub[7];
  assign _0278_ = _0277_ ^ _0272_;
  assign _0016_[0] = ld_r ? _0271_ : _0278_;
  assign _0279_ = w2[1] ^ text_in_r[33];
  assign _0280_ = ~sa02_sr[1];
  assign _0281_ = _0274_ ^ _0280_;
  assign _0282_ = _0281_ ^ sa12_sr[1];
  assign _0283_ = _0282_ ^ sa20_sub[1];
  assign _0284_ = ~sa31_sub[0];
  assign _0285_ = sa31_sub[7] ^ _0284_;
  assign _0286_ = _0285_ ^ _0283_;
  assign _0287_ = _0286_ ^ w2[1];
  assign _0016_[1] = ld_r ? _0279_ : _0287_;
  assign _0288_ = w2[2] ^ text_in_r[34];
  assign _0289_ = ~w2[2];
  assign _0290_ = ~sa12_sr[2];
  assign _0291_ = sa02_sr[2] ^ sa02_sr[1];
  assign _0292_ = _0291_ ^ _0290_;
  assign _0293_ = _0292_ ^ sa20_sub[2];
  assign _0294_ = _0293_ ^ sa31_sub[1];
  assign _0295_ = _0294_ ^ _0289_;
  assign _0016_[2] = ld_r ? _0288_ : _0295_;
  assign _0296_ = w2[3] ^ text_in_r[35];
  assign _0297_ = ~w2[3];
  assign _0298_ = ~sa12_sr[3];
  assign _0299_ = ~sa02_sr[3];
  assign _0300_ = sa02_sr[7] ^ sa02_sr[2];
  assign _0301_ = _0300_ ^ _0299_;
  assign _0302_ = _0301_ ^ _0298_;
  assign _0303_ = _0302_ ^ sa20_sub[3];
  assign _0304_ = ~sa31_sub[2];
  assign _0305_ = sa31_sub[7] ^ _0304_;
  assign _0306_ = _0305_ ^ _0303_;
  assign _0307_ = _0306_ ^ _0297_;
  assign _0016_[3] = ld_r ? _0296_ : _0307_;
  assign _0308_ = w2[4] ^ text_in_r[36];
  assign _0309_ = ~sa02_sr[4];
  assign _0310_ = sa02_sr[7] ^ sa02_sr[3];
  assign _0311_ = _0310_ ^ _0309_;
  assign _0312_ = _0311_ ^ sa12_sr[4];
  assign _0313_ = _0312_ ^ sa20_sub[4];
  assign _0314_ = ~sa31_sub[3];
  assign _0315_ = sa31_sub[7] ^ _0314_;
  assign _0316_ = _0315_ ^ _0313_;
  assign _0317_ = _0316_ ^ w2[4];
  assign _0016_[4] = ld_r ? _0308_ : _0317_;
  assign _0318_ = w2[5] ^ text_in_r[37];
  assign _0319_ = ~w2[5];
  assign _0320_ = ~sa12_sr[5];
  assign _0321_ = sa02_sr[5] ^ sa02_sr[4];
  assign _0322_ = _0321_ ^ _0320_;
  assign _0323_ = _0322_ ^ sa20_sub[5];
  assign _0324_ = _0323_ ^ sa31_sub[4];
  assign _0325_ = _0324_ ^ _0319_;
  assign _0016_[5] = ld_r ? _0318_ : _0325_;
  assign _0326_ = w2[6] ^ text_in_r[38];
  assign _0327_ = ~w2[6];
  assign _0328_ = ~sa12_sr[6];
  assign _0329_ = sa02_sr[6] ^ sa02_sr[5];
  assign _0330_ = _0329_ ^ _0328_;
  assign _0331_ = _0330_ ^ sa20_sub[6];
  assign _0332_ = _0331_ ^ sa31_sub[5];
  assign _0333_ = _0332_ ^ _0327_;
  assign _0016_[6] = ld_r ? _0326_ : _0333_;
  assign _0334_ = w2[7] ^ text_in_r[39];
  assign _0335_ = ~w2[7];
  assign _0336_ = ~sa12_sr[7];
  assign _0337_ = sa02_sr[7] ^ sa02_sr[6];
  assign _0338_ = _0337_ ^ _0336_;
  assign _0339_ = _0338_ ^ sa20_sub[7];
  assign _0340_ = _0339_ ^ sa31_sub[6];
  assign _0341_ = _0340_ ^ _0335_;
  assign _0016_[7] = ld_r ? _0334_ : _0341_;
  assign _0342_ = w2[8] ^ text_in_r[40];
  assign _0343_ = ~sa20_sub[7];
  assign _0344_ = sa12_sr[0] ^ sa02_sr[0];
  assign _0345_ = _0344_ ^ _0343_;
  assign _0346_ = _0345_ ^ sa31_sub[7];
  assign _0347_ = _0346_ ^ _0284_;
  assign _0348_ = _0347_ ^ w2[8];
  assign _0012_[0] = ld_r ? _0342_ : _0348_;
  assign _0349_ = w2[9] ^ text_in_r[41];
  assign _0350_ = ~w2[9];
  assign _0351_ = sa12_sr[1] ^ sa02_sr[1];
  assign _0352_ = sa20_sub[7] ^ sa20_sub[0];
  assign _0353_ = _0352_ ^ _0351_;
  assign _0354_ = _0353_ ^ _0285_;
  assign _0355_ = _0354_ ^ sa31_sub[1];
  assign _0356_ = _0355_ ^ _0350_;
  assign _0012_[1] = ld_r ? _0349_ : _0356_;
  assign _0357_ = w2[10] ^ text_in_r[42];
  assign _0358_ = ~sa20_sub[1];
  assign _0359_ = sa12_sr[2] ^ sa02_sr[2];
  assign _0360_ = _0359_ ^ _0358_;
  assign _0361_ = _0360_ ^ sa31_sub[1];
  assign _0362_ = _0361_ ^ _0304_;
  assign _0363_ = _0362_ ^ w2[10];
  assign _0012_[2] = ld_r ? _0357_ : _0363_;
  assign _0364_ = w2[11] ^ text_in_r[43];
  assign _0365_ = sa12_sr[3] ^ sa02_sr[3];
  assign _0366_ = sa20_sub[7] ^ sa20_sub[2];
  assign _0367_ = _0366_ ^ _0365_;
  assign _0368_ = _0367_ ^ _0305_;
  assign _0369_ = _0368_ ^ _0314_;
  assign _0370_ = _0369_ ^ w2[11];
  assign _0012_[3] = ld_r ? _0364_ : _0370_;
  assign _0371_ = w2[12] ^ text_in_r[44];
  assign _0372_ = ~w2[12];
  assign _0373_ = sa12_sr[4] ^ sa02_sr[4];
  assign _0374_ = sa20_sub[7] ^ sa20_sub[3];
  assign _0375_ = _0374_ ^ _0373_;
  assign _0376_ = _0375_ ^ _0315_;
  assign _0377_ = _0376_ ^ sa31_sub[4];
  assign _0378_ = _0377_ ^ _0372_;
  assign _0012_[4] = ld_r ? _0371_ : _0378_;
  assign _0379_ = w2[13] ^ text_in_r[45];
  assign _0380_ = ~w2[13];
  assign _0381_ = ~sa20_sub[4];
  assign _0382_ = sa12_sr[5] ^ sa02_sr[5];
  assign _0383_ = _0382_ ^ _0381_;
  assign _0384_ = _0383_ ^ sa31_sub[4];
  assign _0385_ = _0384_ ^ sa31_sub[5];
  assign _0386_ = _0385_ ^ _0380_;
  assign _0012_[5] = ld_r ? _0379_ : _0386_;
  assign _0387_ = w2[14] ^ text_in_r[46];
  assign _0388_ = ~w2[14];
  assign _0389_ = ~sa20_sub[5];
  assign _0390_ = sa12_sr[6] ^ sa02_sr[6];
  assign _0391_ = _0390_ ^ _0389_;
  assign _0392_ = _0391_ ^ sa31_sub[5];
  assign _0393_ = _0392_ ^ sa31_sub[6];
  assign _0394_ = _0393_ ^ _0388_;
  assign _0012_[6] = ld_r ? _0387_ : _0394_;
  assign _0395_ = w2[15] ^ text_in_r[47];
  assign _0396_ = ~w2[15];
  assign _0397_ = ~sa20_sub[6];
  assign _0398_ = sa12_sr[7] ^ sa02_sr[7];
  assign _0399_ = _0398_ ^ _0397_;
  assign _0400_ = _0399_ ^ sa31_sub[6];
  assign _0401_ = _0400_ ^ sa31_sub[7];
  assign _0402_ = _0401_ ^ _0396_;
  assign _0012_[7] = ld_r ? _0395_ : _0402_;
  assign _0403_ = w2[16] ^ text_in_r[48];
  assign _0404_ = sa12_sr[7] ^ sa02_sr[0];
  assign _0405_ = _0404_ ^ _0343_;
  assign _0406_ = _0405_ ^ sa20_sub[0];
  assign _0407_ = _0406_ ^ _0284_;
  assign _0408_ = _0407_ ^ w2[16];
  assign _0008_[0] = ld_r ? _0403_ : _0408_;
  assign _0409_ = w2[17] ^ text_in_r[49];
  assign _0410_ = ~w2[17];
  assign _0411_ = sa12_sr[7] ^ sa12_sr[0];
  assign _0412_ = _0411_ ^ _0280_;
  assign _0413_ = _0412_ ^ _0352_;
  assign _0414_ = _0413_ ^ sa20_sub[1];
  assign _0415_ = _0414_ ^ sa31_sub[1];
  assign _0416_ = _0415_ ^ _0410_;
  assign _0008_[1] = ld_r ? _0409_ : _0416_;
  assign _0417_ = w2[18] ^ text_in_r[50];
  assign _0418_ = sa12_sr[1] ^ sa02_sr[2];
  assign _0419_ = _0418_ ^ _0358_;
  assign _0420_ = _0419_ ^ sa20_sub[2];
  assign _0421_ = _0420_ ^ _0304_;
  assign _0422_ = _0421_ ^ w2[18];
  assign _0008_[2] = ld_r ? _0417_ : _0422_;
  assign _0423_ = w2[19] ^ text_in_r[51];
  assign _0424_ = sa12_sr[7] ^ sa12_sr[2];
  assign _0425_ = _0424_ ^ _0299_;
  assign _0426_ = _0425_ ^ _0366_;
  assign _0427_ = _0426_ ^ sa20_sub[3];
  assign _0428_ = _0427_ ^ _0314_;
  assign _0429_ = _0428_ ^ w2[19];
  assign _0008_[3] = ld_r ? _0423_ : _0429_;
  assign _0430_ = w2[20] ^ text_in_r[52];
  assign _0431_ = ~w2[20];
  assign _0432_ = sa12_sr[7] ^ sa12_sr[3];
  assign _0433_ = _0432_ ^ _0309_;
  assign _0434_ = _0433_ ^ _0374_;
  assign _0435_ = _0434_ ^ sa20_sub[4];
  assign _0436_ = _0435_ ^ sa31_sub[4];
  assign _0437_ = _0436_ ^ _0431_;
  assign _0008_[4] = ld_r ? _0430_ : _0437_;
  assign _0438_ = w2[21] ^ text_in_r[53];
  assign _0439_ = ~w2[21];
  assign _0440_ = sa12_sr[4] ^ sa02_sr[5];
  assign _0441_ = _0440_ ^ _0381_;
  assign _0442_ = _0441_ ^ sa20_sub[5];
  assign _0443_ = _0442_ ^ sa31_sub[5];
  assign _0444_ = _0443_ ^ _0439_;
  assign _0008_[5] = ld_r ? _0438_ : _0444_;
  assign _0445_ = w2[22] ^ text_in_r[54];
  assign _0446_ = ~w2[22];
  assign _0447_ = sa12_sr[5] ^ sa02_sr[6];
  assign _0448_ = _0447_ ^ _0389_;
  assign _0449_ = _0448_ ^ sa20_sub[6];
  assign _0450_ = _0449_ ^ sa31_sub[6];
  assign _0451_ = _0450_ ^ _0446_;
  assign _0008_[6] = ld_r ? _0445_ : _0451_;
  assign _0452_ = w2[23] ^ text_in_r[55];
  assign _0453_ = ~w2[23];
  assign _0454_ = sa12_sr[6] ^ sa02_sr[7];
  assign _0455_ = _0454_ ^ _0397_;
  assign _0456_ = _0455_ ^ sa20_sub[7];
  assign _0457_ = _0456_ ^ sa31_sub[7];
  assign _0458_ = _0457_ ^ _0453_;
  assign _0008_[7] = ld_r ? _0452_ : _0458_;
  assign _0459_ = w2[24] ^ text_in_r[56];
  assign _0460_ = _0398_ ^ _0273_;
  assign _0461_ = _0460_ ^ sa20_sub[0];
  assign _0462_ = _0461_ ^ _0284_;
  assign _0463_ = _0462_ ^ w2[24];
  assign _0004_[0] = ld_r ? _0459_ : _0463_;
  assign _0464_ = w2[25] ^ text_in_r[57];
  assign _0465_ = ~w2[25];
  assign _0466_ = _0411_ ^ _0274_;
  assign _0467_ = _0466_ ^ sa12_sr[1];
  assign _0468_ = _0467_ ^ _0358_;
  assign _0469_ = _0468_ ^ sa31_sub[1];
  assign _0470_ = _0469_ ^ _0465_;
  assign _0004_[1] = ld_r ? _0464_ : _0470_;
  assign _0471_ = w2[26] ^ text_in_r[58];
  assign _0472_ = _0351_ ^ _0290_;
  assign _0473_ = _0472_ ^ sa20_sub[2];
  assign _0474_ = _0473_ ^ _0304_;
  assign _0475_ = _0474_ ^ w2[26];
  assign _0004_[2] = ld_r ? _0471_ : _0475_;
  assign _0476_ = w2[27] ^ text_in_r[59];
  assign _0477_ = _0424_ ^ _0300_;
  assign _0478_ = _0477_ ^ _0298_;
  assign _0479_ = _0478_ ^ sa20_sub[3];
  assign _0480_ = _0479_ ^ _0314_;
  assign _0481_ = _0480_ ^ w2[27];
  assign _0004_[3] = ld_r ? _0476_ : _0481_;
  assign _0482_ = w2[28] ^ text_in_r[60];
  assign _0483_ = ~w2[28];
  assign _0484_ = _0432_ ^ _0310_;
  assign _0485_ = _0484_ ^ sa12_sr[4];
  assign _0486_ = _0485_ ^ _0381_;
  assign _0487_ = _0486_ ^ sa31_sub[4];
  assign _0488_ = _0487_ ^ _0483_;
  assign _0004_[4] = ld_r ? _0482_ : _0488_;
  assign _0489_ = w2[29] ^ text_in_r[61];
  assign _0490_ = ~w2[29];
  assign _0491_ = _0373_ ^ _0320_;
  assign _0492_ = _0491_ ^ sa20_sub[5];
  assign _0493_ = _0492_ ^ sa31_sub[5];
  assign _0494_ = _0493_ ^ _0490_;
  assign _0004_[5] = ld_r ? _0489_ : _0494_;
  assign _0495_ = w2[30] ^ text_in_r[62];
  assign _0496_ = ~w2[30];
  assign _0497_ = _0382_ ^ _0328_;
  assign _0498_ = _0497_ ^ sa20_sub[6];
  assign _0499_ = _0498_ ^ sa31_sub[6];
  assign _0500_ = _0499_ ^ _0496_;
  assign _0004_[6] = ld_r ? _0495_ : _0500_;
  assign _0501_ = w2[31] ^ text_in_r[63];
  assign _0502_ = ~w2[31];
  assign _0503_ = _0390_ ^ _0336_;
  assign _0504_ = _0503_ ^ sa20_sub[7];
  assign _0505_ = _0504_ ^ sa31_sub[7];
  assign _0506_ = _0505_ ^ _0502_;
  assign _0004_[7] = ld_r ? _0501_ : _0506_;
  assign _0507_ = w1[0] ^ text_in_r[64];
  assign _0508_ = ~w1[0];
  assign _0509_ = ~sa11_sr[0];
  assign _0510_ = sa01_sr[7] ^ sa01_sr[0];
  assign _0511_ = _0510_ ^ _0509_;
  assign _0512_ = _0511_ ^ sa21_sr[0];
  assign _0513_ = _0512_ ^ sa30_sub[7];
  assign _0514_ = _0513_ ^ _0508_;
  assign _0015_[0] = ld_r ? _0507_ : _0514_;
  assign _0515_ = w1[1] ^ text_in_r[65];
  assign _0516_ = ~sa01_sr[1];
  assign _0517_ = _0510_ ^ _0516_;
  assign _0518_ = _0517_ ^ sa11_sr[1];
  assign _0519_ = _0518_ ^ sa21_sr[1];
  assign _0520_ = ~sa30_sub[0];
  assign _0521_ = sa30_sub[7] ^ _0520_;
  assign _0522_ = _0521_ ^ _0519_;
  assign _0523_ = _0522_ ^ w1[1];
  assign _0015_[1] = ld_r ? _0515_ : _0523_;
  assign _0524_ = w1[2] ^ text_in_r[66];
  assign _0525_ = ~w1[2];
  assign _0526_ = ~sa11_sr[2];
  assign _0527_ = sa01_sr[2] ^ sa01_sr[1];
  assign _0528_ = _0527_ ^ _0526_;
  assign _0529_ = _0528_ ^ sa21_sr[2];
  assign _0530_ = _0529_ ^ sa30_sub[1];
  assign _0531_ = _0530_ ^ _0525_;
  assign _0015_[2] = ld_r ? _0524_ : _0531_;
  assign _0532_ = w1[3] ^ text_in_r[67];
  assign _0533_ = ~w1[3];
  assign _0534_ = ~sa11_sr[3];
  assign _0535_ = ~sa01_sr[3];
  assign _0536_ = sa01_sr[7] ^ sa01_sr[2];
  assign _0537_ = _0536_ ^ _0535_;
  assign _0538_ = _0537_ ^ _0534_;
  assign _0539_ = _0538_ ^ sa21_sr[3];
  assign _0540_ = ~sa30_sub[2];
  assign _0541_ = sa30_sub[7] ^ _0540_;
  assign _0542_ = _0541_ ^ _0539_;
  assign _0543_ = _0542_ ^ _0533_;
  assign _0015_[3] = ld_r ? _0532_ : _0543_;
  assign _0544_ = w1[4] ^ text_in_r[68];
  assign _0545_ = ~sa01_sr[4];
  assign _0546_ = sa01_sr[7] ^ sa01_sr[3];
  assign _0547_ = _0546_ ^ _0545_;
  assign _0548_ = _0547_ ^ sa11_sr[4];
  assign _0549_ = _0548_ ^ sa21_sr[4];
  assign _0550_ = ~sa30_sub[3];
  assign _0551_ = sa30_sub[7] ^ _0550_;
  assign _0552_ = _0551_ ^ _0549_;
  assign _0553_ = _0552_ ^ w1[4];
  assign _0015_[4] = ld_r ? _0544_ : _0553_;
  assign _0554_ = w1[5] ^ text_in_r[69];
  assign _0555_ = ~w1[5];
  assign _0556_ = ~sa11_sr[5];
  assign _0557_ = sa01_sr[5] ^ sa01_sr[4];
  assign _0558_ = _0557_ ^ _0556_;
  assign _0559_ = _0558_ ^ sa21_sr[5];
  assign _0560_ = _0559_ ^ sa30_sub[4];
  assign _0561_ = _0560_ ^ _0555_;
  assign _0015_[5] = ld_r ? _0554_ : _0561_;
  assign _0562_ = w1[6] ^ text_in_r[70];
  assign _0563_ = ~w1[6];
  assign _0564_ = ~sa11_sr[6];
  assign _0565_ = sa01_sr[6] ^ sa01_sr[5];
  assign _0566_ = _0565_ ^ _0564_;
  assign _0567_ = _0566_ ^ sa21_sr[6];
  assign _0568_ = _0567_ ^ sa30_sub[5];
  assign _0569_ = _0568_ ^ _0563_;
  assign _0015_[6] = ld_r ? _0562_ : _0569_;
  assign _0570_ = w1[7] ^ text_in_r[71];
  assign _0571_ = ~w1[7];
  assign _0572_ = ~sa11_sr[7];
  assign _0573_ = sa01_sr[7] ^ sa01_sr[6];
  assign _0574_ = _0573_ ^ _0572_;
  assign _0575_ = _0574_ ^ sa21_sr[7];
  assign _0576_ = _0575_ ^ sa30_sub[6];
  assign _0577_ = _0576_ ^ _0571_;
  assign _0015_[7] = ld_r ? _0570_ : _0577_;
  assign _0578_ = w1[8] ^ text_in_r[72];
  assign _0579_ = ~sa21_sr[7];
  assign _0580_ = sa11_sr[0] ^ sa01_sr[0];
  assign _0581_ = _0580_ ^ _0579_;
  assign _0582_ = _0581_ ^ sa30_sub[7];
  assign _0583_ = _0582_ ^ _0520_;
  assign _0584_ = _0583_ ^ w1[8];
  assign _0011_[0] = ld_r ? _0578_ : _0584_;
  assign _0585_ = w1[9] ^ text_in_r[73];
  assign _0586_ = ~w1[9];
  assign _0587_ = sa11_sr[1] ^ sa01_sr[1];
  assign _0588_ = sa21_sr[7] ^ sa21_sr[0];
  assign _0589_ = _0588_ ^ _0587_;
  assign _0590_ = _0589_ ^ _0521_;
  assign _0591_ = _0590_ ^ sa30_sub[1];
  assign _0592_ = _0591_ ^ _0586_;
  assign _0011_[1] = ld_r ? _0585_ : _0592_;
  assign _0593_ = w1[10] ^ text_in_r[74];
  assign _0594_ = ~sa21_sr[1];
  assign _0595_ = sa11_sr[2] ^ sa01_sr[2];
  assign _0596_ = _0595_ ^ _0594_;
  assign _0597_ = _0596_ ^ sa30_sub[1];
  assign _0598_ = _0597_ ^ _0540_;
  assign _0599_ = _0598_ ^ w1[10];
  assign _0011_[2] = ld_r ? _0593_ : _0599_;
  assign _0600_ = w1[11] ^ text_in_r[75];
  assign _0601_ = sa11_sr[3] ^ sa01_sr[3];
  assign _0602_ = sa21_sr[7] ^ sa21_sr[2];
  assign _0603_ = _0602_ ^ _0601_;
  assign _0604_ = _0603_ ^ _0541_;
  assign _0605_ = _0604_ ^ _0550_;
  assign _0606_ = _0605_ ^ w1[11];
  assign _0011_[3] = ld_r ? _0600_ : _0606_;
  assign _0607_ = w1[12] ^ text_in_r[76];
  assign _0608_ = ~w1[12];
  assign _0609_ = sa11_sr[4] ^ sa01_sr[4];
  assign _0610_ = sa21_sr[7] ^ sa21_sr[3];
  assign _0611_ = _0610_ ^ _0609_;
  assign _0612_ = _0611_ ^ _0551_;
  assign _0613_ = _0612_ ^ sa30_sub[4];
  assign _0614_ = _0613_ ^ _0608_;
  assign _0011_[4] = ld_r ? _0607_ : _0614_;
  assign _0615_ = w1[13] ^ text_in_r[77];
  assign _0616_ = ~w1[13];
  assign _0617_ = ~sa21_sr[4];
  assign _0618_ = sa11_sr[5] ^ sa01_sr[5];
  assign _0619_ = _0618_ ^ _0617_;
  assign _0620_ = _0619_ ^ sa30_sub[4];
  assign _0621_ = _0620_ ^ sa30_sub[5];
  assign _0622_ = _0621_ ^ _0616_;
  assign _0011_[5] = ld_r ? _0615_ : _0622_;
  assign _0623_ = w1[14] ^ text_in_r[78];
  assign _0624_ = ~w1[14];
  assign _0625_ = ~sa21_sr[5];
  assign _0626_ = sa11_sr[6] ^ sa01_sr[6];
  assign _0627_ = _0626_ ^ _0625_;
  assign _0628_ = _0627_ ^ sa30_sub[5];
  assign _0629_ = _0628_ ^ sa30_sub[6];
  assign _0630_ = _0629_ ^ _0624_;
  assign _0011_[6] = ld_r ? _0623_ : _0630_;
  assign _0631_ = w1[15] ^ text_in_r[79];
  assign _0632_ = ~w1[15];
  assign _0633_ = ~sa21_sr[6];
  assign _0634_ = sa11_sr[7] ^ sa01_sr[7];
  assign _0635_ = _0634_ ^ _0633_;
  assign _0636_ = _0635_ ^ sa30_sub[6];
  assign _0637_ = _0636_ ^ sa30_sub[7];
  assign _0638_ = _0637_ ^ _0632_;
  assign _0011_[7] = ld_r ? _0631_ : _0638_;
  assign _0639_ = w1[16] ^ text_in_r[80];
  assign _0640_ = sa11_sr[7] ^ sa01_sr[0];
  assign _0641_ = _0640_ ^ _0579_;
  assign _0642_ = _0641_ ^ sa21_sr[0];
  assign _0643_ = _0642_ ^ _0520_;
  assign _0644_ = _0643_ ^ w1[16];
  assign _0007_[0] = ld_r ? _0639_ : _0644_;
  assign _0645_ = w1[17] ^ text_in_r[81];
  assign _0646_ = ~w1[17];
  assign _0647_ = sa11_sr[7] ^ sa11_sr[0];
  assign _0648_ = _0647_ ^ _0516_;
  assign _0649_ = _0648_ ^ _0588_;
  assign _0650_ = _0649_ ^ sa21_sr[1];
  assign _0651_ = _0650_ ^ sa30_sub[1];
  assign _0652_ = _0651_ ^ _0646_;
  assign _0007_[1] = ld_r ? _0645_ : _0652_;
  assign _0653_ = w1[18] ^ text_in_r[82];
  assign _0654_ = sa11_sr[1] ^ sa01_sr[2];
  assign _0655_ = _0654_ ^ _0594_;
  assign _0656_ = _0655_ ^ sa21_sr[2];
  assign _0657_ = _0656_ ^ _0540_;
  assign _0658_ = _0657_ ^ w1[18];
  assign _0007_[2] = ld_r ? _0653_ : _0658_;
  assign _0659_ = w1[19] ^ text_in_r[83];
  assign _0660_ = sa11_sr[7] ^ sa11_sr[2];
  assign _0661_ = _0660_ ^ _0535_;
  assign _0662_ = _0661_ ^ _0602_;
  assign _0663_ = _0662_ ^ sa21_sr[3];
  assign _0664_ = _0663_ ^ _0550_;
  assign _0665_ = _0664_ ^ w1[19];
  assign _0007_[3] = ld_r ? _0659_ : _0665_;
  assign _0666_ = w1[20] ^ text_in_r[84];
  assign _0667_ = ~w1[20];
  assign _0668_ = sa11_sr[7] ^ sa11_sr[3];
  assign _0669_ = _0668_ ^ _0545_;
  assign _0670_ = _0669_ ^ _0610_;
  assign _0671_ = _0670_ ^ sa21_sr[4];
  assign _0672_ = _0671_ ^ sa30_sub[4];
  assign _0673_ = _0672_ ^ _0667_;
  assign _0007_[4] = ld_r ? _0666_ : _0673_;
  assign _0674_ = w1[21] ^ text_in_r[85];
  assign _0675_ = ~w1[21];
  assign _0676_ = sa11_sr[4] ^ sa01_sr[5];
  assign _0677_ = _0676_ ^ _0617_;
  assign _0678_ = _0677_ ^ sa21_sr[5];
  assign _0679_ = _0678_ ^ sa30_sub[5];
  assign _0680_ = _0679_ ^ _0675_;
  assign _0007_[5] = ld_r ? _0674_ : _0680_;
  assign _0681_ = w1[22] ^ text_in_r[86];
  assign _0682_ = ~w1[22];
  assign _0683_ = sa11_sr[5] ^ sa01_sr[6];
  assign _0684_ = _0683_ ^ _0625_;
  assign _0685_ = _0684_ ^ sa21_sr[6];
  assign _0686_ = _0685_ ^ sa30_sub[6];
  assign _0687_ = _0686_ ^ _0682_;
  assign _0007_[6] = ld_r ? _0681_ : _0687_;
  assign _0688_ = w1[23] ^ text_in_r[87];
  assign _0689_ = ~w1[23];
  assign _0690_ = sa11_sr[6] ^ sa01_sr[7];
  assign _0691_ = _0690_ ^ _0633_;
  assign _0692_ = _0691_ ^ sa21_sr[7];
  assign _0693_ = _0692_ ^ sa30_sub[7];
  assign _0694_ = _0693_ ^ _0689_;
  assign _0007_[7] = ld_r ? _0688_ : _0694_;
  assign _0695_ = w1[24] ^ text_in_r[88];
  assign _0696_ = _0634_ ^ _0509_;
  assign _0697_ = _0696_ ^ sa21_sr[0];
  assign _0698_ = _0697_ ^ _0520_;
  assign _0699_ = _0698_ ^ w1[24];
  assign _0003_[0] = ld_r ? _0695_ : _0699_;
  assign _0700_ = w1[25] ^ text_in_r[89];
  assign _0701_ = ~w1[25];
  assign _0702_ = _0647_ ^ _0510_;
  assign _0703_ = _0702_ ^ sa11_sr[1];
  assign _0704_ = _0703_ ^ _0594_;
  assign _0705_ = _0704_ ^ sa30_sub[1];
  assign _0706_ = _0705_ ^ _0701_;
  assign _0003_[1] = ld_r ? _0700_ : _0706_;
  assign _0707_ = w1[26] ^ text_in_r[90];
  assign _0708_ = _0587_ ^ _0526_;
  assign _0709_ = _0708_ ^ sa21_sr[2];
  assign _0710_ = _0709_ ^ _0540_;
  assign _0711_ = _0710_ ^ w1[26];
  assign _0003_[2] = ld_r ? _0707_ : _0711_;
  assign _0712_ = w1[27] ^ text_in_r[91];
  assign _0713_ = _0660_ ^ _0536_;
  assign _0714_ = _0713_ ^ _0534_;
  assign _0715_ = _0714_ ^ sa21_sr[3];
  assign _0716_ = _0715_ ^ _0550_;
  assign _0717_ = _0716_ ^ w1[27];
  assign _0003_[3] = ld_r ? _0712_ : _0717_;
  assign _0718_ = w1[28] ^ text_in_r[92];
  assign _0719_ = ~w1[28];
  assign _0720_ = _0668_ ^ _0546_;
  assign _0721_ = _0720_ ^ sa11_sr[4];
  assign _0722_ = _0721_ ^ _0617_;
  assign _0723_ = _0722_ ^ sa30_sub[4];
  assign _0724_ = _0723_ ^ _0719_;
  assign _0003_[4] = ld_r ? _0718_ : _0724_;
  assign _0725_ = w1[29] ^ text_in_r[93];
  assign _0726_ = ~w1[29];
  assign _0727_ = _0609_ ^ _0556_;
  assign _0728_ = _0727_ ^ sa21_sr[5];
  assign _0729_ = _0728_ ^ sa30_sub[5];
  assign _0730_ = _0729_ ^ _0726_;
  assign _0003_[5] = ld_r ? _0725_ : _0730_;
  assign _0731_ = w1[30] ^ text_in_r[94];
  assign _0732_ = ~w1[30];
  assign _0733_ = _0618_ ^ _0564_;
  assign _0734_ = _0733_ ^ sa21_sr[6];
  assign _0735_ = _0734_ ^ sa30_sub[6];
  assign _0736_ = _0735_ ^ _0732_;
  assign _0003_[6] = ld_r ? _0731_ : _0736_;
  assign _0737_ = w1[31] ^ text_in_r[95];
  assign _0738_ = ~w1[31];
  assign _0739_ = _0626_ ^ _0572_;
  assign _0740_ = _0739_ ^ sa21_sr[7];
  assign _0741_ = _0740_ ^ sa30_sub[7];
  assign _0742_ = _0741_ ^ _0738_;
  assign _0003_[7] = ld_r ? _0737_ : _0742_;
  assign _0743_ = w0[0] ^ text_in_r[96];
  assign _0744_ = ~w0[0];
  assign _0745_ = ~sa10_sr[0];
  assign _0746_ = sa00_sr[7] ^ sa00_sr[0];
  assign _0747_ = _0746_ ^ _0745_;
  assign _0748_ = _0747_ ^ sa20_sr[0];
  assign _0749_ = _0748_ ^ sa30_sr[7];
  assign _0750_ = _0749_ ^ _0744_;
  assign _0014_[0] = ld_r ? _0743_ : _0750_;
  assign _0751_ = w0[1] ^ text_in_r[97];
  assign _0752_ = ~sa00_sr[1];
  assign _0753_ = _0746_ ^ _0752_;
  assign _0754_ = _0753_ ^ sa10_sr[1];
  assign _0755_ = _0754_ ^ sa20_sr[1];
  assign _0756_ = ~sa30_sr[0];
  assign _0757_ = sa30_sr[7] ^ _0756_;
  assign _0758_ = _0757_ ^ _0755_;
  assign _0759_ = _0758_ ^ w0[1];
  assign _0014_[1] = ld_r ? _0751_ : _0759_;
  assign _0760_ = w0[2] ^ text_in_r[98];
  assign _0761_ = ~w0[2];
  assign _0762_ = ~sa10_sr[2];
  assign _0763_ = sa00_sr[2] ^ sa00_sr[1];
  assign _0764_ = _0763_ ^ _0762_;
  assign _0765_ = _0764_ ^ sa20_sr[2];
  assign _0766_ = _0765_ ^ sa30_sr[1];
  assign _0767_ = _0766_ ^ _0761_;
  assign _0014_[2] = ld_r ? _0760_ : _0767_;
  assign _0768_ = w0[3] ^ text_in_r[99];
  assign _0769_ = ~w0[3];
  assign _0770_ = ~sa10_sr[3];
  assign _0771_ = ~sa00_sr[3];
  assign _0772_ = sa00_sr[7] ^ sa00_sr[2];
  assign _0773_ = _0772_ ^ _0771_;
  assign _0774_ = _0773_ ^ _0770_;
  assign _0775_ = _0774_ ^ sa20_sr[3];
  assign _0776_ = ~sa30_sr[2];
  assign _0777_ = sa30_sr[7] ^ _0776_;
  assign _0778_ = _0777_ ^ _0775_;
  assign _0779_ = _0778_ ^ _0769_;
  assign _0014_[3] = ld_r ? _0768_ : _0779_;
  assign _0780_ = w0[4] ^ text_in_r[100];
  assign _0781_ = ~sa00_sr[4];
  assign _0782_ = sa00_sr[7] ^ sa00_sr[3];
  assign _0783_ = _0782_ ^ _0781_;
  assign _0784_ = _0783_ ^ sa10_sr[4];
  assign _0785_ = _0784_ ^ sa20_sr[4];
  assign _0786_ = ~sa30_sr[3];
  assign _0787_ = sa30_sr[7] ^ _0786_;
  assign _0788_ = _0787_ ^ _0785_;
  assign _0789_ = _0788_ ^ w0[4];
  assign _0014_[4] = ld_r ? _0780_ : _0789_;
  assign _0790_ = w0[5] ^ text_in_r[101];
  assign _0791_ = ~w0[5];
  assign _0792_ = ~sa10_sr[5];
  assign _0793_ = sa00_sr[5] ^ sa00_sr[4];
  assign _0794_ = _0793_ ^ _0792_;
  assign _0795_ = _0794_ ^ sa20_sr[5];
  assign _0796_ = _0795_ ^ sa30_sr[4];
  assign _0797_ = _0796_ ^ _0791_;
  assign _0014_[5] = ld_r ? _0790_ : _0797_;
  assign _0798_ = w0[6] ^ text_in_r[102];
  assign _0799_ = ~w0[6];
  assign _0800_ = ~sa10_sr[6];
  assign _0801_ = sa00_sr[6] ^ sa00_sr[5];
  assign _0802_ = _0801_ ^ _0800_;
  assign _0803_ = _0802_ ^ sa20_sr[6];
  assign _0804_ = _0803_ ^ sa30_sr[5];
  assign _0805_ = _0804_ ^ _0799_;
  assign _0014_[6] = ld_r ? _0798_ : _0805_;
  assign _0806_ = w0[7] ^ text_in_r[103];
  assign _0807_ = ~w0[7];
  assign _0808_ = ~sa10_sr[7];
  assign _0809_ = sa00_sr[7] ^ sa00_sr[6];
  assign _0810_ = _0809_ ^ _0808_;
  assign _0811_ = _0810_ ^ sa20_sr[7];
  assign _0812_ = _0811_ ^ sa30_sr[6];
  assign _0813_ = _0812_ ^ _0807_;
  assign _0014_[7] = ld_r ? _0806_ : _0813_;
  assign _0814_ = w0[8] ^ text_in_r[104];
  assign _0815_ = ~sa20_sr[7];
  assign _0816_ = sa10_sr[0] ^ sa00_sr[0];
  assign _0817_ = _0816_ ^ _0815_;
  assign _0818_ = _0817_ ^ sa30_sr[7];
  assign _0819_ = _0818_ ^ _0756_;
  assign _0820_ = _0819_ ^ w0[8];
  assign _0010_[0] = ld_r ? _0814_ : _0820_;
  assign _0821_ = w0[9] ^ text_in_r[105];
  assign _0822_ = ~w0[9];
  assign _0823_ = sa10_sr[1] ^ sa00_sr[1];
  assign _0824_ = sa20_sr[7] ^ sa20_sr[0];
  assign _0825_ = _0824_ ^ _0823_;
  assign _0826_ = _0825_ ^ _0757_;
  assign _0827_ = _0826_ ^ sa30_sr[1];
  assign _0828_ = _0827_ ^ _0822_;
  assign _0010_[1] = ld_r ? _0821_ : _0828_;
  assign _0829_ = w0[10] ^ text_in_r[106];
  assign _0830_ = ~sa20_sr[1];
  assign _0831_ = sa10_sr[2] ^ sa00_sr[2];
  assign _0832_ = _0831_ ^ _0830_;
  assign _0833_ = _0832_ ^ sa30_sr[1];
  assign _0834_ = _0833_ ^ _0776_;
  assign _0835_ = _0834_ ^ w0[10];
  assign _0010_[2] = ld_r ? _0829_ : _0835_;
  assign _0836_ = w0[11] ^ text_in_r[107];
  assign _0837_ = sa10_sr[3] ^ sa00_sr[3];
  assign _0838_ = sa20_sr[7] ^ sa20_sr[2];
  assign _0839_ = _0838_ ^ _0837_;
  assign _0840_ = _0839_ ^ _0777_;
  assign _0841_ = _0840_ ^ _0786_;
  assign _0842_ = _0841_ ^ w0[11];
  assign _0010_[3] = ld_r ? _0836_ : _0842_;
  assign _0843_ = w0[12] ^ text_in_r[108];
  assign _0844_ = ~w0[12];
  assign _0845_ = sa10_sr[4] ^ sa00_sr[4];
  assign _0846_ = sa20_sr[7] ^ sa20_sr[3];
  assign _0847_ = _0846_ ^ _0845_;
  assign _0848_ = _0847_ ^ _0787_;
  assign _0849_ = _0848_ ^ sa30_sr[4];
  assign _0850_ = _0849_ ^ _0844_;
  assign _0010_[4] = ld_r ? _0843_ : _0850_;
  assign _0851_ = w0[13] ^ text_in_r[109];
  assign _0852_ = ~w0[13];
  assign _0853_ = ~sa20_sr[4];
  assign _0854_ = sa10_sr[5] ^ sa00_sr[5];
  assign _0855_ = _0854_ ^ _0853_;
  assign _0856_ = _0855_ ^ sa30_sr[4];
  assign _0857_ = _0856_ ^ sa30_sr[5];
  assign _0858_ = _0857_ ^ _0852_;
  assign _0010_[5] = ld_r ? _0851_ : _0858_;
  assign _0859_ = w0[14] ^ text_in_r[110];
  assign _0860_ = ~w0[14];
  assign _0861_ = ~sa20_sr[5];
  assign _0862_ = sa10_sr[6] ^ sa00_sr[6];
  assign _0863_ = _0862_ ^ _0861_;
  assign _0864_ = _0863_ ^ sa30_sr[5];
  assign _0865_ = _0864_ ^ sa30_sr[6];
  assign _0866_ = _0865_ ^ _0860_;
  assign _0010_[6] = ld_r ? _0859_ : _0866_;
  assign _0867_ = w0[15] ^ text_in_r[111];
  assign _0868_ = ~w0[15];
  assign _0869_ = ~sa20_sr[6];
  assign _0870_ = sa10_sr[7] ^ sa00_sr[7];
  assign _0871_ = _0870_ ^ _0869_;
  assign _0872_ = _0871_ ^ sa30_sr[6];
  assign _0873_ = _0872_ ^ sa30_sr[7];
  assign _0874_ = _0873_ ^ _0868_;
  assign _0010_[7] = ld_r ? _0867_ : _0874_;
  assign _0875_ = w0[16] ^ text_in_r[112];
  assign _0876_ = sa10_sr[7] ^ sa00_sr[0];
  assign _0877_ = _0876_ ^ _0815_;
  assign _0878_ = _0877_ ^ sa20_sr[0];
  assign _0879_ = _0878_ ^ _0756_;
  assign _0880_ = _0879_ ^ w0[16];
  assign _0006_[0] = ld_r ? _0875_ : _0880_;
  assign _0881_ = w0[17] ^ text_in_r[113];
  assign _0882_ = ~w0[17];
  assign _0883_ = sa10_sr[7] ^ sa10_sr[0];
  assign _0884_ = _0883_ ^ _0752_;
  assign _0885_ = _0884_ ^ _0824_;
  assign _0886_ = _0885_ ^ sa20_sr[1];
  assign _0887_ = _0886_ ^ sa30_sr[1];
  assign _0888_ = _0887_ ^ _0882_;
  assign _0006_[1] = ld_r ? _0881_ : _0888_;
  assign _0889_ = w0[18] ^ text_in_r[114];
  assign _0890_ = sa10_sr[1] ^ sa00_sr[2];
  assign _0891_ = _0890_ ^ _0830_;
  assign _0892_ = _0891_ ^ sa20_sr[2];
  assign _0893_ = _0892_ ^ _0776_;
  assign _0894_ = _0893_ ^ w0[18];
  assign _0006_[2] = ld_r ? _0889_ : _0894_;
  assign _0895_ = w0[19] ^ text_in_r[115];
  assign _0896_ = sa10_sr[7] ^ sa10_sr[2];
  assign _0897_ = _0896_ ^ _0771_;
  assign _0898_ = _0897_ ^ _0838_;
  assign _0899_ = _0898_ ^ sa20_sr[3];
  assign _0900_ = _0899_ ^ _0786_;
  assign _0901_ = _0900_ ^ w0[19];
  assign _0006_[3] = ld_r ? _0895_ : _0901_;
  assign _0902_ = w0[20] ^ text_in_r[116];
  assign _0903_ = ~w0[20];
  assign _0904_ = sa10_sr[7] ^ sa10_sr[3];
  assign _0905_ = _0904_ ^ _0781_;
  assign _0906_ = _0905_ ^ _0846_;
  assign _0907_ = _0906_ ^ sa20_sr[4];
  assign _0908_ = _0907_ ^ sa30_sr[4];
  assign _0909_ = _0908_ ^ _0903_;
  assign _0006_[4] = ld_r ? _0902_ : _0909_;
  assign _0910_ = w0[21] ^ text_in_r[117];
  assign _0911_ = ~w0[21];
  assign _0912_ = sa10_sr[4] ^ sa00_sr[5];
  assign _0913_ = _0912_ ^ _0853_;
  assign _0914_ = _0913_ ^ sa20_sr[5];
  assign _0915_ = _0914_ ^ sa30_sr[5];
  assign _0916_ = _0915_ ^ _0911_;
  assign _0006_[5] = ld_r ? _0910_ : _0916_;
  assign _0917_ = w0[22] ^ text_in_r[118];
  assign _0918_ = ~w0[22];
  assign _0919_ = sa10_sr[5] ^ sa00_sr[6];
  assign _0920_ = _0919_ ^ _0861_;
  assign _0921_ = _0920_ ^ sa20_sr[6];
  assign _0922_ = _0921_ ^ sa30_sr[6];
  assign _0923_ = _0922_ ^ _0918_;
  assign _0006_[6] = ld_r ? _0917_ : _0923_;
  assign _0924_ = w0[23] ^ text_in_r[119];
  assign _0925_ = ~w0[23];
  assign _0926_ = sa10_sr[6] ^ sa00_sr[7];
  assign _0927_ = _0926_ ^ _0869_;
  assign _0928_ = _0927_ ^ sa20_sr[7];
  assign _0929_ = _0928_ ^ sa30_sr[7];
  assign _0930_ = _0929_ ^ _0925_;
  assign _0006_[7] = ld_r ? _0924_ : _0930_;
  assign _0931_ = w0[24] ^ text_in_r[120];
  assign _0932_ = _0870_ ^ _0745_;
  assign _0933_ = _0932_ ^ sa20_sr[0];
  assign _0934_ = _0933_ ^ _0756_;
  assign _0935_ = _0934_ ^ w0[24];
  assign _0002_[0] = ld_r ? _0931_ : _0935_;
  assign _0936_ = w0[25] ^ text_in_r[121];
  assign _0937_ = ~w0[25];
  assign _0938_ = _0883_ ^ _0746_;
  assign _0939_ = _0938_ ^ sa10_sr[1];
  assign _0940_ = _0939_ ^ _0830_;
  assign _0941_ = _0940_ ^ sa30_sr[1];
  assign _0942_ = _0941_ ^ _0937_;
  assign _0002_[1] = ld_r ? _0936_ : _0942_;
  assign _0943_ = w0[26] ^ text_in_r[122];
  assign _0944_ = _0823_ ^ _0762_;
  assign _0945_ = _0944_ ^ sa20_sr[2];
  assign _0946_ = _0945_ ^ _0776_;
  assign _0947_ = _0946_ ^ w0[26];
  assign _0002_[2] = ld_r ? _0943_ : _0947_;
  assign _0948_ = w0[27] ^ text_in_r[123];
  assign _0949_ = _0896_ ^ _0772_;
  assign _0950_ = _0949_ ^ _0770_;
  assign _0951_ = _0950_ ^ sa20_sr[3];
  assign _0952_ = _0951_ ^ _0786_;
  assign _0953_ = _0952_ ^ w0[27];
  assign _0002_[3] = ld_r ? _0948_ : _0953_;
  assign _0954_ = w0[28] ^ text_in_r[124];
  assign _0955_ = ~w0[28];
  assign _0956_ = _0904_ ^ _0782_;
  assign _0957_ = _0956_ ^ sa10_sr[4];
  assign _0958_ = _0957_ ^ _0853_;
  assign _0959_ = _0958_ ^ sa30_sr[4];
  assign _0960_ = _0959_ ^ _0955_;
  assign _0002_[4] = ld_r ? _0954_ : _0960_;
  assign _0961_ = w0[29] ^ text_in_r[125];
  assign _0962_ = ~w0[29];
  assign _0963_ = _0845_ ^ _0792_;
  assign _0964_ = _0963_ ^ sa20_sr[5];
  assign _0965_ = _0964_ ^ sa30_sr[5];
  assign _0966_ = _0965_ ^ _0962_;
  assign _0002_[5] = ld_r ? _0961_ : _0966_;
  assign _0967_ = w0[30] ^ text_in_r[126];
  assign _0968_ = ~w0[30];
  assign _0969_ = _0854_ ^ _0800_;
  assign _0970_ = _0969_ ^ sa20_sr[6];
  assign _0971_ = _0970_ ^ sa30_sr[6];
  assign _0972_ = _0971_ ^ _0968_;
  assign _0002_[6] = ld_r ? _0967_ : _0972_;
  assign _0973_ = w0[31] ^ text_in_r[127];
  assign _0974_ = ~w0[31];
  assign _0975_ = _0862_ ^ _0808_;
  assign _0976_ = _0975_ ^ sa20_sr[7];
  assign _0977_ = _0976_ ^ sa30_sr[7];
  assign _0978_ = _0977_ ^ _0974_;
  assign _0002_[7] = ld_r ? _0973_ : _0978_;
  assign _0022_[0] = sa00_sr[0] ^ w0[24];
  assign _0022_[1] = sa00_sr[1] ^ w0[25];
  assign _0022_[2] = sa00_sr[2] ^ w0[26];
  assign _0022_[3] = sa00_sr[3] ^ w0[27];
  assign _0022_[4] = sa00_sr[4] ^ w0[28];
  assign _0022_[5] = sa00_sr[5] ^ w0[29];
  assign _0022_[6] = sa00_sr[6] ^ w0[30];
  assign _0022_[7] = sa00_sr[7] ^ w0[31];
  assign _0034_[0] = sa01_sr[0] ^ w1[24];
  assign _0034_[1] = sa01_sr[1] ^ w1[25];
  assign _0034_[2] = sa01_sr[2] ^ w1[26];
  assign _0034_[3] = sa01_sr[3] ^ w1[27];
  assign _0034_[4] = sa01_sr[4] ^ w1[28];
  assign _0034_[5] = sa01_sr[5] ^ w1[29];
  assign _0034_[6] = sa01_sr[6] ^ w1[30];
  assign _0034_[7] = sa01_sr[7] ^ w1[31];
  assign _0029_[0] = sa02_sr[0] ^ w2[24];
  assign _0029_[1] = sa02_sr[1] ^ w2[25];
  assign _0029_[2] = sa02_sr[2] ^ w2[26];
  assign _0029_[3] = sa02_sr[3] ^ w2[27];
  assign _0029_[4] = sa02_sr[4] ^ w2[28];
  assign _0029_[5] = sa02_sr[5] ^ w2[29];
  assign _0029_[6] = sa02_sr[6] ^ w2[30];
  assign _0029_[7] = sa02_sr[7] ^ w2[31];
  assign _0025_[0] = sa03_sr[0] ^ w3[24];
  assign _0025_[1] = sa03_sr[1] ^ w3[25];
  assign _0025_[2] = sa03_sr[2] ^ w3[26];
  assign _0025_[3] = sa03_sr[3] ^ w3[27];
  assign _0025_[4] = sa03_sr[4] ^ w3[28];
  assign _0025_[5] = sa03_sr[5] ^ w3[29];
  assign _0025_[6] = sa03_sr[6] ^ w3[30];
  assign _0025_[7] = sa03_sr[7] ^ w3[31];
  assign _0021_[0] = sa10_sr[0] ^ w0[16];
  assign _0021_[1] = sa10_sr[1] ^ w0[17];
  assign _0021_[2] = sa10_sr[2] ^ w0[18];
  assign _0021_[3] = sa10_sr[3] ^ w0[19];
  assign _0021_[4] = sa10_sr[4] ^ w0[20];
  assign _0021_[5] = sa10_sr[5] ^ w0[21];
  assign _0021_[6] = sa10_sr[6] ^ w0[22];
  assign _0021_[7] = sa10_sr[7] ^ w0[23];
  assign _0033_[0] = sa11_sr[0] ^ w1[16];
  assign _0033_[1] = sa11_sr[1] ^ w1[17];
  assign _0033_[2] = sa11_sr[2] ^ w1[18];
  assign _0033_[3] = sa11_sr[3] ^ w1[19];
  assign _0033_[4] = sa11_sr[4] ^ w1[20];
  assign _0033_[5] = sa11_sr[5] ^ w1[21];
  assign _0033_[6] = sa11_sr[6] ^ w1[22];
  assign _0033_[7] = sa11_sr[7] ^ w1[23];
  assign _0028_[0] = sa12_sr[0] ^ w2[16];
  assign _0028_[1] = sa12_sr[1] ^ w2[17];
  assign _0028_[2] = sa12_sr[2] ^ w2[18];
  assign _0028_[3] = sa12_sr[3] ^ w2[19];
  assign _0028_[4] = sa12_sr[4] ^ w2[20];
  assign _0028_[5] = sa12_sr[5] ^ w2[21];
  assign _0028_[6] = sa12_sr[6] ^ w2[22];
  assign _0028_[7] = sa12_sr[7] ^ w2[23];
  assign _0024_[0] = sa10_sub[0] ^ w3[16];
  assign _0024_[1] = sa10_sub[1] ^ w3[17];
  assign _0024_[2] = sa10_sub[2] ^ w3[18];
  assign _0024_[3] = sa10_sub[3] ^ w3[19];
  assign _0024_[4] = sa10_sub[4] ^ w3[20];
  assign _0024_[5] = sa10_sub[5] ^ w3[21];
  assign _0024_[6] = sa10_sub[6] ^ w3[22];
  assign _0024_[7] = sa10_sub[7] ^ w3[23];
  assign _0020_[0] = sa20_sr[0] ^ w0[8];
  assign _0020_[1] = sa20_sr[1] ^ w0[9];
  assign _0020_[2] = sa20_sr[2] ^ w0[10];
  assign _0020_[3] = sa20_sr[3] ^ w0[11];
  assign _0020_[4] = sa20_sr[4] ^ w0[12];
  assign _0020_[5] = sa20_sr[5] ^ w0[13];
  assign _0020_[6] = sa20_sr[6] ^ w0[14];
  assign _0020_[7] = sa20_sr[7] ^ w0[15];
  assign _0031_[0] = sa21_sr[0] ^ w1[8];
  assign _0031_[1] = sa21_sr[1] ^ w1[9];
  assign _0031_[2] = sa21_sr[2] ^ w1[10];
  assign _0031_[3] = sa21_sr[3] ^ w1[11];
  assign _0031_[4] = sa21_sr[4] ^ w1[12];
  assign _0031_[5] = sa21_sr[5] ^ w1[13];
  assign _0031_[6] = sa21_sr[6] ^ w1[14];
  assign _0031_[7] = sa21_sr[7] ^ w1[15];
  assign _0027_[0] = sa20_sub[0] ^ w2[8];
  assign _0027_[1] = sa20_sub[1] ^ w2[9];
  assign _0027_[2] = sa20_sub[2] ^ w2[10];
  assign _0027_[3] = sa20_sub[3] ^ w2[11];
  assign _0027_[4] = sa20_sub[4] ^ w2[12];
  assign _0027_[5] = sa20_sub[5] ^ w2[13];
  assign _0027_[6] = sa20_sub[6] ^ w2[14];
  assign _0027_[7] = sa20_sub[7] ^ w2[15];
  assign _0023_[0] = sa21_sub[0] ^ w3[8];
  assign _0023_[1] = sa21_sub[1] ^ w3[9];
  assign _0023_[2] = sa21_sub[2] ^ w3[10];
  assign _0023_[3] = sa21_sub[3] ^ w3[11];
  assign _0023_[4] = sa21_sub[4] ^ w3[12];
  assign _0023_[5] = sa21_sub[5] ^ w3[13];
  assign _0023_[6] = sa21_sub[6] ^ w3[14];
  assign _0023_[7] = sa21_sub[7] ^ w3[15];
  assign _0019_[0] = sa30_sr[0] ^ w0[0];
  assign _0019_[1] = sa30_sr[1] ^ w0[1];
  assign _0019_[2] = sa30_sr[2] ^ w0[2];
  assign _0019_[3] = sa30_sr[3] ^ w0[3];
  assign _0019_[4] = sa30_sr[4] ^ w0[4];
  assign _0019_[5] = sa30_sr[5] ^ w0[5];
  assign _0019_[6] = sa30_sr[6] ^ w0[6];
  assign _0019_[7] = sa30_sr[7] ^ w0[7];
  assign _0030_[0] = sa30_sub[0] ^ w1[0];
  assign _0030_[1] = sa30_sub[1] ^ w1[1];
  assign _0030_[2] = sa30_sub[2] ^ w1[2];
  assign _0030_[3] = sa30_sub[3] ^ w1[3];
  assign _0030_[4] = sa30_sub[4] ^ w1[4];
  assign _0030_[5] = sa30_sub[5] ^ w1[5];
  assign _0030_[6] = sa30_sub[6] ^ w1[6];
  assign _0030_[7] = sa30_sub[7] ^ w1[7];
  assign _0026_[0] = sa31_sub[0] ^ w2[0];
  assign _0026_[1] = sa31_sub[1] ^ w2[1];
  assign _0026_[2] = sa31_sub[2] ^ w2[2];
  assign _0026_[3] = sa31_sub[3] ^ w2[3];
  assign _0026_[4] = sa31_sub[4] ^ w2[4];
  assign _0026_[5] = sa31_sub[5] ^ w2[5];
  assign _0026_[6] = sa31_sub[6] ^ w2[6];
  assign _0026_[7] = sa31_sub[7] ^ w2[7];
  assign _0032_[0] = sa32_sub[0] ^ w3[0];
  assign _0032_[1] = sa32_sub[1] ^ w3[1];
  assign _0032_[2] = sa32_sub[2] ^ w3[2];
  assign _0032_[3] = sa32_sub[3] ^ w3[3];
  assign _0032_[4] = sa32_sub[4] ^ w3[4];
  assign _0032_[5] = sa32_sub[5] ^ w3[5];
  assign _0032_[6] = sa32_sub[6] ^ w3[6];
  assign _0032_[7] = sa32_sub[7] ^ w3[7];
  always @(posedge clk)
      dcnt[0] <= _0000_[0];
  always @(posedge clk)
      dcnt[1] <= _0000_[1];
  always @(posedge clk)
      dcnt[2] <= _0000_[2];
  always @(posedge clk)
      dcnt[3] <= _0000_[3];
  always @(posedge clk)
      done <= _0001_;
  always @(posedge clk)
      text_in_r[0] <= _0018_[0];
  always @(posedge clk)
      text_in_r[100] <= _0018_[100];
  always @(posedge clk)
      text_in_r[101] <= _0018_[101];
  always @(posedge clk)
      text_in_r[102] <= _0018_[102];
  always @(posedge clk)
      text_in_r[103] <= _0018_[103];
  always @(posedge clk)
      text_in_r[104] <= _0018_[104];
  always @(posedge clk)
      text_in_r[105] <= _0018_[105];
  always @(posedge clk)
      text_in_r[106] <= _0018_[106];
  always @(posedge clk)
      text_in_r[107] <= _0018_[107];
  always @(posedge clk)
      text_in_r[108] <= _0018_[108];
  always @(posedge clk)
      text_in_r[109] <= _0018_[109];
  always @(posedge clk)
      text_in_r[10] <= _0018_[10];
  always @(posedge clk)
      text_in_r[110] <= _0018_[110];
  always @(posedge clk)
      text_in_r[111] <= _0018_[111];
  always @(posedge clk)
      text_in_r[112] <= _0018_[112];
  always @(posedge clk)
      text_in_r[113] <= _0018_[113];
  always @(posedge clk)
      text_in_r[114] <= _0018_[114];
  always @(posedge clk)
      text_in_r[115] <= _0018_[115];
  always @(posedge clk)
      text_in_r[116] <= _0018_[116];
  always @(posedge clk)
      text_in_r[117] <= _0018_[117];
  always @(posedge clk)
      text_in_r[118] <= _0018_[118];
  always @(posedge clk)
      text_in_r[119] <= _0018_[119];
  always @(posedge clk)
      text_in_r[11] <= _0018_[11];
  always @(posedge clk)
      text_in_r[120] <= _0018_[120];
  always @(posedge clk)
      text_in_r[121] <= _0018_[121];
  always @(posedge clk)
      text_in_r[122] <= _0018_[122];
  always @(posedge clk)
      text_in_r[123] <= _0018_[123];
  always @(posedge clk)
      text_in_r[124] <= _0018_[124];
  always @(posedge clk)
      text_in_r[125] <= _0018_[125];
  always @(posedge clk)
      text_in_r[126] <= _0018_[126];
  always @(posedge clk)
      text_in_r[127] <= _0018_[127];
  always @(posedge clk)
      text_in_r[12] <= _0018_[12];
  always @(posedge clk)
      text_in_r[13] <= _0018_[13];
  always @(posedge clk)
      text_in_r[14] <= _0018_[14];
  always @(posedge clk)
      text_in_r[15] <= _0018_[15];
  always @(posedge clk)
      text_in_r[16] <= _0018_[16];
  always @(posedge clk)
      text_in_r[17] <= _0018_[17];
  always @(posedge clk)
      text_in_r[18] <= _0018_[18];
  always @(posedge clk)
      text_in_r[19] <= _0018_[19];
  always @(posedge clk)
      text_in_r[1] <= _0018_[1];
  always @(posedge clk)
      text_in_r[20] <= _0018_[20];
  always @(posedge clk)
      text_in_r[21] <= _0018_[21];
  always @(posedge clk)
      text_in_r[22] <= _0018_[22];
  always @(posedge clk)
      text_in_r[23] <= _0018_[23];
  always @(posedge clk)
      text_in_r[24] <= _0018_[24];
  always @(posedge clk)
      text_in_r[25] <= _0018_[25];
  always @(posedge clk)
      text_in_r[26] <= _0018_[26];
  always @(posedge clk)
      text_in_r[27] <= _0018_[27];
  always @(posedge clk)
      text_in_r[28] <= _0018_[28];
  always @(posedge clk)
      text_in_r[29] <= _0018_[29];
  always @(posedge clk)
      text_in_r[2] <= _0018_[2];
  always @(posedge clk)
      text_in_r[30] <= _0018_[30];
  always @(posedge clk)
      text_in_r[31] <= _0018_[31];
  always @(posedge clk)
      text_in_r[32] <= _0018_[32];
  always @(posedge clk)
      text_in_r[33] <= _0018_[33];
  always @(posedge clk)
      text_in_r[34] <= _0018_[34];
  always @(posedge clk)
      text_in_r[35] <= _0018_[35];
  always @(posedge clk)
      text_in_r[36] <= _0018_[36];
  always @(posedge clk)
      text_in_r[37] <= _0018_[37];
  always @(posedge clk)
      text_in_r[38] <= _0018_[38];
  always @(posedge clk)
      text_in_r[39] <= _0018_[39];
  always @(posedge clk)
      text_in_r[3] <= _0018_[3];
  always @(posedge clk)
      text_in_r[40] <= _0018_[40];
  always @(posedge clk)
      text_in_r[41] <= _0018_[41];
  always @(posedge clk)
      text_in_r[42] <= _0018_[42];
  always @(posedge clk)
      text_in_r[43] <= _0018_[43];
  always @(posedge clk)
      text_in_r[44] <= _0018_[44];
  always @(posedge clk)
      text_in_r[45] <= _0018_[45];
  always @(posedge clk)
      text_in_r[46] <= _0018_[46];
  always @(posedge clk)
      text_in_r[47] <= _0018_[47];
  always @(posedge clk)
      text_in_r[48] <= _0018_[48];
  always @(posedge clk)
      text_in_r[49] <= _0018_[49];
  always @(posedge clk)
      text_in_r[4] <= _0018_[4];
  always @(posedge clk)
      text_in_r[50] <= _0018_[50];
  always @(posedge clk)
      text_in_r[51] <= _0018_[51];
  always @(posedge clk)
      text_in_r[52] <= _0018_[52];
  always @(posedge clk)
      text_in_r[53] <= _0018_[53];
  always @(posedge clk)
      text_in_r[54] <= _0018_[54];
  always @(posedge clk)
      text_in_r[55] <= _0018_[55];
  always @(posedge clk)
      text_in_r[56] <= _0018_[56];
  always @(posedge clk)
      text_in_r[57] <= _0018_[57];
  always @(posedge clk)
      text_in_r[58] <= _0018_[58];
  always @(posedge clk)
      text_in_r[59] <= _0018_[59];
  always @(posedge clk)
      text_in_r[5] <= _0018_[5];
  always @(posedge clk)
      text_in_r[60] <= _0018_[60];
  always @(posedge clk)
      text_in_r[61] <= _0018_[61];
  always @(posedge clk)
      text_in_r[62] <= _0018_[62];
  always @(posedge clk)
      text_in_r[63] <= _0018_[63];
  always @(posedge clk)
      text_in_r[64] <= _0018_[64];
  always @(posedge clk)
      text_in_r[65] <= _0018_[65];
  always @(posedge clk)
      text_in_r[66] <= _0018_[66];
  always @(posedge clk)
      text_in_r[67] <= _0018_[67];
  always @(posedge clk)
      text_in_r[68] <= _0018_[68];
  always @(posedge clk)
      text_in_r[69] <= _0018_[69];
  always @(posedge clk)
      text_in_r[6] <= _0018_[6];
  always @(posedge clk)
      text_in_r[70] <= _0018_[70];
  always @(posedge clk)
      text_in_r[71] <= _0018_[71];
  always @(posedge clk)
      text_in_r[72] <= _0018_[72];
  always @(posedge clk)
      text_in_r[73] <= _0018_[73];
  always @(posedge clk)
      text_in_r[74] <= _0018_[74];
  always @(posedge clk)
      text_in_r[75] <= _0018_[75];
  always @(posedge clk)
      text_in_r[76] <= _0018_[76];
  always @(posedge clk)
      text_in_r[77] <= _0018_[77];
  always @(posedge clk)
      text_in_r[78] <= _0018_[78];
  always @(posedge clk)
      text_in_r[79] <= _0018_[79];
  always @(posedge clk)
      text_in_r[7] <= _0018_[7];
  always @(posedge clk)
      text_in_r[80] <= _0018_[80];
  always @(posedge clk)
      text_in_r[81] <= _0018_[81];
  always @(posedge clk)
      text_in_r[82] <= _0018_[82];
  always @(posedge clk)
      text_in_r[83] <= _0018_[83];
  always @(posedge clk)
      text_in_r[84] <= _0018_[84];
  always @(posedge clk)
      text_in_r[85] <= _0018_[85];
  always @(posedge clk)
      text_in_r[86] <= _0018_[86];
  always @(posedge clk)
      text_in_r[87] <= _0018_[87];
  always @(posedge clk)
      text_in_r[88] <= _0018_[88];
  always @(posedge clk)
      text_in_r[89] <= _0018_[89];
  always @(posedge clk)
      text_in_r[8] <= _0018_[8];
  always @(posedge clk)
      text_in_r[90] <= _0018_[90];
  always @(posedge clk)
      text_in_r[91] <= _0018_[91];
  always @(posedge clk)
      text_in_r[92] <= _0018_[92];
  always @(posedge clk)
      text_in_r[93] <= _0018_[93];
  always @(posedge clk)
      text_in_r[94] <= _0018_[94];
  always @(posedge clk)
      text_in_r[95] <= _0018_[95];
  always @(posedge clk)
      text_in_r[96] <= _0018_[96];
  always @(posedge clk)
      text_in_r[97] <= _0018_[97];
  always @(posedge clk)
      text_in_r[98] <= _0018_[98];
  always @(posedge clk)
      text_in_r[99] <= _0018_[99];
  always @(posedge clk)
      text_in_r[9] <= _0018_[9];
  always @(posedge clk)
      ld_r <= ld;
  always @(posedge clk)
      sa33[0] <= _0017_[0];
  always @(posedge clk)
      sa33[1] <= _0017_[1];
  always @(posedge clk)
      sa33[2] <= _0017_[2];
  always @(posedge clk)
      sa33[3] <= _0017_[3];
  always @(posedge clk)
      sa33[4] <= _0017_[4];
  always @(posedge clk)
      sa33[5] <= _0017_[5];
  always @(posedge clk)
      sa33[6] <= _0017_[6];
  always @(posedge clk)
      sa33[7] <= _0017_[7];
  always @(posedge clk)
      sa23[0] <= _0013_[0];
  always @(posedge clk)
      sa23[1] <= _0013_[1];
  always @(posedge clk)
      sa23[2] <= _0013_[2];
  always @(posedge clk)
      sa23[3] <= _0013_[3];
  always @(posedge clk)
      sa23[4] <= _0013_[4];
  always @(posedge clk)
      sa23[5] <= _0013_[5];
  always @(posedge clk)
      sa23[6] <= _0013_[6];
  always @(posedge clk)
      sa23[7] <= _0013_[7];
  always @(posedge clk)
      sa13[0] <= _0009_[0];
  always @(posedge clk)
      sa13[1] <= _0009_[1];
  always @(posedge clk)
      sa13[2] <= _0009_[2];
  always @(posedge clk)
      sa13[3] <= _0009_[3];
  always @(posedge clk)
      sa13[4] <= _0009_[4];
  always @(posedge clk)
      sa13[5] <= _0009_[5];
  always @(posedge clk)
      sa13[6] <= _0009_[6];
  always @(posedge clk)
      sa13[7] <= _0009_[7];
  always @(posedge clk)
      sa03[0] <= _0005_[0];
  always @(posedge clk)
      sa03[1] <= _0005_[1];
  always @(posedge clk)
      sa03[2] <= _0005_[2];
  always @(posedge clk)
      sa03[3] <= _0005_[3];
  always @(posedge clk)
      sa03[4] <= _0005_[4];
  always @(posedge clk)
      sa03[5] <= _0005_[5];
  always @(posedge clk)
      sa03[6] <= _0005_[6];
  always @(posedge clk)
      sa03[7] <= _0005_[7];
  always @(posedge clk)
      sa32[0] <= _0016_[0];
  always @(posedge clk)
      sa32[1] <= _0016_[1];
  always @(posedge clk)
      sa32[2] <= _0016_[2];
  always @(posedge clk)
      sa32[3] <= _0016_[3];
  always @(posedge clk)
      sa32[4] <= _0016_[4];
  always @(posedge clk)
      sa32[5] <= _0016_[5];
  always @(posedge clk)
      sa32[6] <= _0016_[6];
  always @(posedge clk)
      sa32[7] <= _0016_[7];
  always @(posedge clk)
      sa22[0] <= _0012_[0];
  always @(posedge clk)
      sa22[1] <= _0012_[1];
  always @(posedge clk)
      sa22[2] <= _0012_[2];
  always @(posedge clk)
      sa22[3] <= _0012_[3];
  always @(posedge clk)
      sa22[4] <= _0012_[4];
  always @(posedge clk)
      sa22[5] <= _0012_[5];
  always @(posedge clk)
      sa22[6] <= _0012_[6];
  always @(posedge clk)
      sa22[7] <= _0012_[7];
  always @(posedge clk)
      sa12[0] <= _0008_[0];
  always @(posedge clk)
      sa12[1] <= _0008_[1];
  always @(posedge clk)
      sa12[2] <= _0008_[2];
  always @(posedge clk)
      sa12[3] <= _0008_[3];
  always @(posedge clk)
      sa12[4] <= _0008_[4];
  always @(posedge clk)
      sa12[5] <= _0008_[5];
  always @(posedge clk)
      sa12[6] <= _0008_[6];
  always @(posedge clk)
      sa12[7] <= _0008_[7];
  always @(posedge clk)
      sa02[0] <= _0004_[0];
  always @(posedge clk)
      sa02[1] <= _0004_[1];
  always @(posedge clk)
      sa02[2] <= _0004_[2];
  always @(posedge clk)
      sa02[3] <= _0004_[3];
  always @(posedge clk)
      sa02[4] <= _0004_[4];
  always @(posedge clk)
      sa02[5] <= _0004_[5];
  always @(posedge clk)
      sa02[6] <= _0004_[6];
  always @(posedge clk)
      sa02[7] <= _0004_[7];
  always @(posedge clk)
      sa31[0] <= _0015_[0];
  always @(posedge clk)
      sa31[1] <= _0015_[1];
  always @(posedge clk)
      sa31[2] <= _0015_[2];
  always @(posedge clk)
      sa31[3] <= _0015_[3];
  always @(posedge clk)
      sa31[4] <= _0015_[4];
  always @(posedge clk)
      sa31[5] <= _0015_[5];
  always @(posedge clk)
      sa31[6] <= _0015_[6];
  always @(posedge clk)
      sa31[7] <= _0015_[7];
  always @(posedge clk)
      sa21[0] <= _0011_[0];
  always @(posedge clk)
      sa21[1] <= _0011_[1];
  always @(posedge clk)
      sa21[2] <= _0011_[2];
  always @(posedge clk)
      sa21[3] <= _0011_[3];
  always @(posedge clk)
      sa21[4] <= _0011_[4];
  always @(posedge clk)
      sa21[5] <= _0011_[5];
  always @(posedge clk)
      sa21[6] <= _0011_[6];
  always @(posedge clk)
      sa21[7] <= _0011_[7];
  always @(posedge clk)
      sa11[0] <= _0007_[0];
  always @(posedge clk)
      sa11[1] <= _0007_[1];
  always @(posedge clk)
      sa11[2] <= _0007_[2];
  always @(posedge clk)
      sa11[3] <= _0007_[3];
  always @(posedge clk)
      sa11[4] <= _0007_[4];
  always @(posedge clk)
      sa11[5] <= _0007_[5];
  always @(posedge clk)
      sa11[6] <= _0007_[6];
  always @(posedge clk)
      sa11[7] <= _0007_[7];
  always @(posedge clk)
      sa01[0] <= _0003_[0];
  always @(posedge clk)
      sa01[1] <= _0003_[1];
  always @(posedge clk)
      sa01[2] <= _0003_[2];
  always @(posedge clk)
      sa01[3] <= _0003_[3];
  always @(posedge clk)
      sa01[4] <= _0003_[4];
  always @(posedge clk)
      sa01[5] <= _0003_[5];
  always @(posedge clk)
      sa01[6] <= _0003_[6];
  always @(posedge clk)
      sa01[7] <= _0003_[7];
  always @(posedge clk)
      sa30[0] <= _0014_[0];
  always @(posedge clk)
      sa30[1] <= _0014_[1];
  always @(posedge clk)
      sa30[2] <= _0014_[2];
  always @(posedge clk)
      sa30[3] <= _0014_[3];
  always @(posedge clk)
      sa30[4] <= _0014_[4];
  always @(posedge clk)
      sa30[5] <= _0014_[5];
  always @(posedge clk)
      sa30[6] <= _0014_[6];
  always @(posedge clk)
      sa30[7] <= _0014_[7];
  always @(posedge clk)
      sa20[0] <= _0010_[0];
  always @(posedge clk)
      sa20[1] <= _0010_[1];
  always @(posedge clk)
      sa20[2] <= _0010_[2];
  always @(posedge clk)
      sa20[3] <= _0010_[3];
  always @(posedge clk)
      sa20[4] <= _0010_[4];
  always @(posedge clk)
      sa20[5] <= _0010_[5];
  always @(posedge clk)
      sa20[6] <= _0010_[6];
  always @(posedge clk)
      sa20[7] <= _0010_[7];
  always @(posedge clk)
      sa10[0] <= _0006_[0];
  always @(posedge clk)
      sa10[1] <= _0006_[1];
  always @(posedge clk)
      sa10[2] <= _0006_[2];
  always @(posedge clk)
      sa10[3] <= _0006_[3];
  always @(posedge clk)
      sa10[4] <= _0006_[4];
  always @(posedge clk)
      sa10[5] <= _0006_[5];
  always @(posedge clk)
      sa10[6] <= _0006_[6];
  always @(posedge clk)
      sa10[7] <= _0006_[7];
  always @(posedge clk)
      sa00[0] <= _0002_[0];
  always @(posedge clk)
      sa00[1] <= _0002_[1];
  always @(posedge clk)
      sa00[2] <= _0002_[2];
  always @(posedge clk)
      sa00[3] <= _0002_[3];
  always @(posedge clk)
      sa00[4] <= _0002_[4];
  always @(posedge clk)
      sa00[5] <= _0002_[5];
  always @(posedge clk)
      sa00[6] <= _0002_[6];
  always @(posedge clk)
      sa00[7] <= _0002_[7];
  always @(posedge clk)
      text_out[120] <= _0022_[0];
  always @(posedge clk)
      text_out[121] <= _0022_[1];
  always @(posedge clk)
      text_out[122] <= _0022_[2];
  always @(posedge clk)
      text_out[123] <= _0022_[3];
  always @(posedge clk)
      text_out[124] <= _0022_[4];
  always @(posedge clk)
      text_out[125] <= _0022_[5];
  always @(posedge clk)
      text_out[126] <= _0022_[6];
  always @(posedge clk)
      text_out[127] <= _0022_[7];
  always @(posedge clk)
      text_out[88] <= _0034_[0];
  always @(posedge clk)
      text_out[89] <= _0034_[1];
  always @(posedge clk)
      text_out[90] <= _0034_[2];
  always @(posedge clk)
      text_out[91] <= _0034_[3];
  always @(posedge clk)
      text_out[92] <= _0034_[4];
  always @(posedge clk)
      text_out[93] <= _0034_[5];
  always @(posedge clk)
      text_out[94] <= _0034_[6];
  always @(posedge clk)
      text_out[95] <= _0034_[7];
  always @(posedge clk)
      text_out[56] <= _0029_[0];
  always @(posedge clk)
      text_out[57] <= _0029_[1];
  always @(posedge clk)
      text_out[58] <= _0029_[2];
  always @(posedge clk)
      text_out[59] <= _0029_[3];
  always @(posedge clk)
      text_out[60] <= _0029_[4];
  always @(posedge clk)
      text_out[61] <= _0029_[5];
  always @(posedge clk)
      text_out[62] <= _0029_[6];
  always @(posedge clk)
      text_out[63] <= _0029_[7];
  always @(posedge clk)
      text_out[24] <= _0025_[0];
  always @(posedge clk)
      text_out[25] <= _0025_[1];
  always @(posedge clk)
      text_out[26] <= _0025_[2];
  always @(posedge clk)
      text_out[27] <= _0025_[3];
  always @(posedge clk)
      text_out[28] <= _0025_[4];
  always @(posedge clk)
      text_out[29] <= _0025_[5];
  always @(posedge clk)
      text_out[30] <= _0025_[6];
  always @(posedge clk)
      text_out[31] <= _0025_[7];
  always @(posedge clk)
      text_out[112] <= _0021_[0];
  always @(posedge clk)
      text_out[113] <= _0021_[1];
  always @(posedge clk)
      text_out[114] <= _0021_[2];
  always @(posedge clk)
      text_out[115] <= _0021_[3];
  always @(posedge clk)
      text_out[116] <= _0021_[4];
  always @(posedge clk)
      text_out[117] <= _0021_[5];
  always @(posedge clk)
      text_out[118] <= _0021_[6];
  always @(posedge clk)
      text_out[119] <= _0021_[7];
  always @(posedge clk)
      text_out[80] <= _0033_[0];
  always @(posedge clk)
      text_out[81] <= _0033_[1];
  always @(posedge clk)
      text_out[82] <= _0033_[2];
  always @(posedge clk)
      text_out[83] <= _0033_[3];
  always @(posedge clk)
      text_out[84] <= _0033_[4];
  always @(posedge clk)
      text_out[85] <= _0033_[5];
  always @(posedge clk)
      text_out[86] <= _0033_[6];
  always @(posedge clk)
      text_out[87] <= _0033_[7];
  always @(posedge clk)
      text_out[48] <= _0028_[0];
  always @(posedge clk)
      text_out[49] <= _0028_[1];
  always @(posedge clk)
      text_out[50] <= _0028_[2];
  always @(posedge clk)
      text_out[51] <= _0028_[3];
  always @(posedge clk)
      text_out[52] <= _0028_[4];
  always @(posedge clk)
      text_out[53] <= _0028_[5];
  always @(posedge clk)
      text_out[54] <= _0028_[6];
  always @(posedge clk)
      text_out[55] <= _0028_[7];
  always @(posedge clk)
      text_out[16] <= _0024_[0];
  always @(posedge clk)
      text_out[17] <= _0024_[1];
  always @(posedge clk)
      text_out[18] <= _0024_[2];
  always @(posedge clk)
      text_out[19] <= _0024_[3];
  always @(posedge clk)
      text_out[20] <= _0024_[4];
  always @(posedge clk)
      text_out[21] <= _0024_[5];
  always @(posedge clk)
      text_out[22] <= _0024_[6];
  always @(posedge clk)
      text_out[23] <= _0024_[7];
  always @(posedge clk)
      text_out[104] <= _0020_[0];
  always @(posedge clk)
      text_out[105] <= _0020_[1];
  always @(posedge clk)
      text_out[106] <= _0020_[2];
  always @(posedge clk)
      text_out[107] <= _0020_[3];
  always @(posedge clk)
      text_out[108] <= _0020_[4];
  always @(posedge clk)
      text_out[109] <= _0020_[5];
  always @(posedge clk)
      text_out[110] <= _0020_[6];
  always @(posedge clk)
      text_out[111] <= _0020_[7];
  always @(posedge clk)
      text_out[72] <= _0031_[0];
  always @(posedge clk)
      text_out[73] <= _0031_[1];
  always @(posedge clk)
      text_out[74] <= _0031_[2];
  always @(posedge clk)
      text_out[75] <= _0031_[3];
  always @(posedge clk)
      text_out[76] <= _0031_[4];
  always @(posedge clk)
      text_out[77] <= _0031_[5];
  always @(posedge clk)
      text_out[78] <= _0031_[6];
  always @(posedge clk)
      text_out[79] <= _0031_[7];
  always @(posedge clk)
      text_out[40] <= _0027_[0];
  always @(posedge clk)
      text_out[41] <= _0027_[1];
  always @(posedge clk)
      text_out[42] <= _0027_[2];
  always @(posedge clk)
      text_out[43] <= _0027_[3];
  always @(posedge clk)
      text_out[44] <= _0027_[4];
  always @(posedge clk)
      text_out[45] <= _0027_[5];
  always @(posedge clk)
      text_out[46] <= _0027_[6];
  always @(posedge clk)
      text_out[47] <= _0027_[7];
  always @(posedge clk)
      text_out[8] <= _0023_[0];
  always @(posedge clk)
      text_out[9] <= _0023_[1];
  always @(posedge clk)
      text_out[10] <= _0023_[2];
  always @(posedge clk)
      text_out[11] <= _0023_[3];
  always @(posedge clk)
      text_out[12] <= _0023_[4];
  always @(posedge clk)
      text_out[13] <= _0023_[5];
  always @(posedge clk)
      text_out[14] <= _0023_[6];
  always @(posedge clk)
      text_out[15] <= _0023_[7];
  always @(posedge clk)
      text_out[96] <= _0019_[0];
  always @(posedge clk)
      text_out[97] <= _0019_[1];
  always @(posedge clk)
      text_out[98] <= _0019_[2];
  always @(posedge clk)
      text_out[99] <= _0019_[3];
  always @(posedge clk)
      text_out[100] <= _0019_[4];
  always @(posedge clk)
      text_out[101] <= _0019_[5];
  always @(posedge clk)
      text_out[102] <= _0019_[6];
  always @(posedge clk)
      text_out[103] <= _0019_[7];
  always @(posedge clk)
      text_out[64] <= _0030_[0];
  always @(posedge clk)
      text_out[65] <= _0030_[1];
  always @(posedge clk)
      text_out[66] <= _0030_[2];
  always @(posedge clk)
      text_out[67] <= _0030_[3];
  always @(posedge clk)
      text_out[68] <= _0030_[4];
  always @(posedge clk)
      text_out[69] <= _0030_[5];
  always @(posedge clk)
      text_out[70] <= _0030_[6];
  always @(posedge clk)
      text_out[71] <= _0030_[7];
  always @(posedge clk)
      text_out[32] <= _0026_[0];
  always @(posedge clk)
      text_out[33] <= _0026_[1];
  always @(posedge clk)
      text_out[34] <= _0026_[2];
  always @(posedge clk)
      text_out[35] <= _0026_[3];
  always @(posedge clk)
      text_out[36] <= _0026_[4];
  always @(posedge clk)
      text_out[37] <= _0026_[5];
  always @(posedge clk)
      text_out[38] <= _0026_[6];
  always @(posedge clk)
      text_out[39] <= _0026_[7];
  always @(posedge clk)
      text_out[0] <= _0032_[0];
  always @(posedge clk)
      text_out[1] <= _0032_[1];
  always @(posedge clk)
      text_out[2] <= _0032_[2];
  always @(posedge clk)
      text_out[3] <= _0032_[3];
  always @(posedge clk)
      text_out[4] <= _0032_[4];
  always @(posedge clk)
      text_out[5] <= _0032_[5];
  always @(posedge clk)
      text_out[6] <= _0032_[6];
  always @(posedge clk)
      text_out[7] <= _0032_[7];
  aes_key_expand_128 u0 (
    .clk(clk),
    .key(key),
    .kld(ld),
    .wo_0(w0),
    .wo_1(w1),
    .wo_2(w2),
    .wo_3(w3)
  );
  aes_sbox us00 (
    .a(sa00),
    .d(sa00_sr)
  );
  aes_sbox us01 (
    .a(sa01),
    .d(sa01_sr)
  );
  aes_sbox us02 (
    .a(sa02),
    .d(sa02_sr)
  );
  aes_sbox us03 (
    .a(sa03),
    .d(sa03_sr)
  );
  aes_sbox us10 (
    .a(sa10),
    .d(sa10_sub)
  );
  aes_sbox us11 (
    .a(sa11),
    .d(sa10_sr)
  );
  aes_sbox us12 (
    .a(sa12),
    .d(sa11_sr)
  );
  aes_sbox us13 (
    .a(sa13),
    .d(sa12_sr)
  );
  aes_sbox us20 (
    .a(sa20),
    .d(sa20_sub)
  );
  aes_sbox us21 (
    .a(sa21),
    .d(sa21_sub)
  );
  aes_sbox us22 (
    .a(sa22),
    .d(sa20_sr)
  );
  aes_sbox us23 (
    .a(sa23),
    .d(sa21_sr)
  );
  aes_sbox us30 (
    .a(sa30),
    .d(sa30_sub)
  );
  aes_sbox us31 (
    .a(sa31),
    .d(sa31_sub)
  );
  aes_sbox us32 (
    .a(sa32),
    .d(sa32_sub)
  );
  aes_sbox us33 (
    .a(sa33),
    .d(sa30_sr)
  );
  assign sa00_sub = sa00_sr;
  assign sa01_sub = sa01_sr;
  assign sa02_sub = sa02_sr;
  assign sa03_sub = sa03_sr;
  assign sa11_sub = sa10_sr;
  assign sa12_sub = sa11_sr;
  assign sa13_sr = sa10_sub;
  assign sa13_sub = sa12_sr;
  assign sa22_sr = sa20_sub;
  assign sa22_sub = sa20_sr;
  assign sa23_sr = sa21_sub;
  assign sa23_sub = sa21_sr;
  assign sa31_sr = sa30_sub;
  assign sa32_sr = sa31_sub;
  assign sa33_sr = sa32_sub;
  assign sa33_sub = sa30_sr;
endmodule

module aes_key_expand_128(clk, kld, key, wo_0, wo_1, wo_2, wo_3);
  wire [31:0] _0000_;
  wire [31:0] _0001_;
  wire [31:0] _0002_;
  wire [31:0] _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  input clk;
  input [127:0] key;
  input kld;
  wire [31:0] rcon;
  wire [31:0] subword;
  reg [31:0] tmp_w;
  output [31:0] wo_0;
  reg [31:0] wo_0;
  output [31:0] wo_1;
  reg [31:0] wo_1;
  output [31:0] wo_2;
  reg [31:0] wo_2;
  output [31:0] wo_3;
  assign _0078_ = wo_0[0] ^ subword[0];
  assign _0079_ = _0078_ ^ rcon[0];
  assign _0000_[0] = kld ? key[96] : _0079_;
  assign _0080_ = wo_0[10] ^ subword[10];
  assign _0081_ = _0080_ ^ rcon[10];
  assign _0000_[10] = kld ? key[106] : _0081_;
  assign _0082_ = wo_0[11] ^ subword[11];
  assign _0083_ = _0082_ ^ rcon[11];
  assign _0000_[11] = kld ? key[107] : _0083_;
  assign _0084_ = wo_0[12] ^ subword[12];
  assign _0085_ = _0084_ ^ rcon[12];
  assign _0000_[12] = kld ? key[108] : _0085_;
  assign _0086_ = wo_0[13] ^ subword[13];
  assign _0087_ = _0086_ ^ rcon[13];
  assign _0000_[13] = kld ? key[109] : _0087_;
  assign _0088_ = wo_0[14] ^ subword[14];
  assign _0089_ = _0088_ ^ rcon[14];
  assign _0000_[14] = kld ? key[110] : _0089_;
  assign _0090_ = wo_0[15] ^ subword[15];
  assign _0091_ = _0090_ ^ rcon[15];
  assign _0000_[15] = kld ? key[111] : _0091_;
  assign _0092_ = wo_0[16] ^ subword[16];
  assign _0093_ = _0092_ ^ rcon[16];
  assign _0000_[16] = kld ? key[112] : _0093_;
  assign _0094_ = wo_0[17] ^ subword[17];
  assign _0095_ = _0094_ ^ rcon[17];
  assign _0000_[17] = kld ? key[113] : _0095_;
  assign _0096_ = wo_0[18] ^ subword[18];
  assign _0097_ = _0096_ ^ rcon[18];
  assign _0000_[18] = kld ? key[114] : _0097_;
  assign _0098_ = wo_0[19] ^ subword[19];
  assign _0099_ = _0098_ ^ rcon[19];
  assign _0000_[19] = kld ? key[115] : _0099_;
  assign _0100_ = wo_0[1] ^ subword[1];
  assign _0101_ = _0100_ ^ rcon[1];
  assign _0000_[1] = kld ? key[97] : _0101_;
  assign _0102_ = wo_0[20] ^ subword[20];
  assign _0103_ = _0102_ ^ rcon[20];
  assign _0000_[20] = kld ? key[116] : _0103_;
  assign _0104_ = wo_0[21] ^ subword[21];
  assign _0105_ = _0104_ ^ rcon[21];
  assign _0000_[21] = kld ? key[117] : _0105_;
  assign _0106_ = wo_0[22] ^ subword[22];
  assign _0107_ = _0106_ ^ rcon[22];
  assign _0000_[22] = kld ? key[118] : _0107_;
  assign _0108_ = wo_0[23] ^ subword[23];
  assign _0109_ = _0108_ ^ rcon[23];
  assign _0000_[23] = kld ? key[119] : _0109_;
  assign _0110_ = wo_0[24] ^ subword[24];
  assign _0111_ = _0110_ ^ rcon[24];
  assign _0000_[24] = kld ? key[120] : _0111_;
  assign _0112_ = wo_0[25] ^ subword[25];
  assign _0113_ = _0112_ ^ rcon[25];
  assign _0000_[25] = kld ? key[121] : _0113_;
  assign _0114_ = wo_0[26] ^ subword[26];
  assign _0115_ = _0114_ ^ rcon[26];
  assign _0000_[26] = kld ? key[122] : _0115_;
  assign _0116_ = wo_0[27] ^ subword[27];
  assign _0117_ = _0116_ ^ rcon[27];
  assign _0000_[27] = kld ? key[123] : _0117_;
  assign _0118_ = wo_0[28] ^ subword[28];
  assign _0119_ = _0118_ ^ rcon[28];
  assign _0000_[28] = kld ? key[124] : _0119_;
  assign _0120_ = wo_0[29] ^ subword[29];
  assign _0121_ = _0120_ ^ rcon[29];
  assign _0000_[29] = kld ? key[125] : _0121_;
  assign _0122_ = wo_0[2] ^ subword[2];
  assign _0123_ = _0122_ ^ rcon[2];
  assign _0000_[2] = kld ? key[98] : _0123_;
  assign _0124_ = wo_0[30] ^ subword[30];
  assign _0125_ = _0124_ ^ rcon[30];
  assign _0000_[30] = kld ? key[126] : _0125_;
  assign _0126_ = wo_0[31] ^ subword[31];
  assign _0127_ = _0126_ ^ rcon[31];
  assign _0000_[31] = kld ? key[127] : _0127_;
  assign _0128_ = wo_0[3] ^ subword[3];
  assign _0129_ = _0128_ ^ rcon[3];
  assign _0000_[3] = kld ? key[99] : _0129_;
  assign _0130_ = wo_0[4] ^ subword[4];
  assign _0131_ = _0130_ ^ rcon[4];
  assign _0000_[4] = kld ? key[100] : _0131_;
  assign _0132_ = wo_0[5] ^ subword[5];
  assign _0133_ = _0132_ ^ rcon[5];
  assign _0000_[5] = kld ? key[101] : _0133_;
  assign _0134_ = wo_0[6] ^ subword[6];
  assign _0135_ = _0134_ ^ rcon[6];
  assign _0000_[6] = kld ? key[102] : _0135_;
  assign _0136_ = wo_0[7] ^ subword[7];
  assign _0137_ = _0136_ ^ rcon[7];
  assign _0000_[7] = kld ? key[103] : _0137_;
  assign _0138_ = wo_0[8] ^ subword[8];
  assign _0139_ = _0138_ ^ rcon[8];
  assign _0000_[8] = kld ? key[104] : _0139_;
  assign _0140_ = wo_0[9] ^ subword[9];
  assign _0141_ = _0140_ ^ rcon[9];
  assign _0000_[9] = kld ? key[105] : _0141_;
  assign _0142_ = wo_1[0] ^ wo_0[0];
  assign _0143_ = _0142_ ^ subword[0];
  assign _0144_ = _0143_ ^ rcon[0];
  assign _0001_[0] = kld ? key[64] : _0144_;
  assign _0145_ = wo_1[10] ^ wo_0[10];
  assign _0146_ = _0145_ ^ subword[10];
  assign _0147_ = _0146_ ^ rcon[10];
  assign _0001_[10] = kld ? key[74] : _0147_;
  assign _0148_ = wo_1[11] ^ wo_0[11];
  assign _0149_ = _0148_ ^ subword[11];
  assign _0150_ = _0149_ ^ rcon[11];
  assign _0001_[11] = kld ? key[75] : _0150_;
  assign _0151_ = wo_1[12] ^ wo_0[12];
  assign _0152_ = _0151_ ^ subword[12];
  assign _0153_ = _0152_ ^ rcon[12];
  assign _0001_[12] = kld ? key[76] : _0153_;
  assign _0154_ = wo_1[13] ^ wo_0[13];
  assign _0155_ = _0154_ ^ subword[13];
  assign _0156_ = _0155_ ^ rcon[13];
  assign _0001_[13] = kld ? key[77] : _0156_;
  assign _0157_ = wo_1[14] ^ wo_0[14];
  assign _0158_ = _0157_ ^ subword[14];
  assign _0159_ = _0158_ ^ rcon[14];
  assign _0001_[14] = kld ? key[78] : _0159_;
  assign _0160_ = wo_1[15] ^ wo_0[15];
  assign _0161_ = _0160_ ^ subword[15];
  assign _0162_ = _0161_ ^ rcon[15];
  assign _0001_[15] = kld ? key[79] : _0162_;
  assign _0163_ = wo_1[16] ^ wo_0[16];
  assign _0164_ = _0163_ ^ subword[16];
  assign _0165_ = _0164_ ^ rcon[16];
  assign _0001_[16] = kld ? key[80] : _0165_;
  assign _0166_ = wo_1[17] ^ wo_0[17];
  assign _0167_ = _0166_ ^ subword[17];
  assign _0168_ = _0167_ ^ rcon[17];
  assign _0001_[17] = kld ? key[81] : _0168_;
  assign _0169_ = wo_1[18] ^ wo_0[18];
  assign _0170_ = _0169_ ^ subword[18];
  assign _0171_ = _0170_ ^ rcon[18];
  assign _0001_[18] = kld ? key[82] : _0171_;
  assign _0172_ = wo_1[19] ^ wo_0[19];
  assign _0173_ = _0172_ ^ subword[19];
  assign _0174_ = _0173_ ^ rcon[19];
  assign _0001_[19] = kld ? key[83] : _0174_;
  assign _0175_ = wo_1[1] ^ wo_0[1];
  assign _0176_ = _0175_ ^ subword[1];
  assign _0177_ = _0176_ ^ rcon[1];
  assign _0001_[1] = kld ? key[65] : _0177_;
  assign _0178_ = wo_1[20] ^ wo_0[20];
  assign _0179_ = _0178_ ^ subword[20];
  assign _0180_ = _0179_ ^ rcon[20];
  assign _0001_[20] = kld ? key[84] : _0180_;
  assign _0181_ = wo_1[21] ^ wo_0[21];
  assign _0182_ = _0181_ ^ subword[21];
  assign _0183_ = _0182_ ^ rcon[21];
  assign _0001_[21] = kld ? key[85] : _0183_;
  assign _0184_ = wo_1[22] ^ wo_0[22];
  assign _0185_ = _0184_ ^ subword[22];
  assign _0186_ = _0185_ ^ rcon[22];
  assign _0001_[22] = kld ? key[86] : _0186_;
  assign _0187_ = wo_1[23] ^ wo_0[23];
  assign _0188_ = _0187_ ^ subword[23];
  assign _0189_ = _0188_ ^ rcon[23];
  assign _0001_[23] = kld ? key[87] : _0189_;
  assign _0190_ = wo_1[24] ^ wo_0[24];
  assign _0191_ = _0190_ ^ subword[24];
  assign _0192_ = _0191_ ^ rcon[24];
  assign _0001_[24] = kld ? key[88] : _0192_;
  assign _0193_ = wo_1[25] ^ wo_0[25];
  assign _0194_ = _0193_ ^ subword[25];
  assign _0195_ = _0194_ ^ rcon[25];
  assign _0001_[25] = kld ? key[89] : _0195_;
  assign _0196_ = wo_1[26] ^ wo_0[26];
  assign _0197_ = _0196_ ^ subword[26];
  assign _0198_ = _0197_ ^ rcon[26];
  assign _0001_[26] = kld ? key[90] : _0198_;
  assign _0199_ = wo_1[27] ^ wo_0[27];
  assign _0200_ = _0199_ ^ subword[27];
  assign _0201_ = _0200_ ^ rcon[27];
  assign _0001_[27] = kld ? key[91] : _0201_;
  assign _0202_ = wo_1[28] ^ wo_0[28];
  assign _0203_ = _0202_ ^ subword[28];
  assign _0204_ = _0203_ ^ rcon[28];
  assign _0001_[28] = kld ? key[92] : _0204_;
  assign _0205_ = wo_1[29] ^ wo_0[29];
  assign _0206_ = _0205_ ^ subword[29];
  assign _0207_ = _0206_ ^ rcon[29];
  assign _0001_[29] = kld ? key[93] : _0207_;
  assign _0208_ = wo_1[2] ^ wo_0[2];
  assign _0209_ = _0208_ ^ subword[2];
  assign _0210_ = _0209_ ^ rcon[2];
  assign _0001_[2] = kld ? key[66] : _0210_;
  assign _0211_ = wo_1[30] ^ wo_0[30];
  assign _0212_ = _0211_ ^ subword[30];
  assign _0213_ = _0212_ ^ rcon[30];
  assign _0001_[30] = kld ? key[94] : _0213_;
  assign _0214_ = wo_1[31] ^ wo_0[31];
  assign _0215_ = _0214_ ^ subword[31];
  assign _0216_ = _0215_ ^ rcon[31];
  assign _0001_[31] = kld ? key[95] : _0216_;
  assign _0217_ = wo_1[3] ^ wo_0[3];
  assign _0218_ = _0217_ ^ subword[3];
  assign _0219_ = _0218_ ^ rcon[3];
  assign _0001_[3] = kld ? key[67] : _0219_;
  assign _0220_ = wo_1[4] ^ wo_0[4];
  assign _0221_ = _0220_ ^ subword[4];
  assign _0222_ = _0221_ ^ rcon[4];
  assign _0001_[4] = kld ? key[68] : _0222_;
  assign _0223_ = wo_1[5] ^ wo_0[5];
  assign _0224_ = _0223_ ^ subword[5];
  assign _0225_ = _0224_ ^ rcon[5];
  assign _0001_[5] = kld ? key[69] : _0225_;
  assign _0226_ = wo_1[6] ^ wo_0[6];
  assign _0227_ = _0226_ ^ subword[6];
  assign _0228_ = _0227_ ^ rcon[6];
  assign _0001_[6] = kld ? key[70] : _0228_;
  assign _0229_ = wo_1[7] ^ wo_0[7];
  assign _0230_ = _0229_ ^ subword[7];
  assign _0231_ = _0230_ ^ rcon[7];
  assign _0001_[7] = kld ? key[71] : _0231_;
  assign _0232_ = wo_1[8] ^ wo_0[8];
  assign _0233_ = _0232_ ^ subword[8];
  assign _0234_ = _0233_ ^ rcon[8];
  assign _0001_[8] = kld ? key[72] : _0234_;
  assign _0235_ = wo_1[9] ^ wo_0[9];
  assign _0236_ = _0235_ ^ subword[9];
  assign _0237_ = _0236_ ^ rcon[9];
  assign _0001_[9] = kld ? key[73] : _0237_;
  assign _0238_ = ~rcon[0];
  assign _0239_ = ~wo_2[0];
  assign _0240_ = _0239_ ^ wo_0[0];
  assign _0241_ = _0240_ ^ wo_1[0];
  assign _0242_ = _0241_ ^ subword[0];
  assign _0243_ = _0242_ ^ _0238_;
  assign _0002_[0] = kld ? key[32] : _0243_;
  assign _0244_ = ~rcon[10];
  assign _0245_ = ~wo_2[10];
  assign _0246_ = _0245_ ^ wo_0[10];
  assign _0247_ = _0246_ ^ wo_1[10];
  assign _0248_ = _0247_ ^ subword[10];
  assign _0249_ = _0248_ ^ _0244_;
  assign _0002_[10] = kld ? key[42] : _0249_;
  assign _0250_ = ~rcon[11];
  assign _0251_ = ~wo_2[11];
  assign _0252_ = _0251_ ^ wo_0[11];
  assign _0253_ = _0252_ ^ wo_1[11];
  assign _0254_ = _0253_ ^ subword[11];
  assign _0255_ = _0254_ ^ _0250_;
  assign _0002_[11] = kld ? key[43] : _0255_;
  assign _0256_ = ~rcon[12];
  assign _0257_ = ~wo_2[12];
  assign _0258_ = _0257_ ^ wo_0[12];
  assign _0259_ = _0258_ ^ wo_1[12];
  assign _0260_ = _0259_ ^ subword[12];
  assign _0261_ = _0260_ ^ _0256_;
  assign _0002_[12] = kld ? key[44] : _0261_;
  assign _0262_ = ~rcon[13];
  assign _0263_ = ~wo_2[13];
  assign _0264_ = _0263_ ^ wo_0[13];
  assign _0265_ = _0264_ ^ wo_1[13];
  assign _0266_ = _0265_ ^ subword[13];
  assign _0267_ = _0266_ ^ _0262_;
  assign _0002_[13] = kld ? key[45] : _0267_;
  assign _0268_ = ~rcon[14];
  assign _0269_ = ~wo_2[14];
  assign _0270_ = _0269_ ^ wo_0[14];
  assign _0271_ = _0270_ ^ wo_1[14];
  assign _0272_ = _0271_ ^ subword[14];
  assign _0273_ = _0272_ ^ _0268_;
  assign _0002_[14] = kld ? key[46] : _0273_;
  assign _0274_ = ~rcon[15];
  assign _0275_ = ~wo_2[15];
  assign _0276_ = _0275_ ^ wo_0[15];
  assign _0277_ = _0276_ ^ wo_1[15];
  assign _0278_ = _0277_ ^ subword[15];
  assign _0279_ = _0278_ ^ _0274_;
  assign _0002_[15] = kld ? key[47] : _0279_;
  assign _0280_ = ~rcon[16];
  assign _0281_ = ~wo_2[16];
  assign _0282_ = _0281_ ^ wo_0[16];
  assign _0283_ = _0282_ ^ wo_1[16];
  assign _0284_ = _0283_ ^ subword[16];
  assign _0285_ = _0284_ ^ _0280_;
  assign _0002_[16] = kld ? key[48] : _0285_;
  assign _0286_ = ~rcon[17];
  assign _0287_ = ~wo_2[17];
  assign _0288_ = _0287_ ^ wo_0[17];
  assign _0289_ = _0288_ ^ wo_1[17];
  assign _0290_ = _0289_ ^ subword[17];
  assign _0291_ = _0290_ ^ _0286_;
  assign _0002_[17] = kld ? key[49] : _0291_;
  assign _0292_ = ~rcon[18];
  assign _0293_ = ~wo_2[18];
  assign _0294_ = _0293_ ^ wo_0[18];
  assign _0295_ = _0294_ ^ wo_1[18];
  assign _0296_ = _0295_ ^ subword[18];
  assign _0297_ = _0296_ ^ _0292_;
  assign _0002_[18] = kld ? key[50] : _0297_;
  assign _0298_ = ~rcon[19];
  assign _0299_ = ~wo_2[19];
  assign _0300_ = _0299_ ^ wo_0[19];
  assign _0301_ = _0300_ ^ wo_1[19];
  assign _0302_ = _0301_ ^ subword[19];
  assign _0303_ = _0302_ ^ _0298_;
  assign _0002_[19] = kld ? key[51] : _0303_;
  assign _0304_ = ~rcon[1];
  assign _0305_ = ~wo_2[1];
  assign _0306_ = _0305_ ^ wo_0[1];
  assign _0307_ = _0306_ ^ wo_1[1];
  assign _0308_ = _0307_ ^ subword[1];
  assign _0309_ = _0308_ ^ _0304_;
  assign _0002_[1] = kld ? key[33] : _0309_;
  assign _0310_ = ~rcon[20];
  assign _0311_ = ~wo_2[20];
  assign _0312_ = _0311_ ^ wo_0[20];
  assign _0313_ = _0312_ ^ wo_1[20];
  assign _0314_ = _0313_ ^ subword[20];
  assign _0315_ = _0314_ ^ _0310_;
  assign _0002_[20] = kld ? key[52] : _0315_;
  assign _0316_ = ~rcon[21];
  assign _0317_ = ~wo_2[21];
  assign _0318_ = _0317_ ^ wo_0[21];
  assign _0319_ = _0318_ ^ wo_1[21];
  assign _0320_ = _0319_ ^ subword[21];
  assign _0321_ = _0320_ ^ _0316_;
  assign _0002_[21] = kld ? key[53] : _0321_;
  assign _0322_ = ~rcon[22];
  assign _0323_ = ~wo_2[22];
  assign _0324_ = _0323_ ^ wo_0[22];
  assign _0325_ = _0324_ ^ wo_1[22];
  assign _0326_ = _0325_ ^ subword[22];
  assign _0327_ = _0326_ ^ _0322_;
  assign _0002_[22] = kld ? key[54] : _0327_;
  assign _0328_ = ~rcon[23];
  assign _0329_ = ~wo_2[23];
  assign _0330_ = _0329_ ^ wo_0[23];
  assign _0331_ = _0330_ ^ wo_1[23];
  assign _0332_ = _0331_ ^ subword[23];
  assign _0333_ = _0332_ ^ _0328_;
  assign _0002_[23] = kld ? key[55] : _0333_;
  assign _0334_ = ~rcon[24];
  assign _0335_ = ~wo_2[24];
  assign _0336_ = _0335_ ^ wo_0[24];
  assign _0337_ = _0336_ ^ wo_1[24];
  assign _0338_ = _0337_ ^ subword[24];
  assign _0339_ = _0338_ ^ _0334_;
  assign _0002_[24] = kld ? key[56] : _0339_;
  assign _0340_ = ~rcon[25];
  assign _0341_ = ~wo_2[25];
  assign _0342_ = _0341_ ^ wo_0[25];
  assign _0343_ = _0342_ ^ wo_1[25];
  assign _0344_ = _0343_ ^ subword[25];
  assign _0345_ = _0344_ ^ _0340_;
  assign _0002_[25] = kld ? key[57] : _0345_;
  assign _0346_ = ~rcon[26];
  assign _0347_ = ~wo_2[26];
  assign _0348_ = _0347_ ^ wo_0[26];
  assign _0349_ = _0348_ ^ wo_1[26];
  assign _0350_ = _0349_ ^ subword[26];
  assign _0351_ = _0350_ ^ _0346_;
  assign _0002_[26] = kld ? key[58] : _0351_;
  assign _0352_ = ~rcon[27];
  assign _0353_ = ~wo_2[27];
  assign _0354_ = _0353_ ^ wo_0[27];
  assign _0355_ = _0354_ ^ wo_1[27];
  assign _0356_ = _0355_ ^ subword[27];
  assign _0357_ = _0356_ ^ _0352_;
  assign _0002_[27] = kld ? key[59] : _0357_;
  assign _0358_ = ~rcon[28];
  assign _0359_ = ~wo_2[28];
  assign _0360_ = _0359_ ^ wo_0[28];
  assign _0361_ = _0360_ ^ wo_1[28];
  assign _0362_ = _0361_ ^ subword[28];
  assign _0363_ = _0362_ ^ _0358_;
  assign _0002_[28] = kld ? key[60] : _0363_;
  assign _0364_ = ~rcon[29];
  assign _0365_ = ~wo_2[29];
  assign _0366_ = _0365_ ^ wo_0[29];
  assign _0367_ = _0366_ ^ wo_1[29];
  assign _0368_ = _0367_ ^ subword[29];
  assign _0369_ = _0368_ ^ _0364_;
  assign _0002_[29] = kld ? key[61] : _0369_;
  assign _0370_ = ~rcon[2];
  assign _0371_ = ~wo_2[2];
  assign _0372_ = _0371_ ^ wo_0[2];
  assign _0373_ = _0372_ ^ wo_1[2];
  assign _0374_ = _0373_ ^ subword[2];
  assign _0375_ = _0374_ ^ _0370_;
  assign _0002_[2] = kld ? key[34] : _0375_;
  assign _0376_ = ~rcon[30];
  assign _0377_ = ~wo_2[30];
  assign _0378_ = _0377_ ^ wo_0[30];
  assign _0379_ = _0378_ ^ wo_1[30];
  assign _0380_ = _0379_ ^ subword[30];
  assign _0381_ = _0380_ ^ _0376_;
  assign _0002_[30] = kld ? key[62] : _0381_;
  assign _0382_ = ~rcon[31];
  assign _0383_ = ~wo_2[31];
  assign _0384_ = _0383_ ^ wo_0[31];
  assign _0385_ = _0384_ ^ wo_1[31];
  assign _0386_ = _0385_ ^ subword[31];
  assign _0387_ = _0386_ ^ _0382_;
  assign _0002_[31] = kld ? key[63] : _0387_;
  assign _0388_ = ~rcon[3];
  assign _0389_ = ~wo_2[3];
  assign _0390_ = _0389_ ^ wo_0[3];
  assign _0391_ = _0390_ ^ wo_1[3];
  assign _0392_ = _0391_ ^ subword[3];
  assign _0393_ = _0392_ ^ _0388_;
  assign _0002_[3] = kld ? key[35] : _0393_;
  assign _0394_ = ~rcon[4];
  assign _0395_ = ~wo_2[4];
  assign _0396_ = _0395_ ^ wo_0[4];
  assign _0397_ = _0396_ ^ wo_1[4];
  assign _0398_ = _0397_ ^ subword[4];
  assign _0399_ = _0398_ ^ _0394_;
  assign _0002_[4] = kld ? key[36] : _0399_;
  assign _0400_ = ~rcon[5];
  assign _0401_ = ~wo_2[5];
  assign _0402_ = _0401_ ^ wo_0[5];
  assign _0403_ = _0402_ ^ wo_1[5];
  assign _0404_ = _0403_ ^ subword[5];
  assign _0405_ = _0404_ ^ _0400_;
  assign _0002_[5] = kld ? key[37] : _0405_;
  assign _0406_ = ~rcon[6];
  assign _0407_ = ~wo_2[6];
  assign _0408_ = _0407_ ^ wo_0[6];
  assign _0409_ = _0408_ ^ wo_1[6];
  assign _0410_ = _0409_ ^ subword[6];
  assign _0411_ = _0410_ ^ _0406_;
  assign _0002_[6] = kld ? key[38] : _0411_;
  assign _0412_ = ~rcon[7];
  assign _0413_ = ~wo_2[7];
  assign _0414_ = _0413_ ^ wo_0[7];
  assign _0415_ = _0414_ ^ wo_1[7];
  assign _0416_ = _0415_ ^ subword[7];
  assign _0417_ = _0416_ ^ _0412_;
  assign _0002_[7] = kld ? key[39] : _0417_;
  assign _0418_ = ~rcon[8];
  assign _0419_ = ~wo_2[8];
  assign _0420_ = _0419_ ^ wo_0[8];
  assign _0421_ = _0420_ ^ wo_1[8];
  assign _0422_ = _0421_ ^ subword[8];
  assign _0423_ = _0422_ ^ _0418_;
  assign _0002_[8] = kld ? key[40] : _0423_;
  assign _0424_ = ~rcon[9];
  assign _0425_ = ~wo_2[9];
  assign _0426_ = _0425_ ^ wo_0[9];
  assign _0427_ = _0426_ ^ wo_1[9];
  assign _0428_ = _0427_ ^ subword[9];
  assign _0429_ = _0428_ ^ _0424_;
  assign _0002_[9] = kld ? key[41] : _0429_;
  assign _0430_ = tmp_w[0] ^ wo_0[0];
  assign _0431_ = _0430_ ^ _0239_;
  assign _0432_ = _0431_ ^ wo_1[0];
  assign _0433_ = _0432_ ^ subword[0];
  assign _0434_ = _0433_ ^ _0238_;
  assign _0003_[0] = kld ? key[0] : _0434_;
  assign _0435_ = tmp_w[10] ^ wo_0[10];
  assign _0436_ = _0435_ ^ _0245_;
  assign _0437_ = _0436_ ^ wo_1[10];
  assign _0438_ = _0437_ ^ subword[10];
  assign _0439_ = _0438_ ^ _0244_;
  assign _0003_[10] = kld ? key[10] : _0439_;
  assign _0440_ = tmp_w[11] ^ wo_0[11];
  assign _0441_ = _0440_ ^ _0251_;
  assign _0442_ = _0441_ ^ wo_1[11];
  assign _0443_ = _0442_ ^ subword[11];
  assign _0444_ = _0443_ ^ _0250_;
  assign _0003_[11] = kld ? key[11] : _0444_;
  assign _0445_ = tmp_w[12] ^ wo_0[12];
  assign _0446_ = _0445_ ^ _0257_;
  assign _0447_ = _0446_ ^ wo_1[12];
  assign _0448_ = _0447_ ^ subword[12];
  assign _0449_ = _0448_ ^ _0256_;
  assign _0003_[12] = kld ? key[12] : _0449_;
  assign _0450_ = tmp_w[13] ^ wo_0[13];
  assign _0451_ = _0450_ ^ _0263_;
  assign _0452_ = _0451_ ^ wo_1[13];
  assign _0453_ = _0452_ ^ subword[13];
  assign _0454_ = _0453_ ^ _0262_;
  assign _0003_[13] = kld ? key[13] : _0454_;
  assign _0455_ = tmp_w[14] ^ wo_0[14];
  assign _0456_ = _0455_ ^ _0269_;
  assign _0457_ = _0456_ ^ wo_1[14];
  assign _0458_ = _0457_ ^ subword[14];
  assign _0459_ = _0458_ ^ _0268_;
  assign _0003_[14] = kld ? key[14] : _0459_;
  assign _0460_ = tmp_w[15] ^ wo_0[15];
  assign _0461_ = _0460_ ^ _0275_;
  assign _0462_ = _0461_ ^ wo_1[15];
  assign _0463_ = _0462_ ^ subword[15];
  assign _0464_ = _0463_ ^ _0274_;
  assign _0003_[15] = kld ? key[15] : _0464_;
  assign _0465_ = tmp_w[16] ^ wo_0[16];
  assign _0466_ = _0465_ ^ _0281_;
  assign _0467_ = _0466_ ^ wo_1[16];
  assign _0468_ = _0467_ ^ subword[16];
  assign _0469_ = _0468_ ^ _0280_;
  assign _0003_[16] = kld ? key[16] : _0469_;
  assign _0470_ = tmp_w[17] ^ wo_0[17];
  assign _0471_ = _0470_ ^ _0287_;
  assign _0472_ = _0471_ ^ wo_1[17];
  assign _0473_ = _0472_ ^ subword[17];
  assign _0474_ = _0473_ ^ _0286_;
  assign _0003_[17] = kld ? key[17] : _0474_;
  assign _0475_ = tmp_w[18] ^ wo_0[18];
  assign _0476_ = _0475_ ^ _0293_;
  assign _0477_ = _0476_ ^ wo_1[18];
  assign _0478_ = _0477_ ^ subword[18];
  assign _0479_ = _0478_ ^ _0292_;
  assign _0003_[18] = kld ? key[18] : _0479_;
  assign _0480_ = tmp_w[19] ^ wo_0[19];
  assign _0481_ = _0480_ ^ _0299_;
  assign _0482_ = _0481_ ^ wo_1[19];
  assign _0483_ = _0482_ ^ subword[19];
  assign _0484_ = _0483_ ^ _0298_;
  assign _0003_[19] = kld ? key[19] : _0484_;
  assign _0485_ = tmp_w[1] ^ wo_0[1];
  assign _0486_ = _0485_ ^ _0305_;
  assign _0487_ = _0486_ ^ wo_1[1];
  assign _0488_ = _0487_ ^ subword[1];
  assign _0489_ = _0488_ ^ _0304_;
  assign _0003_[1] = kld ? key[1] : _0489_;
  assign _0490_ = tmp_w[20] ^ wo_0[20];
  assign _0491_ = _0490_ ^ _0311_;
  assign _0492_ = _0491_ ^ wo_1[20];
  assign _0493_ = _0492_ ^ subword[20];
  assign _0494_ = _0493_ ^ _0310_;
  assign _0003_[20] = kld ? key[20] : _0494_;
  assign _0495_ = tmp_w[21] ^ wo_0[21];
  assign _0496_ = _0495_ ^ _0317_;
  assign _0497_ = _0496_ ^ wo_1[21];
  assign _0498_ = _0497_ ^ subword[21];
  assign _0499_ = _0498_ ^ _0316_;
  assign _0003_[21] = kld ? key[21] : _0499_;
  assign _0500_ = tmp_w[22] ^ wo_0[22];
  assign _0501_ = _0500_ ^ _0323_;
  assign _0502_ = _0501_ ^ wo_1[22];
  assign _0503_ = _0502_ ^ subword[22];
  assign _0504_ = _0503_ ^ _0322_;
  assign _0003_[22] = kld ? key[22] : _0504_;
  assign _0505_ = tmp_w[23] ^ wo_0[23];
  assign _0506_ = _0505_ ^ _0329_;
  assign _0507_ = _0506_ ^ wo_1[23];
  assign _0508_ = _0507_ ^ subword[23];
  assign _0509_ = _0508_ ^ _0328_;
  assign _0003_[23] = kld ? key[23] : _0509_;
  assign _0510_ = tmp_w[24] ^ wo_0[24];
  assign _0511_ = _0510_ ^ _0335_;
  assign _0512_ = _0511_ ^ wo_1[24];
  assign _0513_ = _0512_ ^ subword[24];
  assign _0514_ = _0513_ ^ _0334_;
  assign _0003_[24] = kld ? key[24] : _0514_;
  assign _0515_ = tmp_w[25] ^ wo_0[25];
  assign _0004_ = _0515_ ^ _0341_;
  assign _0005_ = _0004_ ^ wo_1[25];
  assign _0006_ = _0005_ ^ subword[25];
  assign _0007_ = _0006_ ^ _0340_;
  assign _0003_[25] = kld ? key[25] : _0007_;
  assign _0008_ = tmp_w[26] ^ wo_0[26];
  assign _0009_ = _0008_ ^ _0347_;
  assign _0010_ = _0009_ ^ wo_1[26];
  assign _0011_ = _0010_ ^ subword[26];
  assign _0012_ = _0011_ ^ _0346_;
  assign _0003_[26] = kld ? key[26] : _0012_;
  assign _0013_ = tmp_w[27] ^ wo_0[27];
  assign _0014_ = _0013_ ^ _0353_;
  assign _0015_ = _0014_ ^ wo_1[27];
  assign _0016_ = _0015_ ^ subword[27];
  assign _0017_ = _0016_ ^ _0352_;
  assign _0003_[27] = kld ? key[27] : _0017_;
  assign _0018_ = tmp_w[28] ^ wo_0[28];
  assign _0019_ = _0018_ ^ _0359_;
  assign _0020_ = _0019_ ^ wo_1[28];
  assign _0021_ = _0020_ ^ subword[28];
  assign _0022_ = _0021_ ^ _0358_;
  assign _0003_[28] = kld ? key[28] : _0022_;
  assign _0023_ = tmp_w[29] ^ wo_0[29];
  assign _0024_ = _0023_ ^ _0365_;
  assign _0025_ = _0024_ ^ wo_1[29];
  assign _0026_ = _0025_ ^ subword[29];
  assign _0027_ = _0026_ ^ _0364_;
  assign _0003_[29] = kld ? key[29] : _0027_;
  assign _0028_ = tmp_w[2] ^ wo_0[2];
  assign _0029_ = _0028_ ^ _0371_;
  assign _0030_ = _0029_ ^ wo_1[2];
  assign _0031_ = _0030_ ^ subword[2];
  assign _0032_ = _0031_ ^ _0370_;
  assign _0003_[2] = kld ? key[2] : _0032_;
  assign _0033_ = tmp_w[30] ^ wo_0[30];
  assign _0034_ = _0033_ ^ _0377_;
  assign _0035_ = _0034_ ^ wo_1[30];
  assign _0036_ = _0035_ ^ subword[30];
  assign _0037_ = _0036_ ^ _0376_;
  assign _0003_[30] = kld ? key[30] : _0037_;
  assign _0038_ = tmp_w[31] ^ wo_0[31];
  assign _0039_ = _0038_ ^ _0383_;
  assign _0040_ = _0039_ ^ wo_1[31];
  assign _0041_ = _0040_ ^ subword[31];
  assign _0042_ = _0041_ ^ _0382_;
  assign _0003_[31] = kld ? key[31] : _0042_;
  assign _0043_ = tmp_w[3] ^ wo_0[3];
  assign _0044_ = _0043_ ^ _0389_;
  assign _0045_ = _0044_ ^ wo_1[3];
  assign _0046_ = _0045_ ^ subword[3];
  assign _0047_ = _0046_ ^ _0388_;
  assign _0003_[3] = kld ? key[3] : _0047_;
  assign _0048_ = tmp_w[4] ^ wo_0[4];
  assign _0049_ = _0048_ ^ _0395_;
  assign _0050_ = _0049_ ^ wo_1[4];
  assign _0051_ = _0050_ ^ subword[4];
  assign _0052_ = _0051_ ^ _0394_;
  assign _0003_[4] = kld ? key[4] : _0052_;
  assign _0053_ = tmp_w[5] ^ wo_0[5];
  assign _0054_ = _0053_ ^ _0401_;
  assign _0055_ = _0054_ ^ wo_1[5];
  assign _0056_ = _0055_ ^ subword[5];
  assign _0057_ = _0056_ ^ _0400_;
  assign _0003_[5] = kld ? key[5] : _0057_;
  assign _0058_ = tmp_w[6] ^ wo_0[6];
  assign _0059_ = _0058_ ^ _0407_;
  assign _0060_ = _0059_ ^ wo_1[6];
  assign _0061_ = _0060_ ^ subword[6];
  assign _0062_ = _0061_ ^ _0406_;
  assign _0003_[6] = kld ? key[6] : _0062_;
  assign _0063_ = tmp_w[7] ^ wo_0[7];
  assign _0064_ = _0063_ ^ _0413_;
  assign _0065_ = _0064_ ^ wo_1[7];
  assign _0066_ = _0065_ ^ subword[7];
  assign _0067_ = _0066_ ^ _0412_;
  assign _0003_[7] = kld ? key[7] : _0067_;
  assign _0068_ = tmp_w[8] ^ wo_0[8];
  assign _0069_ = _0068_ ^ _0419_;
  assign _0070_ = _0069_ ^ wo_1[8];
  assign _0071_ = _0070_ ^ subword[8];
  assign _0072_ = _0071_ ^ _0418_;
  assign _0003_[8] = kld ? key[8] : _0072_;
  assign _0073_ = tmp_w[9] ^ wo_0[9];
  assign _0074_ = _0073_ ^ _0425_;
  assign _0075_ = _0074_ ^ wo_1[9];
  assign _0076_ = _0075_ ^ subword[9];
  assign _0077_ = _0076_ ^ _0424_;
  assign _0003_[9] = kld ? key[9] : _0077_;
  always @(posedge clk)
      wo_0[0] <= _0000_[0];
  always @(posedge clk)
      wo_0[10] <= _0000_[10];
  always @(posedge clk)
      wo_0[11] <= _0000_[11];
  always @(posedge clk)
      wo_0[12] <= _0000_[12];
  always @(posedge clk)
      wo_0[13] <= _0000_[13];
  always @(posedge clk)
      wo_0[14] <= _0000_[14];
  always @(posedge clk)
      wo_0[15] <= _0000_[15];
  always @(posedge clk)
      wo_0[16] <= _0000_[16];
  always @(posedge clk)
      wo_0[17] <= _0000_[17];
  always @(posedge clk)
      wo_0[18] <= _0000_[18];
  always @(posedge clk)
      wo_0[19] <= _0000_[19];
  always @(posedge clk)
      wo_0[1] <= _0000_[1];
  always @(posedge clk)
      wo_0[20] <= _0000_[20];
  always @(posedge clk)
      wo_0[21] <= _0000_[21];
  always @(posedge clk)
      wo_0[22] <= _0000_[22];
  always @(posedge clk)
      wo_0[23] <= _0000_[23];
  always @(posedge clk)
      wo_0[24] <= _0000_[24];
  always @(posedge clk)
      wo_0[25] <= _0000_[25];
  always @(posedge clk)
      wo_0[26] <= _0000_[26];
  always @(posedge clk)
      wo_0[27] <= _0000_[27];
  always @(posedge clk)
      wo_0[28] <= _0000_[28];
  always @(posedge clk)
      wo_0[29] <= _0000_[29];
  always @(posedge clk)
      wo_0[2] <= _0000_[2];
  always @(posedge clk)
      wo_0[30] <= _0000_[30];
  always @(posedge clk)
      wo_0[31] <= _0000_[31];
  always @(posedge clk)
      wo_0[3] <= _0000_[3];
  always @(posedge clk)
      wo_0[4] <= _0000_[4];
  always @(posedge clk)
      wo_0[5] <= _0000_[5];
  always @(posedge clk)
      wo_0[6] <= _0000_[6];
  always @(posedge clk)
      wo_0[7] <= _0000_[7];
  always @(posedge clk)
      wo_0[8] <= _0000_[8];
  always @(posedge clk)
      wo_0[9] <= _0000_[9];
  always @(posedge clk)
      wo_1[0] <= _0001_[0];
  always @(posedge clk)
      wo_1[10] <= _0001_[10];
  always @(posedge clk)
      wo_1[11] <= _0001_[11];
  always @(posedge clk)
      wo_1[12] <= _0001_[12];
  always @(posedge clk)
      wo_1[13] <= _0001_[13];
  always @(posedge clk)
      wo_1[14] <= _0001_[14];
  always @(posedge clk)
      wo_1[15] <= _0001_[15];
  always @(posedge clk)
      wo_1[16] <= _0001_[16];
  always @(posedge clk)
      wo_1[17] <= _0001_[17];
  always @(posedge clk)
      wo_1[18] <= _0001_[18];
  always @(posedge clk)
      wo_1[19] <= _0001_[19];
  always @(posedge clk)
      wo_1[1] <= _0001_[1];
  always @(posedge clk)
      wo_1[20] <= _0001_[20];
  always @(posedge clk)
      wo_1[21] <= _0001_[21];
  always @(posedge clk)
      wo_1[22] <= _0001_[22];
  always @(posedge clk)
      wo_1[23] <= _0001_[23];
  always @(posedge clk)
      wo_1[24] <= _0001_[24];
  always @(posedge clk)
      wo_1[25] <= _0001_[25];
  always @(posedge clk)
      wo_1[26] <= _0001_[26];
  always @(posedge clk)
      wo_1[27] <= _0001_[27];
  always @(posedge clk)
      wo_1[28] <= _0001_[28];
  always @(posedge clk)
      wo_1[29] <= _0001_[29];
  always @(posedge clk)
      wo_1[2] <= _0001_[2];
  always @(posedge clk)
      wo_1[30] <= _0001_[30];
  always @(posedge clk)
      wo_1[31] <= _0001_[31];
  always @(posedge clk)
      wo_1[3] <= _0001_[3];
  always @(posedge clk)
      wo_1[4] <= _0001_[4];
  always @(posedge clk)
      wo_1[5] <= _0001_[5];
  always @(posedge clk)
      wo_1[6] <= _0001_[6];
  always @(posedge clk)
      wo_1[7] <= _0001_[7];
  always @(posedge clk)
      wo_1[8] <= _0001_[8];
  always @(posedge clk)
      wo_1[9] <= _0001_[9];
  always @(posedge clk)
      wo_2[0] <= _0002_[0];
  always @(posedge clk)
      wo_2[10] <= _0002_[10];
  always @(posedge clk)
      wo_2[11] <= _0002_[11];
  always @(posedge clk)
      wo_2[12] <= _0002_[12];
  always @(posedge clk)
      wo_2[13] <= _0002_[13];
  always @(posedge clk)
      wo_2[14] <= _0002_[14];
  always @(posedge clk)
      wo_2[15] <= _0002_[15];
  always @(posedge clk)
      wo_2[16] <= _0002_[16];
  always @(posedge clk)
      wo_2[17] <= _0002_[17];
  always @(posedge clk)
      wo_2[18] <= _0002_[18];
  always @(posedge clk)
      wo_2[19] <= _0002_[19];
  always @(posedge clk)
      wo_2[1] <= _0002_[1];
  always @(posedge clk)
      wo_2[20] <= _0002_[20];
  always @(posedge clk)
      wo_2[21] <= _0002_[21];
  always @(posedge clk)
      wo_2[22] <= _0002_[22];
  always @(posedge clk)
      wo_2[23] <= _0002_[23];
  always @(posedge clk)
      wo_2[24] <= _0002_[24];
  always @(posedge clk)
      wo_2[25] <= _0002_[25];
  always @(posedge clk)
      wo_2[26] <= _0002_[26];
  always @(posedge clk)
      wo_2[27] <= _0002_[27];
  always @(posedge clk)
      wo_2[28] <= _0002_[28];
  always @(posedge clk)
      wo_2[29] <= _0002_[29];
  always @(posedge clk)
      wo_2[2] <= _0002_[2];
  always @(posedge clk)
      wo_2[30] <= _0002_[30];
  always @(posedge clk)
      wo_2[31] <= _0002_[31];
  always @(posedge clk)
      wo_2[3] <= _0002_[3];
  always @(posedge clk)
      wo_2[4] <= _0002_[4];
  always @(posedge clk)
      wo_2[5] <= _0002_[5];
  always @(posedge clk)
      wo_2[6] <= _0002_[6];
  always @(posedge clk)
      wo_2[7] <= _0002_[7];
  always @(posedge clk)
      wo_2[8] <= _0002_[8];
  always @(posedge clk)
      wo_2[9] <= _0002_[9];
  always @(posedge clk)
      tmp_w[0] <= _0003_[0];
  always @(posedge clk)
      tmp_w[10] <= _0003_[10];
  always @(posedge clk)
      tmp_w[11] <= _0003_[11];
  always @(posedge clk)
      tmp_w[12] <= _0003_[12];
  always @(posedge clk)
      tmp_w[13] <= _0003_[13];
  always @(posedge clk)
      tmp_w[14] <= _0003_[14];
  always @(posedge clk)
      tmp_w[15] <= _0003_[15];
  always @(posedge clk)
      tmp_w[16] <= _0003_[16];
  always @(posedge clk)
      tmp_w[17] <= _0003_[17];
  always @(posedge clk)
      tmp_w[18] <= _0003_[18];
  always @(posedge clk)
      tmp_w[19] <= _0003_[19];
  always @(posedge clk)
      tmp_w[1] <= _0003_[1];
  always @(posedge clk)
      tmp_w[20] <= _0003_[20];
  always @(posedge clk)
      tmp_w[21] <= _0003_[21];
  always @(posedge clk)
      tmp_w[22] <= _0003_[22];
  always @(posedge clk)
      tmp_w[23] <= _0003_[23];
  always @(posedge clk)
      tmp_w[24] <= _0003_[24];
  always @(posedge clk)
      tmp_w[25] <= _0003_[25];
  always @(posedge clk)
      tmp_w[26] <= _0003_[26];
  always @(posedge clk)
      tmp_w[27] <= _0003_[27];
  always @(posedge clk)
      tmp_w[28] <= _0003_[28];
  always @(posedge clk)
      tmp_w[29] <= _0003_[29];
  always @(posedge clk)
      tmp_w[2] <= _0003_[2];
  always @(posedge clk)
      tmp_w[30] <= _0003_[30];
  always @(posedge clk)
      tmp_w[31] <= _0003_[31];
  always @(posedge clk)
      tmp_w[3] <= _0003_[3];
  always @(posedge clk)
      tmp_w[4] <= _0003_[4];
  always @(posedge clk)
      tmp_w[5] <= _0003_[5];
  always @(posedge clk)
      tmp_w[6] <= _0003_[6];
  always @(posedge clk)
      tmp_w[7] <= _0003_[7];
  always @(posedge clk)
      tmp_w[8] <= _0003_[8];
  always @(posedge clk)
      tmp_w[9] <= _0003_[9];
  aes_rcon r0 (
    .clk(clk),
    .kld(kld),
    .out(rcon)
  );
  aes_sbox u0 (
    .a(tmp_w[23:16]),
    .d(subword[31:24])
  );
  aes_sbox u1 (
    .a(tmp_w[15:8]),
    .d(subword[23:16])
  );
  aes_sbox u2 (
    .a(tmp_w[7:0]),
    .d(subword[15:8])
  );
  aes_sbox u3 (
    .a(tmp_w[31:24]),
    .d(subword[7:0])
  );
  assign wo_3 = tmp_w;
endmodule

module aes_rcon(clk, kld, out);
  wire [31:0] _000_;
  wire [3:0] _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  input clk;
  input kld;
  output [31:0] out;
  reg [3:0] rcnt;
  assign _002_ = ~rcnt[3];
  assign _003_ = rcnt[1] & rcnt[0];
  assign _004_ = _003_ & rcnt[2];
  assign _005_ = _004_ ^ _002_;
  assign _006_ = _003_ ^ rcnt[2];
  assign _007_ = _003_ & _006_;
  assign _008_ = _007_ & _005_;
  assign _009_ = ~rcnt[0];
  assign _010_ = ~rcnt[1];
  assign _011_ = _010_ & _009_;
  assign _012_ = _011_ & _006_;
  assign _013_ = _012_ & _005_;
  assign _014_ = _013_ | _008_;
  assign _015_ = _010_ & rcnt[0];
  assign _016_ = _015_ & _006_;
  assign _017_ = _016_ & _005_;
  assign _018_ = rcnt[1] & _009_;
  assign _019_ = _018_ & _006_;
  assign _020_ = _019_ & _005_;
  assign _021_ = _020_ | _017_;
  assign _022_ = _021_ | _014_;
  assign _023_ = _004_ ^ rcnt[3];
  assign _024_ = ~rcnt[2];
  assign _025_ = _003_ ^ _024_;
  assign _026_ = _004_ & _023_;
  assign _027_ = _011_ & _025_;
  assign _028_ = _027_ & _023_;
  assign _029_ = _028_ | _026_;
  assign _030_ = _004_ & _005_;
  assign _031_ = _027_ & _005_;
  assign _032_ = _031_ | _030_;
  assign _033_ = _015_ & _025_;
  assign _034_ = _033_ & _005_;
  assign _035_ = _018_ & _025_;
  assign _036_ = _035_ & _005_;
  assign _037_ = _036_ | _034_;
  assign _038_ = _037_ | _032_;
  assign _039_ = _038_ | _029_;
  assign _040_ = _039_ | _022_;
  assign _041_ = ~kld;
  assign _042_ = _004_ & _041_;
  assign _000_[24] = _042_ | kld;
  assign _043_ = _031_ | _029_;
  assign _044_ = _043_ & _041_;
  assign _000_[25] = _044_ & _040_;
  assign _045_ = _005_ ? _033_ : _027_;
  assign _046_ = _045_ & _041_;
  assign _000_[26] = _046_ & _040_;
  assign _047_ = _023_ ? _004_ : _035_;
  assign _048_ = _047_ & _041_;
  assign _000_[27] = _048_ & _040_;
  assign _049_ = _029_ | _008_;
  assign _050_ = _049_ & _041_;
  assign _000_[28] = _050_ & _040_;
  assign _051_ = _005_ ? _012_ : _027_;
  assign _052_ = _051_ & _041_;
  assign _000_[29] = _052_ & _040_;
  assign _053_ = _017_ & _041_;
  assign _000_[30] = _053_ & _040_;
  assign _054_ = _020_ & _041_;
  assign _000_[31] = _054_ & _040_;
  assign _001_[0] = _041_ & _009_;
  assign _055_ = rcnt[1] ^ rcnt[0];
  assign _001_[1] = _055_ & _041_;
  assign _001_[2] = _006_ & _041_;
  assign _001_[3] = _023_ & _041_;
  reg #~@out_reg[24]#~@;
  always @(posedge clk)
      #~@out_reg[24] #~@<= _000_[24];
  assign out[24] = #~@out_reg[24]#~@;
  reg #~@out_reg[25]#~@;
  always @(posedge clk)
      #~@out_reg[25] #~@<= _000_[25];
  assign out[25] = #~@out_reg[25]#~@;
  reg #~@out_reg[26]#~@;
  always @(posedge clk)
      #~@out_reg[26] #~@<= _000_[26];
  assign out[26] = #~@out_reg[26]#~@;
  reg #~@out_reg[27]#~@;
  always @(posedge clk)
      #~@out_reg[27] #~@<= _000_[27];
  assign out[27] = #~@out_reg[27]#~@;
  reg #~@out_reg[28]#~@;
  always @(posedge clk)
      #~@out_reg[28] #~@<= _000_[28];
  assign out[28] = #~@out_reg[28]#~@;
  reg #~@out_reg[29]#~@;
  always @(posedge clk)
      #~@out_reg[29] #~@<= _000_[29];
  assign out[29] = #~@out_reg[29]#~@;
  reg #~@out_reg[30]#~@;
  always @(posedge clk)
      #~@out_reg[30] #~@<= _000_[30];
  assign out[30] = #~@out_reg[30]#~@;
  reg #~@out_reg[31]#~@;
  always @(posedge clk)
      #~@out_reg[31] #~@<= _000_[31];
  assign out[31] = #~@out_reg[31]#~@;
  always @(posedge clk)
      rcnt[0] <= _001_[0];
  always @(posedge clk)
      rcnt[1] <= _001_[1];
  always @(posedge clk)
      rcnt[2] <= _001_[2];
  always @(posedge clk)
      rcnt[3] <= _001_[3];
  assign out[23:0] = 24'b000000000000000000000000;
endmodule

module aes_sbox(a, d);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire _1892_;
  wire _1893_;
  wire _1894_;
  wire _1895_;
  wire _1896_;
  wire _1897_;
  wire _1898_;
  wire _1899_;
  wire _1900_;
  wire _1901_;
  wire _1902_;
  wire _1903_;
  wire _1904_;
  wire _1905_;
  wire _1906_;
  wire _1907_;
  wire _1908_;
  wire _1909_;
  wire _1910_;
  wire _1911_;
  wire _1912_;
  wire _1913_;
  wire _1914_;
  wire _1915_;
  wire _1916_;
  wire _1917_;
  wire _1918_;
  wire _1919_;
  wire _1920_;
  wire _1921_;
  wire _1922_;
  wire _1923_;
  wire _1924_;
  wire _1925_;
  wire _1926_;
  wire _1927_;
  wire _1928_;
  wire _1929_;
  wire _1930_;
  wire _1931_;
  wire _1932_;
  wire _1933_;
  wire _1934_;
  wire _1935_;
  wire _1936_;
  wire _1937_;
  wire _1938_;
  wire _1939_;
  wire _1940_;
  wire _1941_;
  wire _1942_;
  wire _1943_;
  wire _1944_;
  wire _1945_;
  wire _1946_;
  wire _1947_;
  wire _1948_;
  wire _1949_;
  wire _1950_;
  wire _1951_;
  wire _1952_;
  wire _1953_;
  wire _1954_;
  wire _1955_;
  wire _1956_;
  wire _1957_;
  wire _1958_;
  wire _1959_;
  wire _1960_;
  wire _1961_;
  wire _1962_;
  wire _1963_;
  wire _1964_;
  wire _1965_;
  wire _1966_;
  wire _1967_;
  wire _1968_;
  wire _1969_;
  wire _1970_;
  wire _1971_;
  wire _1972_;
  wire _1973_;
  wire _1974_;
  wire _1975_;
  wire _1976_;
  wire _1977_;
  wire _1978_;
  wire _1979_;
  wire _1980_;
  wire _1981_;
  wire _1982_;
  wire _1983_;
  wire _1984_;
  wire _1985_;
  wire _1986_;
  wire _1987_;
  wire _1988_;
  wire _1989_;
  wire _1990_;
  wire _1991_;
  wire _1992_;
  wire _1993_;
  wire _1994_;
  wire _1995_;
  wire _1996_;
  wire _1997_;
  wire _1998_;
  wire _1999_;
  wire _2000_;
  wire _2001_;
  wire _2002_;
  wire _2003_;
  wire _2004_;
  wire _2005_;
  wire _2006_;
  wire _2007_;
  wire _2008_;
  wire _2009_;
  wire _2010_;
  wire _2011_;
  wire _2012_;
  wire _2013_;
  wire _2014_;
  wire _2015_;
  wire _2016_;
  wire _2017_;
  wire _2018_;
  wire _2019_;
  wire _2020_;
  wire _2021_;
  wire _2022_;
  wire _2023_;
  wire _2024_;
  wire _2025_;
  wire _2026_;
  wire _2027_;
  wire _2028_;
  wire _2029_;
  wire _2030_;
  wire _2031_;
  wire _2032_;
  wire _2033_;
  wire _2034_;
  wire _2035_;
  wire _2036_;
  wire _2037_;
  wire _2038_;
  wire _2039_;
  wire _2040_;
  wire _2041_;
  wire _2042_;
  wire _2043_;
  wire _2044_;
  wire _2045_;
  wire _2046_;
  wire _2047_;
  wire _2048_;
  wire _2049_;
  wire _2050_;
  wire _2051_;
  wire _2052_;
  wire _2053_;
  wire _2054_;
  wire _2055_;
  wire _2056_;
  wire _2057_;
  wire _2058_;
  wire _2059_;
  wire _2060_;
  wire _2061_;
  wire _2062_;
  wire _2063_;
  wire _2064_;
  wire _2065_;
  wire _2066_;
  wire _2067_;
  wire _2068_;
  wire _2069_;
  wire _2070_;
  wire _2071_;
  wire _2072_;
  wire _2073_;
  wire _2074_;
  wire _2075_;
  wire _2076_;
  wire _2077_;
  wire _2078_;
  wire _2079_;
  wire _2080_;
  wire _2081_;
  wire _2082_;
  wire _2083_;
  wire _2084_;
  wire _2085_;
  wire _2086_;
  wire _2087_;
  wire _2088_;
  wire _2089_;
  wire _2090_;
  wire _2091_;
  wire _2092_;
  wire _2093_;
  wire _2094_;
  wire _2095_;
  wire _2096_;
  wire _2097_;
  wire _2098_;
  wire _2099_;
  wire _2100_;
  wire _2101_;
  wire _2102_;
  wire _2103_;
  wire _2104_;
  wire _2105_;
  wire _2106_;
  wire _2107_;
  wire _2108_;
  wire _2109_;
  wire _2110_;
  wire _2111_;
  wire _2112_;
  wire _2113_;
  wire _2114_;
  wire _2115_;
  wire _2116_;
  wire _2117_;
  wire _2118_;
  wire _2119_;
  wire _2120_;
  wire _2121_;
  wire _2122_;
  wire _2123_;
  wire _2124_;
  wire _2125_;
  wire _2126_;
  wire _2127_;
  wire _2128_;
  wire _2129_;
  wire _2130_;
  wire _2131_;
  wire _2132_;
  wire _2133_;
  wire _2134_;
  wire _2135_;
  wire _2136_;
  wire _2137_;
  wire _2138_;
  wire _2139_;
  wire _2140_;
  wire _2141_;
  wire _2142_;
  wire _2143_;
  wire _2144_;
  wire _2145_;
  wire _2146_;
  wire _2147_;
  wire _2148_;
  wire _2149_;
  wire _2150_;
  wire _2151_;
  wire _2152_;
  wire _2153_;
  wire _2154_;
  wire _2155_;
  wire _2156_;
  wire _2157_;
  wire _2158_;
  wire _2159_;
  wire _2160_;
  wire _2161_;
  wire _2162_;
  wire _2163_;
  wire _2164_;
  wire _2165_;
  wire _2166_;
  wire _2167_;
  wire _2168_;
  wire _2169_;
  wire _2170_;
  wire _2171_;
  wire _2172_;
  wire _2173_;
  wire _2174_;
  wire _2175_;
  wire _2176_;
  wire _2177_;
  wire _2178_;
  wire _2179_;
  wire _2180_;
  wire _2181_;
  wire _2182_;
  wire _2183_;
  wire _2184_;
  wire _2185_;
  wire _2186_;
  wire _2187_;
  wire _2188_;
  wire _2189_;
  wire _2190_;
  wire _2191_;
  wire _2192_;
  wire _2193_;
  wire _2194_;
  wire _2195_;
  wire _2196_;
  wire _2197_;
  wire _2198_;
  wire _2199_;
  wire _2200_;
  wire _2201_;
  wire _2202_;
  wire _2203_;
  wire _2204_;
  wire _2205_;
  wire _2206_;
  wire _2207_;
  wire _2208_;
  wire _2209_;
  wire _2210_;
  wire _2211_;
  wire _2212_;
  wire _2213_;
  input [7:0] a;
  output [7:0] d;
  assign _0654_ = ~a[7];
  assign _0762_ = ~a[5];
  assign _0872_ = ~a[3];
  assign _0982_ = ~a[2];
  assign _1091_ = a[1] & a[0];
  assign _1198_ = _1091_ & _0982_;
  assign _1307_ = _1198_ & _0872_;
  assign _1416_ = _1307_ & a[4];
  assign _1445_ = _1416_ & _0762_;
  assign _1453_ = _1445_ & a[6];
  assign _1463_ = _1453_ & _0654_;
  assign _1474_ = ~a[0];
  assign _1482_ = ~a[1];
  assign _1490_ = _1482_ & _1474_;
  assign _1501_ = _1490_ & a[2];
  assign _1510_ = _1501_ & _0872_;
  assign _1520_ = _1510_ & a[4];
  assign _1530_ = _1520_ & _0762_;
  assign _1535_ = _1530_ & a[6];
  assign _1543_ = _1535_ & _0654_;
  assign _1561_ = _1482_ & a[0];
  assign _1570_ = _1561_ & a[2];
  assign _1579_ = _1570_ & _0872_;
  assign _1590_ = _1579_ & a[4];
  assign _1601_ = _1590_ & _0762_;
  assign _1611_ = _1601_ & a[6];
  assign _1621_ = _1611_ & _0654_;
  assign _1627_ = a[1] & _1474_;
  assign _1636_ = _1627_ & a[2];
  assign _1645_ = _1636_ & _0872_;
  assign _1656_ = _1645_ & a[4];
  assign _1664_ = _1656_ & _0762_;
  assign _1674_ = _1664_ & a[6];
  assign _1684_ = _1674_ & _0654_;
  assign _1705_ = ~a[4];
  assign _1715_ = _1091_ & a[2];
  assign _1726_ = _1715_ & a[3];
  assign _1737_ = _1726_ & _1705_;
  assign _1748_ = _1737_ & _0762_;
  assign _1759_ = _1748_ & a[6];
  assign _1770_ = _1759_ & _0654_;
  assign _1781_ = _1490_ & _0982_;
  assign _1792_ = _1781_ & _0872_;
  assign _1803_ = _1792_ & a[4];
  assign _1814_ = _1803_ & _0762_;
  assign _1825_ = _1814_ & a[6];
  assign _1836_ = _1825_ & _0654_;
  assign _1857_ = _1561_ & _0982_;
  assign _1868_ = _1857_ & _0872_;
  assign _1879_ = _1868_ & a[4];
  assign _1890_ = _1879_ & _0762_;
  assign _1901_ = _1890_ & a[6];
  assign _1912_ = _1901_ & _0654_;
  assign _1923_ = _1627_ & _0982_;
  assign _1934_ = _1923_ & _0872_;
  assign _1945_ = _1934_ & a[4];
  assign _1956_ = _1945_ & _0762_;
  assign _1967_ = _1956_ & a[6];
  assign _2018_ = _1198_ & a[3];
  assign _2029_ = _2018_ & a[4];
  assign _2040_ = _2029_ & _0762_;
  assign _2051_ = _2040_ & a[6];
  assign _2062_ = _2051_ & _0654_;
  assign _2073_ = _1501_ & a[3];
  assign _2084_ = _2073_ & a[4];
  assign _2095_ = _2084_ & _0762_;
  assign _2105_ = _2095_ & a[6];
  assign _2116_ = _2105_ & _0654_;
  assign _2137_ = _1570_ & a[3];
  assign _2148_ = _2137_ & a[4];
  assign _2159_ = _2148_ & _0762_;
  assign _2170_ = _2159_ & a[6];
  assign _2181_ = _2170_ & _0654_;
  assign _2192_ = _1636_ & a[3];
  assign _2203_ = _2192_ & a[4];
  assign _0000_ = _2203_ & _0762_;
  assign _0011_ = _0000_ & a[6];
  assign _0022_ = _0011_ & _0654_;
  assign _0033_ = _0022_ | _2181_;
  assign _0054_ = _1715_ & _0872_;
  assign _0065_ = _0054_ & a[4];
  assign _0076_ = _0065_ & _0762_;
  assign _0087_ = _0076_ & a[6];
  assign _0098_ = _0087_ & _0654_;
  assign _0109_ = _1781_ & a[3];
  assign _0120_ = _0109_ & a[4];
  assign _0131_ = _0120_ & _0762_;
  assign _0142_ = _0131_ & a[6];
  assign _0153_ = _0142_ & _0654_;
  assign _0164_ = _0153_ | _0098_;
  assign _0175_ = _1857_ & a[3];
  assign _0186_ = _0175_ & a[4];
  assign _0197_ = _0186_ & _0762_;
  assign _0208_ = _0197_ & a[6];
  assign _0219_ = _0208_ & _0654_;
  assign _0230_ = _1923_ & a[3];
  assign _0241_ = _0230_ & a[4];
  assign _0252_ = _0241_ & _0762_;
  assign _0263_ = _0252_ & a[6];
  assign _0274_ = _0263_ & _0654_;
  assign _0325_ = _1307_ & _1705_;
  assign _0336_ = _0325_ & _0762_;
  assign _0347_ = _0336_ & a[6];
  assign _0358_ = _0347_ & _0654_;
  assign _0369_ = _1510_ & _1705_;
  assign _0380_ = _0369_ & _0762_;
  assign _0391_ = _0380_ & a[6];
  assign _0402_ = _0391_ & _0654_;
  assign _0413_ = _0402_ | _0358_;
  assign _0424_ = _1579_ & _1705_;
  assign _0435_ = _0424_ & _0762_;
  assign _0446_ = _0435_ & a[6];
  assign _0457_ = _0446_ & _0654_;
  assign _0468_ = _1645_ & _1705_;
  assign _0479_ = _0468_ & _0762_;
  assign _0490_ = _0479_ & a[6];
  assign _0501_ = _0490_ & _0654_;
  assign _0512_ = _0501_ | _0457_;
  assign _0523_ = _0512_ | _0413_;
  assign _0534_ = ~a[6];
  assign _0545_ = _1726_ & a[4];
  assign _0556_ = _0545_ & a[5];
  assign _0567_ = _0556_ & _0534_;
  assign _0578_ = _0567_ & _0654_;
  assign _0589_ = _1792_ & _1705_;
  assign _0600_ = _0589_ & _0762_;
  assign _0611_ = _0600_ & a[6];
  assign _0622_ = _0611_ & _0654_;
  assign _0643_ = _1868_ & _1705_;
  assign _0655_ = _0643_ & _0762_;
  assign _0666_ = _0655_ & a[6];
  assign _0677_ = _0666_ & _0654_;
  assign _0688_ = _1934_ & _1705_;
  assign _0699_ = _0688_ & _0762_;
  assign _0710_ = _0699_ & a[6];
  assign _0721_ = _0710_ & _0654_;
  assign _0763_ = _2018_ & _1705_;
  assign _0774_ = _0763_ & _0762_;
  assign _0785_ = _0774_ & a[6];
  assign _0796_ = _0785_ & _0654_;
  assign _0807_ = _2073_ & _1705_;
  assign _0818_ = _0807_ & _0762_;
  assign _0828_ = _0818_ & a[6];
  assign _0839_ = _0828_ & _0654_;
  assign _0850_ = _0839_ | _0796_;
  assign _0861_ = _2137_ & _1705_;
  assign _0873_ = _0861_ & _0762_;
  assign _0884_ = _0873_ & a[6];
  assign _0895_ = _0884_ & _0654_;
  assign _0906_ = _2192_ & _1705_;
  assign _0917_ = _0906_ & _0762_;
  assign _0928_ = _0917_ & a[6];
  assign _0938_ = _0928_ & _0654_;
  assign _0949_ = _0938_ | _0895_;
  assign _0960_ = _0949_ | _0850_;
  assign _0971_ = _0054_ & _1705_;
  assign _0983_ = _0971_ & _0762_;
  assign _0994_ = _0983_ & a[6];
  assign _1005_ = _0994_ & _0654_;
  assign _1016_ = _0109_ & _1705_;
  assign _1027_ = _1016_ & _0762_;
  assign _1038_ = _1027_ & a[6];
  assign _1048_ = _1038_ & _0654_;
  assign _1069_ = _0175_ & _1705_;
  assign _1080_ = _1069_ & _0762_;
  assign _1092_ = _1080_ & a[6];
  assign _1103_ = _1092_ & _0654_;
  assign _1114_ = _0230_ & _1705_;
  assign _1125_ = _1114_ & _0762_;
  assign _1136_ = _1125_ & a[6];
  assign _1147_ = _1136_ & _0654_;
  assign _1157_ = _1147_ | _1103_;
  assign _1209_ = _1416_ & a[5];
  assign _1220_ = _1209_ & a[6];
  assign _1231_ = _1220_ & _0654_;
  assign _1242_ = _1520_ & a[5];
  assign _1252_ = _1242_ & a[6];
  assign _1263_ = _1252_ & _0654_;
  assign _1274_ = _1263_ | _1231_;
  assign _1285_ = _1590_ & a[5];
  assign _1296_ = _1285_ & a[6];
  assign _1308_ = _1296_ & _0654_;
  assign _1319_ = _1656_ & a[5];
  assign _1330_ = _1319_ & a[6];
  assign _1341_ = _1330_ & _0654_;
  assign _1351_ = _1341_ | _1308_;
  assign _1372_ = _1737_ & a[5];
  assign _1383_ = _1372_ & a[6];
  assign _1394_ = _1383_ & _0654_;
  assign _1405_ = _1803_ & a[5];
  assign _1417_ = _1405_ & a[6];
  assign _1428_ = _1417_ & _0654_;
  assign _1439_ = _1879_ & a[5];
  assign _1440_ = _1439_ & a[6];
  assign _1441_ = _1440_ & _0654_;
  assign _1442_ = _1945_ & a[5];
  assign _1443_ = _1442_ & a[6];
  assign _1444_ = _1443_ & _0654_;
  assign _1446_ = _2029_ & a[5];
  assign _1447_ = _1446_ & a[6];
  assign _1448_ = _1447_ & _0654_;
  assign _1449_ = _2084_ & a[5];
  assign _1450_ = _1449_ & a[6];
  assign _1451_ = _1450_ & _0654_;
  assign _1452_ = _2148_ & a[5];
  assign _1454_ = _1452_ & a[6];
  assign _1455_ = _1454_ & _0654_;
  assign _1456_ = _2203_ & a[5];
  assign _1457_ = _1456_ & a[6];
  assign _1458_ = _1457_ & _0654_;
  assign _1459_ = _1458_ | _1455_;
  assign _1460_ = _0065_ & a[5];
  assign _1461_ = _1460_ & a[6];
  assign _1462_ = _1461_ & _0654_;
  assign _1464_ = _0120_ & a[5];
  assign _1465_ = _1464_ & a[6];
  assign _1466_ = _1465_ & _0654_;
  assign _1467_ = _1466_ | _1462_;
  assign _1468_ = _0186_ & a[5];
  assign _1469_ = _1468_ & a[6];
  assign _1470_ = _1469_ & _0654_;
  assign _1471_ = _0241_ & a[5];
  assign _1472_ = _1471_ & a[6];
  assign _1473_ = _1472_ & _0654_;
  assign _1475_ = _1473_ | _1470_;
  assign _1476_ = _0325_ & a[5];
  assign _1477_ = _1476_ & a[6];
  assign _1478_ = _1477_ & _0654_;
  assign _1479_ = _0369_ & a[5];
  assign _1480_ = _1479_ & a[6];
  assign _1481_ = _1480_ & _0654_;
  assign _1483_ = _0424_ & a[5];
  assign _1484_ = _1483_ & a[6];
  assign _1485_ = _1484_ & _0654_;
  assign _1486_ = _0468_ & a[5];
  assign _1487_ = _1486_ & a[6];
  assign _1488_ = _1487_ & _0654_;
  assign _1489_ = _0545_ & _0762_;
  assign _1491_ = _1489_ & a[6];
  assign _1492_ = _1491_ & _0654_;
  assign _1493_ = _0589_ & a[5];
  assign _1494_ = _1493_ & a[6];
  assign _1495_ = _1494_ & _0654_;
  assign _1496_ = _1495_ | _1492_;
  assign _1497_ = _0643_ & a[5];
  assign _1498_ = _1497_ & a[6];
  assign _1499_ = _1498_ & _0654_;
  assign _1500_ = _0688_ & a[5];
  assign _1502_ = _1500_ & a[6];
  assign _1503_ = _1502_ & _0654_;
  assign _1504_ = _1503_ | _1499_;
  assign _1505_ = _0763_ & a[5];
  assign _1506_ = _1505_ & a[6];
  assign _1507_ = _1506_ & _0654_;
  assign _1508_ = _0807_ & a[5];
  assign _1509_ = _1508_ & a[6];
  assign _1511_ = _1509_ & _0654_;
  assign _1512_ = _1511_ | _1507_;
  assign _1513_ = _0861_ & a[5];
  assign _1514_ = _1513_ & a[6];
  assign _1515_ = _1514_ & _0654_;
  assign _1516_ = _0906_ & a[5];
  assign _1517_ = _1516_ & a[6];
  assign _1518_ = _1517_ & _0654_;
  assign _1519_ = _1518_ | _1515_;
  assign _1521_ = _0971_ & a[5];
  assign _1522_ = _1521_ & a[6];
  assign _1523_ = _1522_ & _0654_;
  assign _1524_ = _1016_ & a[5];
  assign _1525_ = _1524_ & a[6];
  assign _1526_ = _1525_ & _0654_;
  assign _1527_ = _1069_ & a[5];
  assign _1528_ = _1527_ & a[6];
  assign _1529_ = _1528_ & _0654_;
  assign _1531_ = _1114_ & a[5];
  assign _1532_ = _1531_ & a[6];
  assign _1533_ = _1532_ & _0654_;
  assign _1534_ = _1445_ & _0534_;
  assign _1536_ = _1534_ & _0654_;
  assign _1537_ = _1530_ & _0534_;
  assign _1538_ = _1537_ & _0654_;
  assign _1539_ = _1601_ & _0534_;
  assign _1540_ = _1539_ & _0654_;
  assign _1541_ = _1664_ & _0534_;
  assign _1542_ = _1541_ & _0654_;
  assign _1544_ = _1748_ & _0534_;
  assign _1545_ = _1544_ & _0654_;
  assign _1546_ = _1814_ & _0534_;
  assign _1547_ = _1546_ & _0654_;
  assign _1548_ = _1547_ | _1545_;
  assign _1549_ = _1890_ & _0534_;
  assign _1550_ = _1549_ & _0654_;
  assign _1551_ = _1956_ & _0534_;
  assign _1552_ = _1551_ & _0654_;
  assign _1553_ = _2040_ & _0534_;
  assign _1554_ = _1553_ & _0654_;
  assign _1555_ = _2095_ & _0534_;
  assign _1556_ = _1555_ & _0654_;
  assign _1557_ = _1556_ | _1554_;
  assign _1558_ = _2159_ & _0534_;
  assign _1559_ = _1558_ & _0654_;
  assign _1560_ = _0000_ & _0534_;
  assign _1562_ = _1560_ & _0654_;
  assign _1563_ = _0076_ & _0534_;
  assign _1564_ = _1563_ & _0654_;
  assign _1565_ = _0131_ & _0534_;
  assign _1566_ = _1565_ & _0654_;
  assign _1567_ = _1566_ | _1564_;
  assign _1568_ = _0197_ & _0534_;
  assign _1569_ = _1568_ & _0654_;
  assign _1571_ = _0252_ & _0534_;
  assign _1572_ = _1571_ & _0654_;
  assign _1573_ = _1572_ | _1569_;
  assign _1574_ = _1573_ | _1567_;
  assign _1575_ = _0336_ & _0534_;
  assign _1576_ = _1575_ & _0654_;
  assign _1577_ = _0380_ & _0534_;
  assign _1578_ = _1577_ & _0654_;
  assign _1580_ = _1578_ | _1576_;
  assign _1581_ = _0435_ & _0534_;
  assign _1582_ = _1581_ & _0654_;
  assign _1583_ = _0479_ & _0534_;
  assign _1584_ = _1583_ & _0654_;
  assign _1585_ = _1584_ | _1582_;
  assign _1586_ = _1585_ | _1580_;
  assign _1587_ = _0600_ & _0534_;
  assign _1588_ = _1587_ & _0654_;
  assign _1589_ = _0654_ & a[6];
  assign _1591_ = _1589_ & _0556_;
  assign _1592_ = _1591_ | _1588_;
  assign _1593_ = _0655_ & _0534_;
  assign _1594_ = _1593_ & _0654_;
  assign _1595_ = _0699_ & _0534_;
  assign _1596_ = _1595_ & _0654_;
  assign _1597_ = _1596_ | _1594_;
  assign _1598_ = _1597_ | _1592_;
  assign _1599_ = _1598_ | _1586_;
  assign _1600_ = _0774_ & _0534_;
  assign _1602_ = _1600_ & _0654_;
  assign _1603_ = _0818_ & _0534_;
  assign _1604_ = _1603_ & _0654_;
  assign _1605_ = _1604_ | _1602_;
  assign _1606_ = _0873_ & _0534_;
  assign _1607_ = _1606_ & _0654_;
  assign _1608_ = _0917_ & _0534_;
  assign _1609_ = _1608_ & _0654_;
  assign _1610_ = _1609_ | _1607_;
  assign _1612_ = _0983_ & _0534_;
  assign _1613_ = _1612_ & _0654_;
  assign _1614_ = _1027_ & _0534_;
  assign _1615_ = _1614_ & _0654_;
  assign _1616_ = _1080_ & _0534_;
  assign _1617_ = _1616_ & _0654_;
  assign _1618_ = _1125_ & _0534_;
  assign _1619_ = _1618_ & _0654_;
  assign _1620_ = _1619_ | _1617_;
  assign _1622_ = _1209_ & _0534_;
  assign _1623_ = _1622_ & _0654_;
  assign _1624_ = _1242_ & _0534_;
  assign _1625_ = _1624_ & _0654_;
  assign _1626_ = _1285_ & _0534_;
  assign _1628_ = _1626_ & _0654_;
  assign _1629_ = _1319_ & _0534_;
  assign _1630_ = _1629_ & _0654_;
  assign _1631_ = _1630_ | _1628_;
  assign _1632_ = _1372_ & _0534_;
  assign _1633_ = _1632_ & _0654_;
  assign _1634_ = _1405_ & _0534_;
  assign _1635_ = _1634_ & _0654_;
  assign _1637_ = _1439_ & _0534_;
  assign _1638_ = _1637_ & _0654_;
  assign _1639_ = _1442_ & _0534_;
  assign _1640_ = _1639_ & _0654_;
  assign _1641_ = _1640_ | _1638_;
  assign _1642_ = _1446_ & _0534_;
  assign _1643_ = _1642_ & _0654_;
  assign _1644_ = _1449_ & _0534_;
  assign _1646_ = _1644_ & _0654_;
  assign _1647_ = _1646_ | _1643_;
  assign _1648_ = _1452_ & _0534_;
  assign _1649_ = _1648_ & _0654_;
  assign _1650_ = _1456_ & _0534_;
  assign _1651_ = _1650_ & _0654_;
  assign _1652_ = _1651_ | _1649_;
  assign _1653_ = _1652_ | _1647_;
  assign _1654_ = _1460_ & _0534_;
  assign _1655_ = _1654_ & _0654_;
  assign _1657_ = _1464_ & _0534_;
  assign _1658_ = _1657_ & _0654_;
  assign _1659_ = _1658_ | _1655_;
  assign _1660_ = _1468_ & _0534_;
  assign _1661_ = _1660_ & _0654_;
  assign _1662_ = _1471_ & _0534_;
  assign _1663_ = _1662_ & _0654_;
  assign _1665_ = _1476_ & _0534_;
  assign _1666_ = _1665_ & _0654_;
  assign _1667_ = _1479_ & _0534_;
  assign _1668_ = _1667_ & _0654_;
  assign _1669_ = _1668_ | _1666_;
  assign _1670_ = _1483_ & _0534_;
  assign _1671_ = _1670_ & _0654_;
  assign _1672_ = _1486_ & _0534_;
  assign _1673_ = _1672_ & _0654_;
  assign _1675_ = _1673_ | _1671_;
  assign _1676_ = _1675_ | _1669_;
  assign _1677_ = _1489_ & _0534_;
  assign _1678_ = _1677_ & _0654_;
  assign _1679_ = _1493_ & _0534_;
  assign _1680_ = _1679_ & _0654_;
  assign _1681_ = _1497_ & _0534_;
  assign _1682_ = _1681_ & _0654_;
  assign _1683_ = _1500_ & _0534_;
  assign _1685_ = _1683_ & _0654_;
  assign _1686_ = _1685_ | _1682_;
  assign _1687_ = _1505_ & _0534_;
  assign _1688_ = _1687_ & _0654_;
  assign _1689_ = _1508_ & _0534_;
  assign _1690_ = _1689_ & _0654_;
  assign _1691_ = _1690_ | _1688_;
  assign _1692_ = _1513_ & _0534_;
  assign _1693_ = _1692_ & _0654_;
  assign _1694_ = _1516_ & _0534_;
  assign _1695_ = _1694_ & _0654_;
  assign _1696_ = _1521_ & _0534_;
  assign _1697_ = _1696_ & _0654_;
  assign _1698_ = _1524_ & _0534_;
  assign _1699_ = _1698_ & _0654_;
  assign _1700_ = _1527_ & _0534_;
  assign _1701_ = _1700_ & _0654_;
  assign _1702_ = _1531_ & _0534_;
  assign _1703_ = _1702_ & _0654_;
  assign _1704_ = _1703_ | _1701_;
  assign _1706_ = _1535_ & a[7];
  assign _1707_ = _1611_ & a[7];
  assign _1708_ = _1707_ | _1706_;
  assign _1709_ = _1674_ & a[7];
  assign _1710_ = _0087_ & a[7];
  assign _1711_ = _1710_ | _1709_;
  assign _1712_ = _1711_ | _1708_;
  assign _1713_ = _1825_ & a[7];
  assign _1714_ = _1901_ & a[7];
  assign _1716_ = _1714_ | _1713_;
  assign _1717_ = _1967_ & a[7];
  assign _1718_ = _1453_ & a[7];
  assign _1719_ = _1718_ | _1717_;
  assign _1720_ = _1719_ | _1716_;
  assign _1721_ = _1720_ | _1712_;
  assign _1722_ = _2105_ & a[7];
  assign _1723_ = _2170_ & a[7];
  assign _1724_ = _1723_ | _1722_;
  assign _1725_ = _0011_ & a[7];
  assign _1727_ = _1491_ & a[7];
  assign _1728_ = _1727_ | _1725_;
  assign _1729_ = _1728_ | _1724_;
  assign _1730_ = _0142_ & a[7];
  assign _1731_ = _0208_ & a[7];
  assign _1732_ = _1731_ | _1730_;
  assign _1733_ = _0263_ & a[7];
  assign _1734_ = _2051_ & a[7];
  assign _1735_ = _1734_ | _1733_;
  assign _1736_ = _1735_ | _1732_;
  assign _1738_ = _1736_ | _1729_;
  assign _1739_ = _1738_ | _1721_;
  assign _1740_ = _0391_ & a[7];
  assign _1741_ = _0446_ & a[7];
  assign _1742_ = _1741_ | _1740_;
  assign _1743_ = _0490_ & a[7];
  assign _1744_ = _0994_ & a[7];
  assign _1745_ = _1744_ | _1743_;
  assign _1746_ = _1745_ | _1742_;
  assign _1747_ = _0611_ & a[7];
  assign _1749_ = _0666_ & a[7];
  assign _1750_ = _1749_ | _1747_;
  assign _1751_ = _0710_ & a[7];
  assign _1752_ = _0347_ & a[7];
  assign _1753_ = _1752_ | _1751_;
  assign _1754_ = _1753_ | _1750_;
  assign _1755_ = _1754_ | _1746_;
  assign _1756_ = _0828_ & a[7];
  assign _1757_ = _0884_ & a[7];
  assign _1758_ = _1757_ | _1756_;
  assign _1760_ = _0928_ & a[7];
  assign _1761_ = _1759_ & a[7];
  assign _1762_ = _1761_ | _1760_;
  assign _1763_ = _1762_ | _1758_;
  assign _1764_ = _1038_ & a[7];
  assign _1765_ = _1092_ & a[7];
  assign _1766_ = _1765_ | _1764_;
  assign _1767_ = _1136_ & a[7];
  assign _1768_ = _0785_ & a[7];
  assign _1769_ = _1768_ | _1767_;
  assign _1771_ = _1769_ | _1766_;
  assign _1772_ = _1771_ | _1763_;
  assign _1773_ = _1772_ | _1755_;
  assign _1774_ = _1773_ | _1739_;
  assign _1775_ = _1252_ & a[7];
  assign _1776_ = _1296_ & a[7];
  assign _1777_ = _1776_ | _1775_;
  assign _1778_ = _1330_ & a[7];
  assign _1779_ = _1461_ & a[7];
  assign _1780_ = _1779_ | _1778_;
  assign _1782_ = _1780_ | _1777_;
  assign _1783_ = _1417_ & a[7];
  assign _1784_ = _1440_ & a[7];
  assign _1785_ = _1784_ | _1783_;
  assign _1786_ = _1443_ & a[7];
  assign _1787_ = _1220_ & a[7];
  assign _1788_ = _1787_ | _1786_;
  assign _1789_ = _1788_ | _1785_;
  assign _1790_ = _1789_ | _1782_;
  assign _1791_ = _1457_ & a[7];
  assign _1793_ = _1450_ & a[7];
  assign _1794_ = _1454_ & a[7];
  assign _1795_ = _1794_ | _1793_;
  assign _1796_ = _1795_ | _1791_;
  assign _1797_ = _1465_ & a[7];
  assign _1798_ = _1469_ & a[7];
  assign _1799_ = _1798_ | _1797_;
  assign _1800_ = _1472_ & a[7];
  assign _1801_ = _1447_ & a[7];
  assign _1802_ = _1801_ | _1800_;
  assign _1804_ = _1802_ | _1799_;
  assign _1805_ = _1804_ | _1796_;
  assign _1806_ = _1805_ | _1790_;
  assign _1807_ = _1480_ & a[7];
  assign _1808_ = _1484_ & a[7];
  assign _1809_ = _1808_ | _1807_;
  assign _1810_ = _1487_ & a[7];
  assign _1811_ = _1522_ & a[7];
  assign _1812_ = _1811_ | _1810_;
  assign _1813_ = _1812_ | _1809_;
  assign _1815_ = _1494_ & a[7];
  assign _1816_ = _1498_ & a[7];
  assign _1817_ = _1816_ | _1815_;
  assign _1818_ = _1502_ & a[7];
  assign _1819_ = _1477_ & a[7];
  assign _1820_ = _1819_ | _1818_;
  assign _1821_ = _1820_ | _1817_;
  assign _1822_ = _1821_ | _1813_;
  assign _1823_ = _1509_ & a[7];
  assign _1824_ = _1514_ & a[7];
  assign _1826_ = _1824_ | _1823_;
  assign _1827_ = _1517_ & a[7];
  assign _1828_ = _1383_ & a[7];
  assign _1829_ = _1828_ | _1827_;
  assign _1830_ = _1829_ | _1826_;
  assign _1831_ = _1525_ & a[7];
  assign _1832_ = _1528_ & a[7];
  assign _1833_ = _1832_ | _1831_;
  assign _1834_ = _1532_ & a[7];
  assign _1835_ = _1506_ & a[7];
  assign _1837_ = _1835_ | _1834_;
  assign _1838_ = _1837_ | _1833_;
  assign _1839_ = _1838_ | _1830_;
  assign _1840_ = _1839_ | _1822_;
  assign _1841_ = _1840_ | _1806_;
  assign _1842_ = _1841_ | _1774_;
  assign _1843_ = _1537_ & a[7];
  assign _1844_ = _1539_ & a[7];
  assign _1845_ = _1844_ | _1843_;
  assign _1846_ = _1541_ & a[7];
  assign _1847_ = _1563_ & a[7];
  assign _1848_ = _1847_ | _1846_;
  assign _1849_ = _1848_ | _1845_;
  assign _1850_ = _1546_ & a[7];
  assign _1851_ = _1549_ & a[7];
  assign _1852_ = _1851_ | _1850_;
  assign _1853_ = _1551_ & a[7];
  assign _1854_ = _1534_ & a[7];
  assign _1855_ = _1854_ | _1853_;
  assign _1856_ = _1855_ | _1852_;
  assign _1858_ = _1856_ | _1849_;
  assign _1859_ = _1555_ & a[7];
  assign _1860_ = _1558_ & a[7];
  assign _1861_ = _1860_ | _1859_;
  assign _1862_ = _1560_ & a[7];
  assign _1863_ = _1677_ & a[7];
  assign _1864_ = _1863_ | _1862_;
  assign _1865_ = _1864_ | _1861_;
  assign _1866_ = _1565_ & a[7];
  assign _1867_ = _1568_ & a[7];
  assign _1869_ = _1867_ | _1866_;
  assign _1870_ = _1571_ & a[7];
  assign _1871_ = _1553_ & a[7];
  assign _1872_ = _1871_ | _1870_;
  assign _1873_ = _1872_ | _1869_;
  assign _1874_ = _1873_ | _1865_;
  assign _1875_ = _1874_ | _1858_;
  assign _1876_ = _1577_ & a[7];
  assign _1877_ = _1581_ & a[7];
  assign _1878_ = _1877_ | _1876_;
  assign _1880_ = _1583_ & a[7];
  assign _1881_ = _1612_ & a[7];
  assign _1882_ = _1881_ | _1880_;
  assign _1883_ = _1882_ | _1878_;
  assign _1884_ = _1587_ & a[7];
  assign _1885_ = _1593_ & a[7];
  assign _1886_ = _1885_ | _1884_;
  assign _1887_ = _1595_ & a[7];
  assign _1888_ = _1575_ & a[7];
  assign _1889_ = _1888_ | _1887_;
  assign _1891_ = _1889_ | _1886_;
  assign _1892_ = _1891_ | _1883_;
  assign _1893_ = _1603_ & a[7];
  assign _1894_ = _1606_ & a[7];
  assign _1895_ = _1894_ | _1893_;
  assign _1896_ = _1608_ & a[7];
  assign _1897_ = _1544_ & a[7];
  assign _1898_ = _1897_ | _1896_;
  assign _1899_ = _1898_ | _1895_;
  assign _1900_ = _1614_ & a[7];
  assign _1902_ = _1616_ & a[7];
  assign _1903_ = _1902_ | _1900_;
  assign _1904_ = _1618_ & a[7];
  assign _1905_ = _1600_ & a[7];
  assign _1906_ = _1905_ | _1904_;
  assign _1907_ = _1906_ | _1903_;
  assign _1908_ = _1907_ | _1899_;
  assign _1909_ = _1908_ | _1892_;
  assign _1910_ = _1909_ | _1875_;
  assign _1911_ = _1624_ & a[7];
  assign _1913_ = _1626_ & a[7];
  assign _1914_ = _1913_ | _1911_;
  assign _1915_ = _1629_ & a[7];
  assign _1916_ = _1654_ & a[7];
  assign _1917_ = _1916_ | _1915_;
  assign _1918_ = _1917_ | _1914_;
  assign _1919_ = _1634_ & a[7];
  assign _1920_ = _1637_ & a[7];
  assign _1921_ = _1920_ | _1919_;
  assign _1922_ = _1639_ & a[7];
  assign _1924_ = _1622_ & a[7];
  assign _1925_ = _1924_ | _1922_;
  assign _1926_ = _1925_ | _1921_;
  assign _1927_ = _1926_ | _1918_;
  assign _1928_ = _1644_ & a[7];
  assign _1929_ = _1648_ & a[7];
  assign _1930_ = _1929_ | _1928_;
  assign _1931_ = _1650_ & a[7];
  assign _1932_ = _0567_ & a[7];
  assign _1933_ = _1932_ | _1931_;
  assign _1935_ = _1933_ | _1930_;
  assign _1936_ = _1657_ & a[7];
  assign _1937_ = _1660_ & a[7];
  assign _1938_ = _1937_ | _1936_;
  assign _1939_ = _1662_ & a[7];
  assign _1940_ = _1642_ & a[7];
  assign _1941_ = _1940_ | _1939_;
  assign _1942_ = _1941_ | _1938_;
  assign _1943_ = _1942_ | _1935_;
  assign _1944_ = _1943_ | _1927_;
  assign _1946_ = _1667_ & a[7];
  assign _1947_ = _1670_ & a[7];
  assign _1948_ = _1947_ | _1946_;
  assign _1949_ = _1672_ & a[7];
  assign _1950_ = _1696_ & a[7];
  assign _1951_ = _1950_ | _1949_;
  assign _1952_ = _1951_ | _1948_;
  assign _1953_ = _1679_ & a[7];
  assign _1954_ = _1681_ & a[7];
  assign _1955_ = _1954_ | _1953_;
  assign _1957_ = _1683_ & a[7];
  assign _1958_ = _1665_ & a[7];
  assign _1959_ = _1958_ | _1957_;
  assign _1960_ = _1959_ | _1955_;
  assign _1961_ = _1960_ | _1952_;
  assign _1962_ = _1689_ & a[7];
  assign _1963_ = _1692_ & a[7];
  assign _1964_ = _1963_ | _1962_;
  assign _1965_ = _1694_ & a[7];
  assign _1966_ = _1632_ & a[7];
  assign _1968_ = _1966_ | _1965_;
  assign _1969_ = _1968_ | _1964_;
  assign _1970_ = _1698_ & a[7];
  assign _1971_ = _1700_ & a[7];
  assign _1972_ = _1971_ | _1970_;
  assign _1973_ = _1702_ & a[7];
  assign _1974_ = _1687_ & a[7];
  assign _1975_ = _1974_ | _1973_;
  assign _1976_ = _1975_ | _1972_;
  assign _1977_ = _1976_ | _1969_;
  assign _1978_ = _1977_ | _1961_;
  assign _1979_ = _1978_ | _1944_;
  assign _1980_ = _1979_ | _1910_;
  assign _1981_ = _1980_ | _1842_;
  assign _1982_ = _1981_ | _0654_;
  assign _1983_ = _1971_ | _1946_;
  assign _1984_ = _1983_ | _1964_;
  assign _1985_ = _1853_ | _1851_;
  assign _1986_ = _1985_ | _1864_;
  assign _1987_ = _1986_ | _1984_;
  assign _1988_ = _1928_ | _1916_;
  assign _1989_ = _1988_ | _1914_;
  assign _1990_ = _1966_ | _1919_;
  assign _1991_ = _1990_ | _1925_;
  assign _1992_ = _1991_ | _1989_;
  assign _1993_ = _1992_ | _1987_;
  assign _1994_ = _1887_ | _1884_;
  assign _1995_ = _1994_ | _1459_;
  assign _1996_ = _1308_ | _1231_;
  assign _1997_ = _1462_ | _1448_;
  assign _1998_ = _1997_ | _1996_;
  assign _1999_ = _1998_ | _1995_;
  assign _2000_ = _1905_ | _1894_;
  assign _2001_ = _2000_ | _1898_;
  assign _2002_ = _1902_ | _1881_;
  assign _2003_ = _2002_ | _1878_;
  assign _2004_ = _2003_ | _2001_;
  assign _2005_ = _2004_ | _1999_;
  assign _2006_ = _2005_ | _1993_;
  assign _2007_ = _1835_ | _1824_;
  assign _2008_ = _1828_ | _1784_;
  assign _2009_ = _2008_ | _2007_;
  assign _2010_ = _1834_ | _1831_;
  assign _2011_ = _2010_ | _1809_;
  assign _2012_ = _2011_ | _2009_;
  assign _2013_ = _1801_ | _1791_;
  assign _2014_ = _1800_ | _1798_;
  assign _2015_ = _2014_ | _2013_;
  assign _2016_ = _1797_ | _1775_;
  assign _2017_ = _2016_ | _1788_;
  assign _2019_ = _2017_ | _2015_;
  assign _2020_ = _2019_ | _2012_;
  assign _2021_ = _1760_ | _1757_;
  assign _2022_ = _1717_ | _1707_;
  assign _2023_ = _2022_ | _2021_;
  assign _2024_ = _1765_ | _1751_;
  assign _2025_ = _1768_ | _1756_;
  assign _2026_ = _2025_ | _2024_;
  assign _2027_ = _2026_ | _2023_;
  assign _2028_ = _1725_ | _1723_;
  assign _2030_ = _1819_ | _1815_;
  assign _2031_ = _2030_ | _2028_;
  assign _2032_ = _2031_ | _1736_;
  assign _2033_ = _2032_ | _2027_;
  assign _2034_ = _2033_ | _2020_;
  assign _2035_ = _2034_ | _2006_;
  assign _2036_ = _1704_ | _1675_;
  assign _2037_ = _1680_ | _1554_;
  assign _2038_ = _2037_ | _1686_;
  assign _2039_ = _2038_ | _2036_;
  assign _2041_ = _1630_ | _1623_;
  assign _2042_ = _2041_ | _1641_;
  assign _2043_ = _1695_ | _1633_;
  assign _2044_ = _2043_ | _1691_;
  assign _2045_ = _2044_ | _2042_;
  assign _2046_ = _2045_ | _2039_;
  assign _2047_ = _1613_ | _1584_;
  assign _2048_ = _2047_ | _1620_;
  assign _2049_ = _1596_ | _1588_;
  assign _2050_ = _1582_ | _1576_;
  assign _2052_ = _2050_ | _2049_;
  assign _2053_ = _2052_ | _2048_;
  assign _2054_ = _1540_ | _1536_;
  assign _2055_ = _1566_ | _1542_;
  assign _2056_ = _2055_ | _2054_;
  assign _2057_ = _1607_ | _1602_;
  assign _2058_ = _1609_ | _1552_;
  assign _2059_ = _2058_ | _2057_;
  assign _2060_ = _2059_ | _2056_;
  assign _2061_ = _2060_ | _2053_;
  assign _2063_ = _2061_ | _2046_;
  assign _2064_ = _1499_ | _1478_;
  assign _2065_ = _1485_ | _1481_;
  assign _2066_ = _2065_ | _2064_;
  assign _2067_ = _0219_ | _0098_;
  assign _2068_ = _1492_ | _2062_;
  assign _2069_ = _2068_ | _2067_;
  assign _2070_ = _2069_ | _2066_;
  assign _2071_ = _1518_ | _1507_;
  assign _2072_ = _1441_ | _1428_;
  assign _2074_ = _2072_ | _2071_;
  assign _2075_ = _1523_ | _1488_;
  assign _2076_ = _1529_ | _1526_;
  assign _2077_ = _2076_ | _2075_;
  assign _2078_ = _2077_ | _2074_;
  assign _2079_ = _2078_ | _2070_;
  assign _2080_ = _0677_ | _0622_;
  assign _2081_ = _1103_ | _0402_;
  assign _2082_ = _2081_ | _2080_;
  assign _2083_ = _1658_ | _1646_;
  assign _2085_ = _1649_ | _0578_;
  assign _2086_ = _2085_ | _2083_;
  assign _2087_ = _2086_ | _2082_;
  assign _2088_ = _1912_ | _1836_;
  assign _2089_ = _1684_ | _1463_;
  assign _2090_ = _2089_ | _2088_;
  assign _2091_ = _2090_ | _0960_;
  assign _2092_ = _2091_ | _2087_;
  assign _2093_ = _2092_ | _2079_;
  assign _2094_ = _2093_ | _2063_;
  assign _2096_ = _2094_ | _2035_;
  assign d[0] = _2096_ & _1982_;
  assign _2097_ = _1482_ | _1474_;
  assign _2098_ = _2097_ | a[2];
  assign _2099_ = _2098_ | a[3];
  assign _2100_ = _2099_ | _1705_;
  assign _2101_ = _2100_ | a[5];
  assign _2102_ = _2101_ | _0534_;
  assign _2103_ = _2102_ | a[7];
  assign _2104_ = a[1] | a[0];
  assign _2106_ = _2104_ | _0982_;
  assign _2107_ = _2106_ | a[3];
  assign _2108_ = _2107_ | _1705_;
  assign _2109_ = _2108_ | a[5];
  assign _2110_ = _2109_ | _0534_;
  assign _2111_ = _2110_ | a[7];
  assign _2112_ = _2111_ & _2103_;
  assign _2113_ = a[1] | _1474_;
  assign _2114_ = _2113_ | _0982_;
  assign _2115_ = _2114_ | a[3];
  assign _2117_ = _2115_ | _1705_;
  assign _2118_ = _2117_ | a[5];
  assign _2119_ = _2118_ | _0534_;
  assign _2120_ = _2119_ | a[7];
  assign _2121_ = _1482_ | a[0];
  assign _2122_ = _2121_ | _0982_;
  assign _2123_ = _2122_ | a[3];
  assign _2124_ = _2123_ | _1705_;
  assign _2125_ = _2124_ | a[5];
  assign _2126_ = _2125_ | _0534_;
  assign _2127_ = _2126_ | a[7];
  assign _2128_ = _2127_ & _2120_;
  assign _2129_ = _2128_ & _2112_;
  assign _2130_ = _2097_ | _0982_;
  assign _2131_ = _2130_ | _0872_;
  assign _2132_ = _2131_ | a[4];
  assign _2133_ = _2132_ | a[5];
  assign _2134_ = _2133_ | _0534_;
  assign _2135_ = _2134_ | a[7];
  assign _2136_ = _2104_ | a[2];
  assign _2138_ = _2136_ | a[3];
  assign _2139_ = _2138_ | _1705_;
  assign _2140_ = _2139_ | a[5];
  assign _2141_ = _2140_ | _0534_;
  assign _2142_ = _2141_ | a[7];
  assign _2143_ = _2142_ & _2135_;
  assign _2144_ = _2113_ | a[2];
  assign _2145_ = _2144_ | a[3];
  assign _2146_ = _2145_ | _1705_;
  assign _2147_ = _2146_ | a[5];
  assign _2149_ = _2147_ | _0534_;
  assign _2150_ = _2149_ | a[7];
  assign _2151_ = _2121_ | a[2];
  assign _2152_ = _2151_ | a[3];
  assign _2153_ = _2152_ | _1705_;
  assign _2154_ = _2153_ | a[5];
  assign _2155_ = _2154_ | _0534_;
  assign _2156_ = _2155_ | a[7];
  assign _2157_ = _2156_ & _2150_;
  assign _2158_ = _2157_ & _2143_;
  assign _2160_ = _2158_ & _2129_;
  assign _2161_ = _2098_ | _0872_;
  assign _2162_ = _2161_ | _1705_;
  assign _2163_ = _2162_ | a[5];
  assign _2164_ = _2163_ | _0534_;
  assign _2165_ = _2164_ | a[7];
  assign _2166_ = _2106_ | _0872_;
  assign _2167_ = _2166_ | _1705_;
  assign _2168_ = _2167_ | a[5];
  assign _2169_ = _2168_ | _0534_;
  assign _2171_ = _2169_ | a[7];
  assign _2172_ = _2171_ & _2165_;
  assign _2173_ = _2114_ | _0872_;
  assign _2174_ = _2173_ | _1705_;
  assign _2175_ = _2174_ | a[5];
  assign _2176_ = _2175_ | _0534_;
  assign _2177_ = _2176_ | a[7];
  assign _2178_ = _2122_ | _0872_;
  assign _2179_ = _2178_ | _1705_;
  assign _2180_ = _2179_ | a[5];
  assign _2182_ = _2180_ | _0534_;
  assign _2183_ = _2182_ | a[7];
  assign _2184_ = _2183_ & _2177_;
  assign _2185_ = _2184_ & _2172_;
  assign _2186_ = _2130_ | a[3];
  assign _2187_ = _2186_ | _1705_;
  assign _2188_ = _2187_ | a[5];
  assign _2189_ = _2188_ | _0534_;
  assign _2190_ = _2189_ | a[7];
  assign _2191_ = _2136_ | _0872_;
  assign _2193_ = _2191_ | _1705_;
  assign _2194_ = _2193_ | a[5];
  assign _2195_ = _2194_ | _0534_;
  assign _2196_ = _2195_ | a[7];
  assign _2197_ = _2196_ & _2190_;
  assign _2198_ = _2144_ | _0872_;
  assign _2199_ = _2198_ | _1705_;
  assign _2200_ = _2199_ | a[5];
  assign _2201_ = _2200_ | _0534_;
  assign _2202_ = _2201_ | a[7];
  assign _2204_ = _2151_ | _0872_;
  assign _2205_ = _2204_ | _1705_;
  assign _2206_ = _2205_ | a[5];
  assign _2207_ = _2206_ | _0534_;
  assign _2208_ = _2207_ | a[7];
  assign _2209_ = _2208_ & _2202_;
  assign _2210_ = _2209_ & _2197_;
  assign _2211_ = _2210_ & _2185_;
  assign _2212_ = _2211_ & _2160_;
  assign _2213_ = _2099_ | a[4];
  assign _0001_ = _2213_ | a[5];
  assign _0002_ = _0001_ | _0534_;
  assign _0003_ = _0002_ | a[7];
  assign _0004_ = _2107_ | a[4];
  assign _0005_ = _0004_ | a[5];
  assign _0006_ = _0005_ | _0534_;
  assign _0007_ = _0006_ | a[7];
  assign _0008_ = _0007_ & _0003_;
  assign _0009_ = _2115_ | a[4];
  assign _0010_ = _0009_ | a[5];
  assign _0012_ = _0010_ | _0534_;
  assign _0013_ = _0012_ | a[7];
  assign _0014_ = _2123_ | a[4];
  assign _0015_ = _0014_ | a[5];
  assign _0016_ = _0015_ | _0534_;
  assign _0017_ = _0016_ | a[7];
  assign _0018_ = _0017_ & _0013_;
  assign _0019_ = _0018_ & _0008_;
  assign _0020_ = _2131_ | _1705_;
  assign _0021_ = _0020_ | _0762_;
  assign _0023_ = _0021_ | a[6];
  assign _0024_ = _0023_ | a[7];
  assign _0025_ = _2138_ | a[4];
  assign _0026_ = _0025_ | a[5];
  assign _0027_ = _0026_ | _0534_;
  assign _0028_ = _0027_ | a[7];
  assign _0029_ = _0028_ & _0024_;
  assign _0030_ = _2145_ | a[4];
  assign _0031_ = _0030_ | a[5];
  assign _0032_ = _0031_ | _0534_;
  assign _0034_ = _0032_ | a[7];
  assign _0035_ = _2152_ | a[4];
  assign _0036_ = _0035_ | a[5];
  assign _0037_ = _0036_ | _0534_;
  assign _0038_ = _0037_ | a[7];
  assign _0039_ = _0038_ & _0034_;
  assign _0040_ = _0039_ & _0029_;
  assign _0041_ = _0040_ & _0019_;
  assign _0042_ = _2161_ | a[4];
  assign _0043_ = _0042_ | a[5];
  assign _0044_ = _0043_ | _0534_;
  assign _0045_ = _0044_ | a[7];
  assign _0046_ = _2166_ | a[4];
  assign _0047_ = _0046_ | a[5];
  assign _0048_ = _0047_ | _0534_;
  assign _0049_ = _0048_ | a[7];
  assign _0050_ = _0049_ & _0045_;
  assign _0051_ = _2173_ | a[4];
  assign _0052_ = _0051_ | a[5];
  assign _0053_ = _0052_ | _0534_;
  assign _0055_ = _0053_ | a[7];
  assign _0056_ = _2178_ | a[4];
  assign _0057_ = _0056_ | a[5];
  assign _0058_ = _0057_ | _0534_;
  assign _0059_ = _0058_ | a[7];
  assign _0060_ = _0059_ & _0055_;
  assign _0061_ = _0060_ & _0050_;
  assign _0062_ = _2186_ | a[4];
  assign _0063_ = _0062_ | a[5];
  assign _0064_ = _0063_ | _0534_;
  assign _0066_ = _0064_ | a[7];
  assign _0067_ = _2191_ | a[4];
  assign _0068_ = _0067_ | a[5];
  assign _0069_ = _0068_ | _0534_;
  assign _0070_ = _0069_ | a[7];
  assign _0071_ = _0070_ & _0066_;
  assign _0072_ = _2198_ | a[4];
  assign _0073_ = _0072_ | a[5];
  assign _0074_ = _0073_ | _0534_;
  assign _0075_ = _0074_ | a[7];
  assign _0077_ = _2204_ | a[4];
  assign _0078_ = _0077_ | a[5];
  assign _0079_ = _0078_ | _0534_;
  assign _0080_ = _0079_ | a[7];
  assign _0081_ = _0080_ & _0075_;
  assign _0082_ = _0081_ & _0071_;
  assign _0083_ = _0082_ & _0061_;
  assign _0084_ = _0083_ & _0041_;
  assign _0085_ = _0084_ & _2212_;
  assign _0086_ = _2100_ | _0762_;
  assign _0088_ = _0086_ | _0534_;
  assign _0089_ = _0088_ | a[7];
  assign _0090_ = _2108_ | _0762_;
  assign _0091_ = _0090_ | _0534_;
  assign _0092_ = _0091_ | a[7];
  assign _0093_ = _0092_ & _0089_;
  assign _0094_ = _2117_ | _0762_;
  assign _0095_ = _0094_ | _0534_;
  assign _0096_ = _0095_ | a[7];
  assign _0097_ = _2124_ | _0762_;
  assign _0099_ = _0097_ | _0534_;
  assign _0100_ = _0099_ | a[7];
  assign _0101_ = _0100_ & _0096_;
  assign _0102_ = _0101_ & _0093_;
  assign _0103_ = _2132_ | _0762_;
  assign _0104_ = _0103_ | _0534_;
  assign _0105_ = _0104_ | a[7];
  assign _0106_ = _2139_ | _0762_;
  assign _0107_ = _0106_ | _0534_;
  assign _0108_ = _0107_ | a[7];
  assign _0110_ = _0108_ & _0105_;
  assign _0111_ = _2146_ | _0762_;
  assign _0112_ = _0111_ | _0534_;
  assign _0113_ = _0112_ | a[7];
  assign _0114_ = _2153_ | _0762_;
  assign _0115_ = _0114_ | _0534_;
  assign _0116_ = _0115_ | a[7];
  assign _0117_ = _0116_ & _0113_;
  assign _0118_ = _0117_ & _0110_;
  assign _0119_ = _0118_ & _0102_;
  assign _0121_ = _2162_ | _0762_;
  assign _0122_ = _0121_ | _0534_;
  assign _0123_ = _0122_ | a[7];
  assign _0124_ = _2167_ | _0762_;
  assign _0125_ = _0124_ | _0534_;
  assign _0126_ = _0125_ | a[7];
  assign _0127_ = _0126_ & _0123_;
  assign _0128_ = _2174_ | _0762_;
  assign _0129_ = _0128_ | _0534_;
  assign _0130_ = _0129_ | a[7];
  assign _0132_ = _2179_ | _0762_;
  assign _0133_ = _0132_ | _0534_;
  assign _0134_ = _0133_ | a[7];
  assign _0135_ = _0134_ & _0130_;
  assign _0136_ = _0135_ & _0127_;
  assign _0137_ = _2187_ | _0762_;
  assign _0138_ = _0137_ | _0534_;
  assign _0139_ = _0138_ | a[7];
  assign _0140_ = _2193_ | _0762_;
  assign _0141_ = _0140_ | _0534_;
  assign _0143_ = _0141_ | a[7];
  assign _0144_ = _0143_ & _0139_;
  assign _0145_ = _2199_ | _0762_;
  assign _0146_ = _0145_ | _0534_;
  assign _0147_ = _0146_ | a[7];
  assign _0148_ = _2205_ | _0762_;
  assign _0149_ = _0148_ | _0534_;
  assign _0150_ = _0149_ | a[7];
  assign _0151_ = _0150_ & _0147_;
  assign _0152_ = _0151_ & _0144_;
  assign _0154_ = _0152_ & _0136_;
  assign _0155_ = _0154_ & _0119_;
  assign _0156_ = _2213_ | _0762_;
  assign _0157_ = _0156_ | _0534_;
  assign _0158_ = _0157_ | a[7];
  assign _0159_ = _0004_ | _0762_;
  assign _0160_ = _0159_ | _0534_;
  assign _0161_ = _0160_ | a[7];
  assign _0162_ = _0161_ & _0158_;
  assign _0163_ = _0009_ | _0762_;
  assign _0165_ = _0163_ | _0534_;
  assign _0166_ = _0165_ | a[7];
  assign _0167_ = _0014_ | _0762_;
  assign _0168_ = _0167_ | _0534_;
  assign _0169_ = _0168_ | a[7];
  assign _0170_ = _0169_ & _0166_;
  assign _0171_ = _0170_ & _0162_;
  assign _0172_ = _0020_ | a[5];
  assign _0173_ = _0172_ | _0534_;
  assign _0174_ = _0173_ | a[7];
  assign _0176_ = _0025_ | _0762_;
  assign _0177_ = _0176_ | _0534_;
  assign _0178_ = _0177_ | a[7];
  assign _0179_ = _0178_ & _0174_;
  assign _0180_ = _0030_ | _0762_;
  assign _0181_ = _0180_ | _0534_;
  assign _0182_ = _0181_ | a[7];
  assign _0183_ = _0035_ | _0762_;
  assign _0184_ = _0183_ | _0534_;
  assign _0185_ = _0184_ | a[7];
  assign _0187_ = _0185_ & _0182_;
  assign _0188_ = _0187_ & _0179_;
  assign _0189_ = _0188_ & _0171_;
  assign _0190_ = _0042_ | _0762_;
  assign _0191_ = _0190_ | _0534_;
  assign _0192_ = _0191_ | a[7];
  assign _0193_ = _0046_ | _0762_;
  assign _0194_ = _0193_ | _0534_;
  assign _0195_ = _0194_ | a[7];
  assign _0196_ = _0195_ & _0192_;
  assign _0198_ = _0051_ | _0762_;
  assign _0199_ = _0198_ | _0534_;
  assign _0200_ = _0199_ | a[7];
  assign _0201_ = _0056_ | _0762_;
  assign _0202_ = _0201_ | _0534_;
  assign _0203_ = _0202_ | a[7];
  assign _0204_ = _0203_ & _0200_;
  assign _0205_ = _0204_ & _0196_;
  assign _0206_ = _0062_ | _0762_;
  assign _0207_ = _0206_ | _0534_;
  assign _0209_ = _0207_ | a[7];
  assign _0210_ = _0067_ | _0762_;
  assign _0211_ = _0210_ | _0534_;
  assign _0212_ = _0211_ | a[7];
  assign _0213_ = _0212_ & _0209_;
  assign _0214_ = _0072_ | _0762_;
  assign _0215_ = _0214_ | _0534_;
  assign _0216_ = _0215_ | a[7];
  assign _0217_ = _0077_ | _0762_;
  assign _0218_ = _0217_ | _0534_;
  assign _0220_ = _0218_ | a[7];
  assign _0221_ = _0220_ & _0216_;
  assign _0222_ = _0221_ & _0213_;
  assign _0223_ = _0222_ & _0205_;
  assign _0224_ = _0223_ & _0189_;
  assign _0225_ = _0224_ & _0155_;
  assign _0226_ = _0225_ & _0085_;
  assign _0227_ = _2101_ | a[6];
  assign _0228_ = _0227_ | a[7];
  assign _0229_ = _2109_ | a[6];
  assign _0231_ = _0229_ | a[7];
  assign _0232_ = _0231_ & _0228_;
  assign _0233_ = _2118_ | a[6];
  assign _0234_ = _0233_ | a[7];
  assign _0235_ = _2125_ | a[6];
  assign _0236_ = _0235_ | a[7];
  assign _0237_ = _0236_ & _0234_;
  assign _0238_ = _0237_ & _0232_;
  assign _0239_ = _2133_ | a[6];
  assign _0240_ = _0239_ | a[7];
  assign _0242_ = _2140_ | a[6];
  assign _0243_ = _0242_ | a[7];
  assign _0244_ = _0243_ & _0240_;
  assign _0245_ = _2147_ | a[6];
  assign _0246_ = _0245_ | a[7];
  assign _0247_ = _2154_ | a[6];
  assign _0248_ = _0247_ | a[7];
  assign _0249_ = _0248_ & _0246_;
  assign _0250_ = _0249_ & _0244_;
  assign _0251_ = _0250_ & _0238_;
  assign _0253_ = _2163_ | a[6];
  assign _0254_ = _0253_ | a[7];
  assign _0255_ = _2168_ | a[6];
  assign _0256_ = _0255_ | a[7];
  assign _0257_ = _0256_ & _0254_;
  assign _0258_ = _2175_ | a[6];
  assign _0259_ = _0258_ | a[7];
  assign _0260_ = _2180_ | a[6];
  assign _0261_ = _0260_ | a[7];
  assign _0262_ = _0261_ & _0259_;
  assign _0264_ = _0262_ & _0257_;
  assign _0265_ = _2188_ | a[6];
  assign _0266_ = _0265_ | a[7];
  assign _0267_ = _2194_ | a[6];
  assign _0268_ = _0267_ | a[7];
  assign _0269_ = _0268_ & _0266_;
  assign _0270_ = _2200_ | a[6];
  assign _0271_ = _0270_ | a[7];
  assign _0272_ = _2206_ | a[6];
  assign _0273_ = _0272_ | a[7];
  assign _0275_ = _0273_ & _0271_;
  assign _0276_ = _0275_ & _0269_;
  assign _0277_ = _0276_ & _0264_;
  assign _0278_ = _0277_ & _0251_;
  assign _0279_ = _0001_ | a[6];
  assign _0280_ = _0279_ | a[7];
  assign _0281_ = _0005_ | a[6];
  assign _0282_ = _0281_ | a[7];
  assign _0283_ = _0282_ & _0280_;
  assign _0284_ = _0010_ | a[6];
  assign _0285_ = _0284_ | a[7];
  assign _0286_ = _0015_ | a[6];
  assign _0287_ = _0286_ | a[7];
  assign _0288_ = _0287_ & _0285_;
  assign _0289_ = _0288_ & _0283_;
  assign _0290_ = _0026_ | a[6];
  assign _0291_ = _0290_ | a[7];
  assign _0292_ = ~_1591_;
  assign _0293_ = _0292_ & _0291_;
  assign _0294_ = _0031_ | a[6];
  assign _0295_ = _0294_ | a[7];
  assign _0296_ = _0036_ | a[6];
  assign _0297_ = _0296_ | a[7];
  assign _0298_ = _0297_ & _0295_;
  assign _0299_ = _0298_ & _0293_;
  assign _0300_ = _0299_ & _0289_;
  assign _0301_ = _0043_ | a[6];
  assign _0302_ = _0301_ | a[7];
  assign _0303_ = _0047_ | a[6];
  assign _0304_ = _0303_ | a[7];
  assign _0305_ = _0304_ & _0302_;
  assign _0306_ = _0052_ | a[6];
  assign _0307_ = _0306_ | a[7];
  assign _0308_ = _0057_ | a[6];
  assign _0309_ = _0308_ | a[7];
  assign _0310_ = _0309_ & _0307_;
  assign _0311_ = _0310_ & _0305_;
  assign _0312_ = _0063_ | a[6];
  assign _0313_ = _0312_ | a[7];
  assign _0314_ = _0068_ | a[6];
  assign _0315_ = _0314_ | a[7];
  assign _0316_ = _0315_ & _0313_;
  assign _0317_ = _0073_ | a[6];
  assign _0318_ = _0317_ | a[7];
  assign _0319_ = _0078_ | a[6];
  assign _0320_ = _0319_ | a[7];
  assign _0321_ = _0320_ & _0318_;
  assign _0322_ = _0321_ & _0316_;
  assign _0323_ = _0322_ & _0311_;
  assign _0324_ = _0323_ & _0300_;
  assign _0326_ = _0324_ & _0278_;
  assign _0327_ = _0086_ | a[6];
  assign _0328_ = _0327_ | a[7];
  assign _0329_ = _0090_ | a[6];
  assign _0330_ = _0329_ | a[7];
  assign _0331_ = _0330_ & _0328_;
  assign _0332_ = _0094_ | a[6];
  assign _0333_ = _0332_ | a[7];
  assign _0334_ = _0097_ | a[6];
  assign _0335_ = _0334_ | a[7];
  assign _0337_ = _0335_ & _0333_;
  assign _0338_ = _0337_ & _0331_;
  assign _0339_ = _0103_ | a[6];
  assign _0340_ = _0339_ | a[7];
  assign _0341_ = _0106_ | a[6];
  assign _0342_ = _0341_ | a[7];
  assign _0343_ = _0342_ & _0340_;
  assign _0344_ = _0111_ | a[6];
  assign _0345_ = _0344_ | a[7];
  assign _0346_ = _0114_ | a[6];
  assign _0348_ = _0346_ | a[7];
  assign _0349_ = _0348_ & _0345_;
  assign _0350_ = _0349_ & _0343_;
  assign _0351_ = _0350_ & _0338_;
  assign _0352_ = _0121_ | a[6];
  assign _0353_ = _0352_ | a[7];
  assign _0354_ = _0124_ | a[6];
  assign _0355_ = _0354_ | a[7];
  assign _0356_ = _0355_ & _0353_;
  assign _0357_ = _0128_ | a[6];
  assign _0359_ = _0357_ | a[7];
  assign _0360_ = _0132_ | a[6];
  assign _0361_ = _0360_ | a[7];
  assign _0362_ = _0361_ & _0359_;
  assign _0363_ = _0362_ & _0356_;
  assign _0364_ = _0137_ | a[6];
  assign _0365_ = _0364_ | a[7];
  assign _0366_ = _0140_ | a[6];
  assign _0367_ = _0366_ | a[7];
  assign _0368_ = _0367_ & _0365_;
  assign _0370_ = _0145_ | a[6];
  assign _0371_ = _0370_ | a[7];
  assign _0372_ = _0148_ | a[6];
  assign _0373_ = _0372_ | a[7];
  assign _0374_ = _0373_ & _0371_;
  assign _0375_ = _0374_ & _0368_;
  assign _0376_ = _0375_ & _0363_;
  assign _0377_ = _0376_ & _0351_;
  assign _0378_ = _0156_ | a[6];
  assign _0379_ = _0378_ | a[7];
  assign _0381_ = _0159_ | a[6];
  assign _0382_ = _0381_ | a[7];
  assign _0383_ = _0382_ & _0379_;
  assign _0384_ = _0163_ | a[6];
  assign _0385_ = _0384_ | a[7];
  assign _0386_ = _0167_ | a[6];
  assign _0387_ = _0386_ | a[7];
  assign _0388_ = _0387_ & _0385_;
  assign _0389_ = _0388_ & _0383_;
  assign _0390_ = _0172_ | a[6];
  assign _0392_ = _0390_ | a[7];
  assign _0393_ = _0176_ | a[6];
  assign _0394_ = _0393_ | a[7];
  assign _0395_ = _0394_ & _0392_;
  assign _0396_ = _0180_ | a[6];
  assign _0397_ = _0396_ | a[7];
  assign _0398_ = _0183_ | a[6];
  assign _0399_ = _0398_ | a[7];
  assign _0400_ = _0399_ & _0397_;
  assign _0401_ = _0400_ & _0395_;
  assign _0403_ = _0401_ & _0389_;
  assign _0404_ = _0190_ | a[6];
  assign _0405_ = _0404_ | a[7];
  assign _0406_ = _0193_ | a[6];
  assign _0407_ = _0406_ | a[7];
  assign _0408_ = _0407_ & _0405_;
  assign _0409_ = _0198_ | a[6];
  assign _0410_ = _0409_ | a[7];
  assign _0411_ = _0201_ | a[6];
  assign _0412_ = _0411_ | a[7];
  assign _0414_ = _0412_ & _0410_;
  assign _0415_ = _0414_ & _0408_;
  assign _0416_ = _0206_ | a[6];
  assign _0417_ = _0416_ | a[7];
  assign _0418_ = _0210_ | a[6];
  assign _0419_ = _0418_ | a[7];
  assign _0420_ = _0419_ & _0417_;
  assign _0421_ = _0214_ | a[6];
  assign _0422_ = _0421_ | a[7];
  assign _0423_ = _0217_ | a[6];
  assign _0425_ = _0423_ | a[7];
  assign _0426_ = _0425_ & _0422_;
  assign _0427_ = _0426_ & _0420_;
  assign _0428_ = _0427_ & _0415_;
  assign _0429_ = _0428_ & _0403_;
  assign _0430_ = _0429_ & _0377_;
  assign _0431_ = _0430_ & _0326_;
  assign _0432_ = _0431_ & _0226_;
  assign _0433_ = _2110_ | _0654_;
  assign _0434_ = _2119_ | _0654_;
  assign _0436_ = _0434_ & _0433_;
  assign _0437_ = _2126_ | _0654_;
  assign _0438_ = _2189_ | _0654_;
  assign _0439_ = _0438_ & _0437_;
  assign _0440_ = _0439_ & _0436_;
  assign _0441_ = _2141_ | _0654_;
  assign _0442_ = _2149_ | _0654_;
  assign _0443_ = _0442_ & _0441_;
  assign _0444_ = _2155_ | _0654_;
  assign _0445_ = _2102_ | _0654_;
  assign _0447_ = _0445_ & _0444_;
  assign _0448_ = _0447_ & _0443_;
  assign _0449_ = _0448_ & _0440_;
  assign _0450_ = _2169_ | _0654_;
  assign _0451_ = _2176_ | _0654_;
  assign _0452_ = _0451_ & _0450_;
  assign _0453_ = _2182_ | _0654_;
  assign _0454_ = _0173_ | _0654_;
  assign _0455_ = _0454_ & _0453_;
  assign _0456_ = _0455_ & _0452_;
  assign _0458_ = _2195_ | _0654_;
  assign _0459_ = _2201_ | _0654_;
  assign _0460_ = _0459_ & _0458_;
  assign _0461_ = _2207_ | _0654_;
  assign _0462_ = _2164_ | _0654_;
  assign _0463_ = _0462_ & _0461_;
  assign _0464_ = _0463_ & _0460_;
  assign _0465_ = _0464_ & _0456_;
  assign _0466_ = _0465_ & _0449_;
  assign _0467_ = _0006_ | _0654_;
  assign _0469_ = _0012_ | _0654_;
  assign _0470_ = _0469_ & _0467_;
  assign _0471_ = _0016_ | _0654_;
  assign _0472_ = _0064_ | _0654_;
  assign _0473_ = _0472_ & _0471_;
  assign _0474_ = _0473_ & _0470_;
  assign _0475_ = _0027_ | _0654_;
  assign _0476_ = _0032_ | _0654_;
  assign _0477_ = _0476_ & _0475_;
  assign _0478_ = _0037_ | _0654_;
  assign _0480_ = _0002_ | _0654_;
  assign _0481_ = _0480_ & _0478_;
  assign _0482_ = _0481_ & _0477_;
  assign _0483_ = _0482_ & _0474_;
  assign _0484_ = _0048_ | _0654_;
  assign _0485_ = _0053_ | _0654_;
  assign _0486_ = _0485_ & _0484_;
  assign _0487_ = _0058_ | _0654_;
  assign _0488_ = _2134_ | _0654_;
  assign _0489_ = _0488_ & _0487_;
  assign _0491_ = _0489_ & _0486_;
  assign _0492_ = _0069_ | _0654_;
  assign _0493_ = _0074_ | _0654_;
  assign _0494_ = _0493_ & _0492_;
  assign _0495_ = _0079_ | _0654_;
  assign _0496_ = _0044_ | _0654_;
  assign _0497_ = _0496_ & _0495_;
  assign _0498_ = _0497_ & _0494_;
  assign _0499_ = _0498_ & _0491_;
  assign _0500_ = _0499_ & _0483_;
  assign _0502_ = _0500_ & _0466_;
  assign _0503_ = _0091_ | _0654_;
  assign _0504_ = _0095_ | _0654_;
  assign _0505_ = _0504_ & _0503_;
  assign _0506_ = _0099_ | _0654_;
  assign _0507_ = _0138_ | _0654_;
  assign _0508_ = _0507_ & _0506_;
  assign _0509_ = _0508_ & _0505_;
  assign _0510_ = _0107_ | _0654_;
  assign _0511_ = _0112_ | _0654_;
  assign _0513_ = _0511_ & _0510_;
  assign _0514_ = _0115_ | _0654_;
  assign _0515_ = _0088_ | _0654_;
  assign _0516_ = _0515_ & _0514_;
  assign _0517_ = _0516_ & _0513_;
  assign _0518_ = _0517_ & _0509_;
  assign _0519_ = _0133_ | _0654_;
  assign _0520_ = _0125_ | _0654_;
  assign _0521_ = _0129_ | _0654_;
  assign _0522_ = _0521_ & _0520_;
  assign _0524_ = _0522_ & _0519_;
  assign _0525_ = _0141_ | _0654_;
  assign _0526_ = _0146_ | _0654_;
  assign _0527_ = _0526_ & _0525_;
  assign _0528_ = _0149_ | _0654_;
  assign _0529_ = _0122_ | _0654_;
  assign _0530_ = _0529_ & _0528_;
  assign _0531_ = _0530_ & _0527_;
  assign _0532_ = _0531_ & _0524_;
  assign _0533_ = _0532_ & _0518_;
  assign _0535_ = _0160_ | _0654_;
  assign _0536_ = _0165_ | _0654_;
  assign _0537_ = _0536_ & _0535_;
  assign _0538_ = _0168_ | _0654_;
  assign _0539_ = _0207_ | _0654_;
  assign _0540_ = _0539_ & _0538_;
  assign _0541_ = _0540_ & _0537_;
  assign _0542_ = _0177_ | _0654_;
  assign _0543_ = _0181_ | _0654_;
  assign _0544_ = _0543_ & _0542_;
  assign _0546_ = _0184_ | _0654_;
  assign _0547_ = _0157_ | _0654_;
  assign _0548_ = _0547_ & _0546_;
  assign _0549_ = _0548_ & _0544_;
  assign _0550_ = _0549_ & _0541_;
  assign _0551_ = _0194_ | _0654_;
  assign _0552_ = _0199_ | _0654_;
  assign _0553_ = _0552_ & _0551_;
  assign _0554_ = _0202_ | _0654_;
  assign _0555_ = _0104_ | _0654_;
  assign _0557_ = _0555_ & _0554_;
  assign _0558_ = _0557_ & _0553_;
  assign _0559_ = _0211_ | _0654_;
  assign _0560_ = _0215_ | _0654_;
  assign _0561_ = _0560_ & _0559_;
  assign _0562_ = _0218_ | _0654_;
  assign _0563_ = _0191_ | _0654_;
  assign _0564_ = _0563_ & _0562_;
  assign _0565_ = _0564_ & _0561_;
  assign _0566_ = _0565_ & _0558_;
  assign _0568_ = _0566_ & _0550_;
  assign _0569_ = _0568_ & _0533_;
  assign _0570_ = _0569_ & _0502_;
  assign _0571_ = _0229_ | _0654_;
  assign _0572_ = _0233_ | _0654_;
  assign _0573_ = _0572_ & _0571_;
  assign _0574_ = _0235_ | _0654_;
  assign _0575_ = _0265_ | _0654_;
  assign _0576_ = _0575_ & _0574_;
  assign _0577_ = _0576_ & _0573_;
  assign _0579_ = _0242_ | _0654_;
  assign _0580_ = _0245_ | _0654_;
  assign _0581_ = _0580_ & _0579_;
  assign _0582_ = _0247_ | _0654_;
  assign _0583_ = _0227_ | _0654_;
  assign _0584_ = _0583_ & _0582_;
  assign _0585_ = _0584_ & _0581_;
  assign _0586_ = _0585_ & _0577_;
  assign _0587_ = _0255_ | _0654_;
  assign _0588_ = _0258_ | _0654_;
  assign _0590_ = _0588_ & _0587_;
  assign _0591_ = _0260_ | _0654_;
  assign _0592_ = _0390_ | _0654_;
  assign _0593_ = _0592_ & _0591_;
  assign _0594_ = _0593_ & _0590_;
  assign _0595_ = _0267_ | _0654_;
  assign _0596_ = _0270_ | _0654_;
  assign _0597_ = _0596_ & _0595_;
  assign _0598_ = _0272_ | _0654_;
  assign _0599_ = _0253_ | _0654_;
  assign _0601_ = _0599_ & _0598_;
  assign _0602_ = _0601_ & _0597_;
  assign _0603_ = _0602_ & _0594_;
  assign _0604_ = _0603_ & _0586_;
  assign _0605_ = _0281_ | _0654_;
  assign _0606_ = _0284_ | _0654_;
  assign _0607_ = _0606_ & _0605_;
  assign _0608_ = _0286_ | _0654_;
  assign _0609_ = _0312_ | _0654_;
  assign _0610_ = _0609_ & _0608_;
  assign _0612_ = _0610_ & _0607_;
  assign _0613_ = _0290_ | _0654_;
  assign _0614_ = _0294_ | _0654_;
  assign _0615_ = _0614_ & _0613_;
  assign _0616_ = _0296_ | _0654_;
  assign _0617_ = _0279_ | _0654_;
  assign _0618_ = _0617_ & _0616_;
  assign _0619_ = _0618_ & _0615_;
  assign _0620_ = _0619_ & _0612_;
  assign _0621_ = _0303_ | _0654_;
  assign _0623_ = _0306_ | _0654_;
  assign _0624_ = _0623_ & _0621_;
  assign _0625_ = _0308_ | _0654_;
  assign _0626_ = _0239_ | _0654_;
  assign _0627_ = _0626_ & _0625_;
  assign _0628_ = _0627_ & _0624_;
  assign _0629_ = _0314_ | _0654_;
  assign _0630_ = _0317_ | _0654_;
  assign _0631_ = _0630_ & _0629_;
  assign _0632_ = _0319_ | _0654_;
  assign _0633_ = _0301_ | _0654_;
  assign _0634_ = _0633_ & _0632_;
  assign _0635_ = _0634_ & _0631_;
  assign _0636_ = _0635_ & _0628_;
  assign _0637_ = _0636_ & _0620_;
  assign _0638_ = _0637_ & _0604_;
  assign _0639_ = _0329_ | _0654_;
  assign _0640_ = _0332_ | _0654_;
  assign _0641_ = _0640_ & _0639_;
  assign _0642_ = _0334_ | _0654_;
  assign _0644_ = _0364_ | _0654_;
  assign _0645_ = _0644_ & _0642_;
  assign _0646_ = _0645_ & _0641_;
  assign _0647_ = _0341_ | _0654_;
  assign _0648_ = _0344_ | _0654_;
  assign _0649_ = _0648_ & _0647_;
  assign _0650_ = _0346_ | _0654_;
  assign _0651_ = _0327_ | _0654_;
  assign _0652_ = _0651_ & _0650_;
  assign _0653_ = _0652_ & _0649_;
  assign _0656_ = _0653_ & _0646_;
  assign _0657_ = _0354_ | _0654_;
  assign _0658_ = _0357_ | _0654_;
  assign _0659_ = _0658_ & _0657_;
  assign _0660_ = _0360_ | _0654_;
  assign _0661_ = _0023_ | _0654_;
  assign _0662_ = _0661_ & _0660_;
  assign _0663_ = _0662_ & _0659_;
  assign _0664_ = _0366_ | _0654_;
  assign _0665_ = _0370_ | _0654_;
  assign _0667_ = _0665_ & _0664_;
  assign _0668_ = _0372_ | _0654_;
  assign _0669_ = _0352_ | _0654_;
  assign _0670_ = _0669_ & _0668_;
  assign _0671_ = _0670_ & _0667_;
  assign _0672_ = _0671_ & _0663_;
  assign _0673_ = _0672_ & _0656_;
  assign _0674_ = _0381_ | _0654_;
  assign _0675_ = _0384_ | _0654_;
  assign _0676_ = _0675_ & _0674_;
  assign _0678_ = _0386_ | _0654_;
  assign _0679_ = _0416_ | _0654_;
  assign _0680_ = _0679_ & _0678_;
  assign _0681_ = _0680_ & _0676_;
  assign _0682_ = _0393_ | _0654_;
  assign _0683_ = _0396_ | _0654_;
  assign _0684_ = _0683_ & _0682_;
  assign _0685_ = _0398_ | _0654_;
  assign _0686_ = _0378_ | _0654_;
  assign _0687_ = _0686_ & _0685_;
  assign _0689_ = _0687_ & _0684_;
  assign _0690_ = _0689_ & _0681_;
  assign _0691_ = _0406_ | _0654_;
  assign _0692_ = _0409_ | _0654_;
  assign _0693_ = _0692_ & _0691_;
  assign _0694_ = _0411_ | _0654_;
  assign _0695_ = _0339_ | _0654_;
  assign _0696_ = _0695_ & _0694_;
  assign _0697_ = _0696_ & _0693_;
  assign _0698_ = _0418_ | _0654_;
  assign _0700_ = _0421_ | _0654_;
  assign _0701_ = _0700_ & _0698_;
  assign _0702_ = _0423_ | _0654_;
  assign _0703_ = _0404_ | _0654_;
  assign _0704_ = _0703_ & _0702_;
  assign _0705_ = _0704_ & _0701_;
  assign _0706_ = _0705_ & _0697_;
  assign _0707_ = _0706_ & _0690_;
  assign _0708_ = _0707_ & _0673_;
  assign _0709_ = _0708_ & _0638_;
  assign _0711_ = _0709_ & _0570_;
  assign _0712_ = _0711_ & _0432_;
  assign _0713_ = _1869_ | _1845_;
  assign _0714_ = _0713_ | _1865_;
  assign _0715_ = _1974_ | _1919_;
  assign _0716_ = _0715_ | _1972_;
  assign _0717_ = _1957_ | _1954_;
  assign _0718_ = _1958_ | _1947_;
  assign _0719_ = _0718_ | _0717_;
  assign _0720_ = _0719_ | _0716_;
  assign _0722_ = _0720_ | _0714_;
  assign _0723_ = _1475_ | _1459_;
  assign _0724_ = _1518_ | _1441_;
  assign _0725_ = _0724_ | _1274_;
  assign _0726_ = _0725_ | _0723_;
  assign _0727_ = _1904_ | _1902_;
  assign _0728_ = _1897_ | _1853_;
  assign _0729_ = _0728_ | _0727_;
  assign _0730_ = _1887_ | _1876_;
  assign _0731_ = _1881_ | _1877_;
  assign _0732_ = _0731_ | _0730_;
  assign _0733_ = _0732_ | _0729_;
  assign _0734_ = _0733_ | _0726_;
  assign _0735_ = _0734_ | _0722_;
  assign _0736_ = _1727_ | _1722_;
  assign _0737_ = _1831_ | _1810_;
  assign _0738_ = _0737_ | _0736_;
  assign _0739_ = _1709_ | _1707_;
  assign _0740_ = _1733_ | _1710_;
  assign _0741_ = _0740_ | _0739_;
  assign _0742_ = _0741_ | _0738_;
  assign _0743_ = _1778_ | _1777_;
  assign _0744_ = _1834_ | _1832_;
  assign _0745_ = _1828_ | _1823_;
  assign _0746_ = _0745_ | _0744_;
  assign _0747_ = _0746_ | _0743_;
  assign _0748_ = _0747_ | _0742_;
  assign _0749_ = _1931_ | _1929_;
  assign _0750_ = _1752_ | _1747_;
  assign _0751_ = _0750_ | _0749_;
  assign _0752_ = _1922_ | _1915_;
  assign _0753_ = _1940_ | _1937_;
  assign _0754_ = _0753_ | _0752_;
  assign _0755_ = _0754_ | _0751_;
  assign _0756_ = _1718_ | _1714_;
  assign _0757_ = _0756_ | _1762_;
  assign _0758_ = _1744_ | _1741_;
  assign _0759_ = _0758_ | _2025_;
  assign _0760_ = _0759_ | _0757_;
  assign _0761_ = _0760_ | _0755_;
  assign _0764_ = _0761_ | _0748_;
  assign _0765_ = _0764_ | _0735_;
  assign _0766_ = _1685_ | _1562_;
  assign _0767_ = _0766_ | _2037_;
  assign _0768_ = _1550_ | _1538_;
  assign _0769_ = _1572_ | _1542_;
  assign _0770_ = _0769_ | _0768_;
  assign _0771_ = _0770_ | _0767_;
  assign _0772_ = _1628_ | _1623_;
  assign _0773_ = _0772_ | _1641_;
  assign _0775_ = _0773_ | _1676_;
  assign _0776_ = _0775_ | _0771_;
  assign _0777_ = _1596_ | _1576_;
  assign _0778_ = _1582_ | _1578_;
  assign _0779_ = _0778_ | _0777_;
  assign _0780_ = _2013_ | _1592_;
  assign _0781_ = _0780_ | _0779_;
  assign _0782_ = _1610_ | _1548_;
  assign _0783_ = _1619_ | _1584_;
  assign _0784_ = _0783_ | _1605_;
  assign _0786_ = _0784_ | _0782_;
  assign _0787_ = _0786_ | _0781_;
  assign _0788_ = _0787_ | _0776_;
  assign _0789_ = _0219_ | _0153_;
  assign _0790_ = _0274_ | _2116_;
  assign _0791_ = _0790_ | _0789_;
  assign _0792_ = _0098_ | _1836_;
  assign _0793_ = _0792_ | _0949_;
  assign _0794_ = _0793_ | _0791_;
  assign _0795_ = _1488_ | _1481_;
  assign _0797_ = _1533_ | _1507_;
  assign _0798_ = _0797_ | _0795_;
  assign _0799_ = _1499_ | _1492_;
  assign _0800_ = _1503_ | _1478_;
  assign _0801_ = _0800_ | _0799_;
  assign _0802_ = _0801_ | _0798_;
  assign _0803_ = _0802_ | _0794_;
  assign _0804_ = _1649_ | _1646_;
  assign _0805_ = _1651_ | _0677_;
  assign _0806_ = _0805_ | _0804_;
  assign _0808_ = _1661_ | _1643_;
  assign _0809_ = _0808_ | _1659_;
  assign _0810_ = _0809_ | _0806_;
  assign _0811_ = _1103_ | _1048_;
  assign _0812_ = _1147_ | _0796_;
  assign _0813_ = _0812_ | _0811_;
  assign _0814_ = _0813_ | _0523_;
  assign _0815_ = _0814_ | _0810_;
  assign _0816_ = _0815_ | _0803_;
  assign _0817_ = _0816_ | _0788_;
  assign _0819_ = _0817_ | _0765_;
  assign d[1] = _0819_ | _0712_;
  assign _0820_ = _1924_ | _1911_;
  assign _0821_ = _1915_ | _1913_;
  assign _0822_ = _0821_ | _0820_;
  assign _0823_ = _1965_ | _1963_;
  assign _0824_ = _1922_ | _1919_;
  assign _0825_ = _0824_ | _0823_;
  assign _0826_ = _0825_ | _0822_;
  assign _0827_ = _1931_ | _1751_;
  assign _0829_ = _1752_ | _1740_;
  assign _0830_ = _0829_ | _0827_;
  assign _0831_ = _1939_ | _1928_;
  assign _0832_ = _0831_ | _1938_;
  assign _0833_ = _0832_ | _0830_;
  assign _0834_ = _0833_ | _0826_;
  assign _0835_ = _1893_ | _1853_;
  assign _0836_ = _1866_ | _1854_;
  assign _0837_ = _0836_ | _0835_;
  assign _0838_ = _0727_ | _2000_;
  assign _0840_ = _0838_ | _0837_;
  assign _0841_ = _1949_ | _1947_;
  assign _0842_ = _1973_ | _1950_;
  assign _0843_ = _0842_ | _0841_;
  assign _0844_ = _1871_ | _1867_;
  assign _0845_ = _0844_ | _1861_;
  assign _0846_ = _0845_ | _0843_;
  assign _0847_ = _0846_ | _0840_;
  assign _0848_ = _0847_ | _0834_;
  assign _0849_ = _1834_ | _1823_;
  assign _0851_ = _1828_ | _1824_;
  assign _0852_ = _0851_ | _0849_;
  assign _0853_ = _1810_ | _1725_;
  assign _0854_ = _1832_ | _1811_;
  assign _0855_ = _0854_ | _0853_;
  assign _0856_ = _0855_ | _0852_;
  assign _0857_ = _1802_ | _1794_;
  assign _0858_ = _1787_ | _1783_;
  assign _0859_ = _0858_ | _1777_;
  assign _0860_ = _0859_ | _0857_;
  assign _0862_ = _0860_ | _0856_;
  assign _0863_ = _1757_ | _1714_;
  assign _0864_ = _0863_ | _1769_;
  assign _0865_ = _1765_ | _1743_;
  assign _0866_ = _0865_ | _0758_;
  assign _0867_ = _0866_ | _0864_;
  assign _0868_ = _1733_ | _1731_;
  assign _0869_ = _0868_ | _0736_;
  assign _0870_ = _1719_ | _1711_;
  assign _0871_ = _0870_ | _0869_;
  assign _0874_ = _0871_ | _0867_;
  assign _0875_ = _0874_ | _0862_;
  assign _0876_ = _0875_ | _0848_;
  assign _0877_ = _1697_ | _1673_;
  assign _0878_ = _1701_ | _1699_;
  assign _0879_ = _0878_ | _0877_;
  assign _0880_ = _1682_ | _1666_;
  assign _0881_ = _1671_ | _1668_;
  assign _0882_ = _0881_ | _0880_;
  assign _0883_ = _0882_ | _0879_;
  assign _0885_ = _1658_ | _1649_;
  assign _0886_ = _0885_ | _1631_;
  assign _0887_ = _1703_ | _1633_;
  assign _0888_ = _1638_ | _1635_;
  assign _0889_ = _0888_ | _0887_;
  assign _0890_ = _0889_ | _0886_;
  assign _0891_ = _0890_ | _0883_;
  assign _0892_ = _1619_ | _1604_;
  assign _0893_ = _1607_ | _1545_;
  assign _0894_ = _0893_ | _0892_;
  assign _0896_ = _2047_ | _1597_;
  assign _0897_ = _0896_ | _0894_;
  assign _0898_ = _1680_ | _1559_;
  assign _0899_ = _0898_ | _1557_;
  assign _0900_ = _1542_ | _1536_;
  assign _0901_ = _1569_ | _1566_;
  assign _0902_ = _0901_ | _0900_;
  assign _0903_ = _0902_ | _0899_;
  assign _0904_ = _0903_ | _0897_;
  assign _0905_ = _0904_ | _0891_;
  assign _0907_ = _1470_ | _1455_;
  assign _0908_ = _0907_ | _1467_;
  assign _0909_ = _1996_ | _1519_;
  assign _0910_ = _0909_ | _0908_;
  assign _0911_ = _1900_ | _1880_;
  assign _0912_ = _0911_ | _0731_;
  assign _0913_ = _1888_ | _1876_;
  assign _0914_ = _0913_ | _1886_;
  assign _0915_ = _0914_ | _0912_;
  assign _0916_ = _0915_ | _0910_;
  assign _0918_ = _0938_ | _1770_;
  assign _0919_ = _1621_ | _1463_;
  assign _0920_ = _0919_ | _0918_;
  assign _0921_ = _0721_ | _0578_;
  assign _0922_ = _1147_ | _0457_;
  assign _0923_ = _0922_ | _0921_;
  assign _0924_ = _0923_ | _0920_;
  assign _0925_ = _1523_ | _1485_;
  assign _0926_ = _1526_ | _1507_;
  assign _0927_ = _0926_ | _0925_;
  assign _0929_ = _0274_ | _2181_;
  assign _0930_ = _0929_ | _0799_;
  assign _0931_ = _0930_ | _0927_;
  assign _0932_ = _0931_ | _0924_;
  assign _0933_ = _0932_ | _0916_;
  assign _0934_ = _0933_ | _0905_;
  assign _0935_ = _0934_ | _0876_;
  assign d[2] = _0935_ | _0712_;
  assign _0936_ = _1940_ | _1936_;
  assign _0937_ = _0936_ | _1917_;
  assign _0939_ = _1966_ | _1920_;
  assign _0940_ = _0939_ | _0820_;
  assign _0941_ = _0940_ | _0937_;
  assign _0942_ = _1752_ | _1749_;
  assign _0943_ = _1764_ | _1740_;
  assign _0944_ = _0943_ | _0942_;
  assign _0945_ = _1932_ | _1747_;
  assign _0946_ = _0945_ | _0749_;
  assign _0947_ = _0946_ | _0944_;
  assign _0948_ = _0947_ | _0941_;
  assign _0950_ = _1867_ | _1847_;
  assign _0951_ = _1870_ | _1859_;
  assign _0952_ = _0951_ | _0950_;
  assign _0953_ = _1896_ | _1853_;
  assign _0954_ = _1854_ | _1844_;
  assign _0955_ = _0954_ | _0953_;
  assign _0956_ = _0955_ | _0952_;
  assign _0957_ = _1958_ | _1946_;
  assign _0958_ = _0957_ | _0842_;
  assign _0959_ = _1862_ | _1860_;
  assign _0961_ = _1957_ | _1863_;
  assign _0962_ = _0961_ | _0959_;
  assign _0963_ = _0962_ | _0958_;
  assign _0964_ = _0963_ | _0956_;
  assign _0965_ = _0964_ | _0948_;
  assign _0966_ = _1827_ | _1783_;
  assign _0967_ = _0966_ | _0745_;
  assign _0968_ = _1835_ | _1832_;
  assign _0969_ = _0968_ | _0737_;
  assign _0970_ = _0969_ | _0967_;
  assign _0972_ = _1779_ | _1775_;
  assign _0973_ = _0972_ | _1788_;
  assign _0974_ = _0973_ | _2015_;
  assign _0975_ = _0974_ | _0970_;
  assign _0976_ = _1714_ | _1706_;
  assign _0977_ = _0976_ | _1762_;
  assign _0978_ = _1768_ | _1765_;
  assign _0979_ = _0978_ | _1758_;
  assign _0980_ = _0979_ | _0977_;
  assign _0981_ = _1818_ | _1816_;
  assign _0984_ = _0981_ | _1809_;
  assign _0985_ = _1734_ | _1710_;
  assign _0986_ = _0985_ | _1728_;
  assign _0987_ = _0986_ | _0984_;
  assign _0988_ = _0987_ | _0980_;
  assign _0989_ = _0988_ | _0975_;
  assign _0990_ = _0989_ | _0965_;
  assign _0991_ = _1655_ | _1646_;
  assign _0992_ = _0721_ | _0622_;
  assign _0993_ = _0992_ | _0991_;
  assign _0995_ = _1697_ | _1671_;
  assign _0996_ = _1693_ | _1625_;
  assign _0997_ = _0996_ | _0995_;
  assign _0998_ = _0997_ | _0993_;
  assign _0999_ = _1103_ | _0839_;
  assign _1000_ = _0938_ | _1463_;
  assign _1001_ = _1000_ | _0999_;
  assign _1002_ = _1001_ | _0523_;
  assign _1003_ = _1002_ | _0998_;
  assign _1004_ = _2058_ | _1605_;
  assign _1006_ = _1594_ | _1576_;
  assign _1007_ = _1006_ | _1585_;
  assign _1008_ = _1007_ | _1004_;
  assign _1009_ = _1566_ | _1554_;
  assign _1010_ = _1682_ | _1556_;
  assign _1011_ = _1010_ | _1009_;
  assign _1012_ = _1547_ | _1536_;
  assign _1013_ = _1540_ | _1538_;
  assign _1014_ = _1013_ | _1012_;
  assign _1015_ = _1014_ | _1011_;
  assign _1017_ = _1015_ | _1008_;
  assign _1018_ = _1017_ | _1003_;
  assign _1019_ = _1473_ | _1466_;
  assign _1020_ = _1019_ | _1351_;
  assign _1021_ = _1394_ | _1231_;
  assign _1022_ = _1021_ | _1519_;
  assign _1023_ = _1022_ | _1020_;
  assign _1024_ = _1904_ | _1876_;
  assign _1025_ = _1024_ | _2000_;
  assign _1026_ = _0654_ ? _1454_ : _1587_;
  assign _1028_ = _1888_ | _1885_;
  assign _1029_ = _1028_ | _1026_;
  assign _1030_ = _1029_ | _1025_;
  assign _1031_ = _1030_ | _1023_;
  assign _1032_ = _0790_ | _2068_;
  assign _1033_ = _0098_ | _1621_;
  assign _1034_ = _1033_ | _0789_;
  assign _1035_ = _1034_ | _1032_;
  assign _1036_ = _1485_ | _1478_;
  assign _1037_ = _1529_ | _1507_;
  assign _1039_ = _1037_ | _1036_;
  assign _1040_ = _1504_ | _0033_;
  assign _1041_ = _1040_ | _1039_;
  assign _1042_ = _1041_ | _1035_;
  assign _1043_ = _1042_ | _1031_;
  assign _1044_ = _1043_ | _1018_;
  assign _1045_ = _1044_ | _0990_;
  assign d[3] = _1045_ & _1982_;
  assign _1046_ = _1971_ | _1950_;
  assign _1047_ = _1046_ | _0717_;
  assign _1049_ = _1871_ | _1859_;
  assign _1050_ = _1863_ | _1860_;
  assign _1051_ = _1050_ | _1049_;
  assign _1052_ = _1051_ | _1047_;
  assign _1053_ = _1937_ | _1913_;
  assign _1054_ = _1939_ | _1929_;
  assign _1055_ = _1054_ | _1053_;
  assign _1056_ = _1966_ | _1922_;
  assign _1057_ = _1056_ | _1964_;
  assign _1058_ = _1057_ | _1055_;
  assign _1059_ = _1058_ | _1052_;
  assign _1060_ = _1458_ | _1451_;
  assign _1061_ = _1060_ | _0907_;
  assign _1062_ = _1061_ | _0732_;
  assign _1063_ = _1897_ | _1854_;
  assign _1064_ = _1870_ | _1846_;
  assign _1065_ = _1064_ | _1063_;
  assign _1066_ = _1896_ | _1894_;
  assign _1067_ = _1066_ | _1906_;
  assign _1068_ = _1067_ | _1065_;
  assign _1070_ = _1068_ | _1062_;
  assign _1071_ = _1070_ | _1059_;
  assign _1072_ = _1811_ | _1808_;
  assign _1073_ = _1072_ | _1833_;
  assign _1074_ = _1816_ | _1727_;
  assign _1075_ = _1074_ | _1820_;
  assign _1076_ = _1075_ | _1073_;
  assign _1077_ = _1798_ | _1775_;
  assign _1078_ = _1077_ | _0851_;
  assign _1079_ = _1078_ | _1796_;
  assign _1081_ = _1079_ | _1076_;
  assign _1082_ = _1767_ | _1757_;
  assign _1083_ = _1082_ | _0978_;
  assign _1084_ = _1743_ | _1740_;
  assign _1085_ = _1084_ | _1750_;
  assign _1086_ = _1085_ | _1083_;
  assign _1087_ = _1734_ | _1725_;
  assign _1088_ = _1087_ | _0868_;
  assign _1089_ = _1717_ | _1709_;
  assign _1090_ = _1089_ | _1716_;
  assign _1093_ = _1090_ | _1088_;
  assign _1094_ = _1093_ | _1086_;
  assign _1095_ = _1094_ | _1081_;
  assign _1096_ = _1095_ | _1071_;
  assign _1097_ = _1699_ | _1688_;
  assign _1098_ = _1097_ | _1675_;
  assign _1099_ = _1680_ | _1562_;
  assign _1100_ = _1685_ | _1668_;
  assign _1101_ = _1100_ | _1099_;
  assign _1102_ = _1101_ | _1098_;
  assign _1104_ = _1628_ | _1625_;
  assign _1105_ = _1661_ | _1655_;
  assign _1106_ = _1105_ | _1104_;
  assign _1107_ = _1693_ | _1690_;
  assign _1108_ = _1107_ | _2043_;
  assign _1109_ = _1108_ | _1106_;
  assign _1110_ = _1109_ | _1102_;
  assign _1111_ = _1615_ | _1578_;
  assign _1112_ = _1607_ | _1604_;
  assign _1113_ = _1112_ | _1111_;
  assign _1115_ = _1594_ | _1591_;
  assign _1116_ = _1115_ | _0777_;
  assign _1117_ = _1116_ | _1113_;
  assign _1118_ = _1569_ | _1564_;
  assign _1119_ = _1118_ | _1010_;
  assign _1120_ = _1545_ | _1536_;
  assign _1121_ = _1120_ | _1013_;
  assign _1122_ = _1121_ | _1119_;
  assign _1123_ = _1122_ | _1117_;
  assign _1124_ = _1123_ | _1110_;
  assign _1126_ = _1515_ | _1511_;
  assign _1127_ = _1126_ | _1037_;
  assign _1128_ = _1495_ | _0022_;
  assign _1129_ = _1488_ | _1478_;
  assign _1130_ = _1129_ | _1128_;
  assign _1131_ = _1130_ | _1127_;
  assign _1132_ = _1462_ | _1341_;
  assign _1133_ = _1132_ | _1019_;
  assign _1134_ = _1518_ | _1428_;
  assign _1135_ = _1308_ | _1263_;
  assign _1137_ = _1135_ | _1134_;
  assign _1138_ = _1137_ | _1133_;
  assign _1139_ = _1138_ | _1131_;
  assign _1140_ = _1048_ | _0501_;
  assign _1141_ = _1140_ | _1157_;
  assign _1142_ = _1651_ | _0578_;
  assign _1143_ = _1142_ | _0413_;
  assign _1144_ = _1143_ | _1141_;
  assign _1145_ = _0098_ | _1684_;
  assign _1146_ = _0274_ | _2062_;
  assign _1148_ = _1146_ | _1145_;
  assign _1149_ = _0796_ | _1836_;
  assign _1150_ = _1912_ | _1621_;
  assign _1151_ = _1150_ | _1149_;
  assign _1152_ = _1151_ | _1148_;
  assign _1153_ = _1152_ | _1144_;
  assign _1154_ = _1153_ | _1139_;
  assign _1155_ = _1154_ | _1124_;
  assign _1156_ = _1155_ | _1096_;
  assign d[4] = _1156_ | _0712_;
  assign _1158_ = _1973_ | _1949_;
  assign _1159_ = _1158_ | _0717_;
  assign _1160_ = _1867_ | _1844_;
  assign _1161_ = _1953_ | _1870_;
  assign _1162_ = _1161_ | _1160_;
  assign _1163_ = _1162_ | _1159_;
  assign _1164_ = _1988_ | _1925_;
  assign _1165_ = _0715_ | _1968_;
  assign _1166_ = _1165_ | _1164_;
  assign _1167_ = _1166_ | _1163_;
  assign _1168_ = _1458_ | _1448_;
  assign _1169_ = _1168_ | _0907_;
  assign _1170_ = _1441_ | _1341_;
  assign _1171_ = _1170_ | _1467_;
  assign _1172_ = _1171_ | _1169_;
  assign _1173_ = _1897_ | _1893_;
  assign _1174_ = _1850_ | _1843_;
  assign _1175_ = _1174_ | _1173_;
  assign _1176_ = _1902_ | _1888_;
  assign _1177_ = _1176_ | _1906_;
  assign _1178_ = _1177_ | _1175_;
  assign _1179_ = _1178_ | _1172_;
  assign _1180_ = _1179_ | _1167_;
  assign _1181_ = _1734_ | _1731_;
  assign _1182_ = _1181_ | _1817_;
  assign _1183_ = _1730_ | _1709_;
  assign _1184_ = _1183_ | _1719_;
  assign _1185_ = _1184_ | _1182_;
  assign _1186_ = _1800_ | _1779_;
  assign _1187_ = _1186_ | _1777_;
  assign _1188_ = _1835_ | _1807_;
  assign _1189_ = _1827_ | _1784_;
  assign _1190_ = _1189_ | _1188_;
  assign _1191_ = _1190_ | _1187_;
  assign _1192_ = _1191_ | _1185_;
  assign _1193_ = _0827_ | _1750_;
  assign _1194_ = _1936_ | _1929_;
  assign _1195_ = _1194_ | _1941_;
  assign _1196_ = _1195_ | _1193_;
  assign _1197_ = _1082_ | _1716_;
  assign _1199_ = _1752_ | _1741_;
  assign _1200_ = _1764_ | _1743_;
  assign _1201_ = _1200_ | _1199_;
  assign _1202_ = _1201_ | _1197_;
  assign _1203_ = _1202_ | _1196_;
  assign _1204_ = _1203_ | _1192_;
  assign _1205_ = _1204_ | _1180_;
  assign _1206_ = _1572_ | _1559_;
  assign _1207_ = _1206_ | _1099_;
  assign _1208_ = _1564_ | _1538_;
  assign _1210_ = _1208_ | _1009_;
  assign _1211_ = _1210_ | _1207_;
  assign _1212_ = _1699_ | _1673_;
  assign _1213_ = _1212_ | _1704_;
  assign _1214_ = _1213_ | _0882_;
  assign _1215_ = _1214_ | _1211_;
  assign _1216_ = _1006_ | _0778_;
  assign _1217_ = _1793_ | _1791_;
  assign _1218_ = _1217_ | _2049_;
  assign _1219_ = _1218_ | _1216_;
  assign _1221_ = _1609_ | _1604_;
  assign _1222_ = _1221_ | _1120_;
  assign _1223_ = _1615_ | _1602_;
  assign _1224_ = _1223_ | _0783_;
  assign _1225_ = _1224_ | _1222_;
  assign _1226_ = _1225_ | _1219_;
  assign _1227_ = _1226_ | _1215_;
  assign _1228_ = _0153_ | _1684_;
  assign _1229_ = _1228_ | _1146_;
  assign _1230_ = _1621_ | _1543_;
  assign _1232_ = _1230_ | _1000_;
  assign _1233_ = _1232_ | _1229_;
  assign _1234_ = _1515_ | _1394_;
  assign _1235_ = _1234_ | _1037_;
  assign _1236_ = _1129_ | _1504_;
  assign _1237_ = _1236_ | _1235_;
  assign _1238_ = _1237_ | _1233_;
  assign _1239_ = _1695_ | _1640_;
  assign _1240_ = _1239_ | _1691_;
  assign _1241_ = _1240_ | _1653_;
  assign _1243_ = _0895_ | _0796_;
  assign _1244_ = _1243_ | _0999_;
  assign _1245_ = _1005_ | _0457_;
  assign _1246_ = _1245_ | _0921_;
  assign _1247_ = _1246_ | _1244_;
  assign _1248_ = _1247_ | _1241_;
  assign _1249_ = _1248_ | _1238_;
  assign _1250_ = _1249_ | _1227_;
  assign _1251_ = _1250_ | _1205_;
  assign d[5] = _1251_ & _1982_;
  assign _1253_ = _1970_ | _1950_;
  assign _1254_ = _1253_ | _1983_;
  assign _1255_ = _1953_ | _1863_;
  assign _1256_ = _1255_ | _1861_;
  assign _1257_ = _1256_ | _1254_;
  assign _1258_ = _1924_ | _1920_;
  assign _1259_ = _1258_ | _0821_;
  assign _1260_ = _1259_ | _1165_;
  assign _1261_ = _1260_ | _1257_;
  assign _1262_ = _1024_ | _0911_;
  assign _1264_ = _1888_ | _1884_;
  assign _1265_ = _1264_ | _1459_;
  assign _1266_ = _1265_ | _1262_;
  assign _1267_ = _1854_ | _1850_;
  assign _1268_ = _1267_ | _1869_;
  assign _1269_ = _0728_ | _1895_;
  assign _1270_ = _1269_ | _1268_;
  assign _1271_ = _1270_ | _1266_;
  assign _1272_ = _1271_ | _1261_;
  assign _1273_ = _1816_ | _1807_;
  assign _1275_ = _1835_ | _1808_;
  assign _1276_ = _1275_ | _1273_;
  assign _1277_ = _1733_ | _1730_;
  assign _1278_ = _1815_ | _1723_;
  assign _1279_ = _1278_ | _1277_;
  assign _1280_ = _1279_ | _1276_;
  assign _1281_ = _1797_ | _1794_;
  assign _1282_ = _1281_ | _1780_;
  assign _1283_ = _1828_ | _1776_;
  assign _1284_ = _1283_ | _1826_;
  assign _1286_ = _1284_ | _1282_;
  assign _1287_ = _1286_ | _1280_;
  assign _1288_ = _1749_ | _1744_;
  assign _1289_ = _1288_ | _1930_;
  assign _1290_ = _1289_ | _1942_;
  assign _1291_ = _1718_ | _1713_;
  assign _1292_ = _1709_ | _1706_;
  assign _1293_ = _1292_ | _1291_;
  assign _1294_ = _1767_ | _1756_;
  assign _1295_ = _1294_ | _1766_;
  assign _1297_ = _1295_ | _1293_;
  assign _1298_ = _1297_ | _1290_;
  assign _1299_ = _1298_ | _1287_;
  assign _1300_ = _1299_ | _1272_;
  assign _1301_ = _1569_ | _1562_;
  assign _1302_ = _1682_ | _1678_;
  assign _1303_ = _1302_ | _1301_;
  assign _1304_ = _1564_ | _1542_;
  assign _1305_ = _1304_ | _1013_;
  assign _1306_ = _1305_ | _1303_;
  assign _1309_ = _1638_ | _1623_;
  assign _1310_ = _1309_ | _1107_;
  assign _1311_ = _1703_ | _1688_;
  assign _1312_ = _1311_ | _0877_;
  assign _1313_ = _1312_ | _1310_;
  assign _1314_ = _1313_ | _1306_;
  assign _1315_ = _1552_ | _1536_;
  assign _1316_ = _1315_ | _1548_;
  assign _1317_ = _1619_ | _1613_;
  assign _1318_ = _1317_ | _1112_;
  assign _1320_ = _1318_ | _1316_;
  assign _1321_ = _1320_ | _1599_;
  assign _1322_ = _1321_ | _1314_;
  assign _1323_ = _1496_ | _0033_;
  assign _1324_ = _1323_ | _2066_;
  assign _1325_ = _1444_ | _1428_;
  assign _1326_ = _1473_ | _1462_;
  assign _1327_ = _1326_ | _1325_;
  assign _1328_ = _2076_ | _1512_;
  assign _1329_ = _1328_ | _1327_;
  assign _1331_ = _1329_ | _1324_;
  assign _1332_ = _1147_ | _0895_;
  assign _1333_ = _1332_ | _1140_;
  assign _1334_ = _0578_ | _0457_;
  assign _1335_ = _1334_ | _1647_;
  assign _1336_ = _1335_ | _1333_;
  assign _1337_ = _0219_ | _2116_;
  assign _1338_ = _1337_ | _0164_;
  assign _1339_ = _0919_ | _2088_;
  assign _1340_ = _1339_ | _1338_;
  assign _1342_ = _1340_ | _1336_;
  assign _1343_ = _1342_ | _1331_;
  assign _1344_ = _1343_ | _1322_;
  assign _1345_ = _1344_ | _1300_;
  assign d[6] = _1345_ & _1982_;
  assign _1346_ = _1973_ | _1962_;
  assign _1347_ = _1346_ | _0823_;
  assign _1348_ = _1255_ | _1972_;
  assign _1349_ = _1348_ | _1347_;
  assign _1350_ = _1939_ | _1916_;
  assign _1352_ = _1940_ | _1931_;
  assign _1353_ = _1352_ | _1350_;
  assign _1354_ = _1921_ | _1914_;
  assign _1355_ = _1354_ | _1353_;
  assign _1356_ = _1355_ | _1349_;
  assign _1357_ = _1900_ | _1877_;
  assign _1358_ = _1357_ | _1264_;
  assign _1359_ = _1358_ | _0723_;
  assign _1360_ = _1902_ | _1851_;
  assign _1361_ = _1854_ | _1846_;
  assign _1362_ = _1361_ | _1360_;
  assign _1363_ = _1362_ | _0952_;
  assign _1364_ = _1363_ | _1359_;
  assign _1365_ = _1364_ | _1356_;
  assign _1366_ = _0737_ | _1837_;
  assign _1367_ = _1818_ | _1815_;
  assign _1368_ = _1367_ | _1072_;
  assign _1369_ = _1368_ | _1366_;
  assign _1370_ = _1786_ | _1775_;
  assign _1371_ = _1798_ | _1776_;
  assign _1373_ = _1371_ | _1370_;
  assign _1374_ = _0745_ | _1785_;
  assign _1375_ = _1374_ | _1373_;
  assign _1376_ = _1375_ | _1369_;
  assign _1377_ = _2021_ | _1766_;
  assign _1378_ = _1747_ | _1741_;
  assign _1379_ = _1378_ | _1745_;
  assign _1380_ = _1379_ | _1377_;
  assign _1381_ = _1074_ | _1724_;
  assign _1382_ = _1761_ | _1717_;
  assign _1384_ = _1734_ | _1709_;
  assign _1385_ = _1384_ | _1382_;
  assign _1386_ = _1385_ | _1381_;
  assign _1387_ = _1386_ | _1380_;
  assign _1388_ = _1387_ | _1376_;
  assign _1389_ = _1388_ | _1365_;
  assign _1390_ = _1685_ | _1673_;
  assign _1391_ = _1390_ | _1302_;
  assign _1392_ = _1391_ | _0899_;
  assign _1393_ = _1693_ | _1638_;
  assign _1395_ = _1393_ | _0772_;
  assign _1396_ = _1701_ | _1697_;
  assign _1397_ = _1396_ | _1311_;
  assign _1398_ = _1397_ | _1395_;
  assign _1399_ = _1398_ | _1392_;
  assign _1400_ = _1613_ | _1604_;
  assign _1401_ = _1400_ | _1610_;
  assign _1402_ = _1591_ | _1578_;
  assign _1403_ = _1402_ | _1217_;
  assign _1404_ = _1403_ | _1401_;
  assign _1406_ = _1550_ | _1547_;
  assign _1407_ = _1552_ | _1538_;
  assign _1408_ = _1407_ | _1406_;
  assign _1409_ = _1408_ | _1574_;
  assign _1410_ = _1409_ | _1404_;
  assign _1411_ = _1410_ | _1399_;
  assign _1412_ = _1529_ | _1523_;
  assign _1413_ = _1412_ | _0800_;
  assign _1414_ = _1492_ | _0274_;
  assign _1415_ = _1499_ | _1495_;
  assign _1418_ = _1415_ | _1414_;
  assign _1419_ = _1418_ | _1413_;
  assign _1420_ = _1135_ | _1467_;
  assign _1421_ = _1021_ | _0724_;
  assign _1422_ = _1421_ | _1420_;
  assign _1423_ = _1422_ | _1419_;
  assign _1424_ = _1147_ | _1005_;
  assign _1425_ = _1424_ | _0805_;
  assign _1426_ = _1663_ | _1643_;
  assign _1427_ = _1426_ | _0991_;
  assign _1429_ = _1427_ | _1425_;
  assign _1430_ = _0219_ | _1684_;
  assign _1431_ = _1430_ | _0919_;
  assign _1432_ = _1912_ | _1770_;
  assign _1433_ = _1432_ | _1243_;
  assign _1434_ = _1433_ | _1431_;
  assign _1435_ = _1434_ | _1429_;
  assign _1436_ = _1435_ | _1423_;
  assign _1437_ = _1436_ | _1411_;
  assign _1438_ = _1437_ | _1389_;
  assign d[7] = _1438_ & _1982_;
endmodule
