/*
:name: parameter_range
:description: parameter with implied range tests
:should_fail: 0
:tags: 6.20.2
*/
module top();
	parameter p = 16'h1234;
endmodule
