/*
:name: 22.11--pragma-number
:description: Test
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_number 123
