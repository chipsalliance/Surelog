(* top *)
module multiclock (input clk, en1, en2, i, output q);
reg [6:0] r;
always @(posedge clk) begin
    if (en1) begin
        r[2:0] <= {r[1:0], i};
        r[6:4] <= r[5:3];
    end
    if (en2)
        r[3] <= r[2];
end
assign q = r[6];
endmodule

`ifndef _AUTOTB
module __test ;
    wire [4095:0] assert_area = "cd multiclock; select t:SRL* -assert-count 2; select t:FD* -assert-count 1";
endmodule
`endif
