module sub ();
endmodule

