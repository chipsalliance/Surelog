/*
:name: string_atooct
:description: string.atooct()  tests
:should_fail: 0
:tags: 6.16.9
*/
module top();
	string a = "777";
	int b = a.atooct();
endmodule
