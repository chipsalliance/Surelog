module top ();
  export "DPI-C" function func_1;
  function int func_1();
    return 1;
  endfunction
endmodule
