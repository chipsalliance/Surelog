/*
:name: class_test_2
:description: Test
:tags: 6.15 8.3
*/
class static Foo; endclass