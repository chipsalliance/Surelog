/*
:name: 22.7--timescale-reset
:description: Test
:tags: 22.7
:type: preprocessing
*/
`timescale 1 ns / 1 ps
`resetall
`timescale 10 us / 100 ns
