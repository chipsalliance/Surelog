`define DDR_ANA_PROG_DLY_CTRL_BIN_RANGE                7:0
`define DDR_ANA_PROG_DLY_GEAR_RANGE                    9:8
`define DDR_ANA_PROG_DLY_EN_RANGE                      10
