module top(b);
input b;
endmodule
