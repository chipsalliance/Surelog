/*
:name: typedef_test_1
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef reg[3:0] quartet;