/*
:name: desc_test_10
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef FPGA
`ifndef DEBUGGER
interface myinterface;
endinterface
`endif
`endif
