
`begin_keywords "1364-2005"
module main;

   reg [3:0] foo, bar;
   reg [1:0] adr;

   reg	     bit, rst, clk;
   reg	     load_enable, write_enable;

endmodule // main
`end_keywords

