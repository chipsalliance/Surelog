module AND();
endmodule // AND
