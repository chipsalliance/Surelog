/*
:name: associative-arrays-wildcard
:description: Test associative arrays support
:should_fail: 0
:tags: 7.8.1 7.8
*/
module top ();

int arr [*];

endmodule
