module top;
   import "DPI-C" function
     chandle test_output();

   import "DPI-C" function
     void test_input(input chandle in);
endmodule
