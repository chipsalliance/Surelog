/*
:name: typedef_test_20
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef enum logic[3:0] {
  Global = 4'h2,
  Local = 4'h3
} myenum_fwd;