module top();
adder a1();
adder a2();

wtop wtop();

endmodule

module m();
// rtl
endmodule
