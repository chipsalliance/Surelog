/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 17448
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_dqs_drvr_w_lpbk_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240, View -
//schematic
// LAST TIME SAVED: Nov 30 15:42:35 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240 (drv_out, vddq, vss, en_dn, en_up, inb_n, 
    inb_p, ncal, pcal);

output  drv_out;

inout  vddq, vss;

input  en_dn, en_up, inb_n, inb_p;

input [5:0]  pcal;
input [4:0]  ncal;

// Buses in the design

wire  [5:0]  nbb;

wire  [6:0]  p1;

wire  [6:0]  pb;

wire  [4:0]  net022;

wire  [6:0]  p;

wire  [5:0]  calp;

wire  [4:0]  dn_code;

wire  [5:0]  net023;

wire  [4:0]  caln;

wire  [5:0]  n1;

wire  [5:0]  n;

wire  [5:0]  up_code;


wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240n I4 ( .out(drv_out), .dn_code(dn_code), 
    .dn_fix(n_fix), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_6 ( .tiehi(vddq), .tielo(vss), .in(pb[6]), 
    .vss(vss), .out(p1[6]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_5 ( .tiehi(vddq), .tielo(vss), .in(pb[5]), 
    .vss(vss), .out(p1[5]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_4 ( .tiehi(vddq), .tielo(vss), .in(pb[4]), 
    .vss(vss), .out(p1[4]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_3 ( .tiehi(vddq), .tielo(vss), .in(pb[3]), 
    .vss(vss), .out(p1[3]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_2 ( .tiehi(vddq), .tielo(vss), .in(pb[2]), 
    .vss(vss), .out(p1[2]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_1 ( .tiehi(vddq), .tielo(vss), .in(pb[1]), 
    .vss(vss), .out(p1[1]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT INV1_0 ( .tiehi(vddq), .tielo(vss), .in(pb[0]), 
    .vss(vss), .out(p1[0]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV5_1 ( .in(p1[6]), .vss(vss), .out(p[6]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV5_0 ( .in(p1[5]), .vss(vss), .out(p[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_5 ( .in(nbb[5]), .vss(vss), .out(n1[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_4 ( .in(nbb[4]), .vss(vss), .out(n1[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_3 ( .in(nbb[3]), .vss(vss), .out(n1[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_2 ( .in(nbb[2]), .vss(vss), .out(n1[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_1 ( .in(nbb[1]), .vss(vss), .out(n1[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV12_0 ( .in(nbb[0]), .vss(vss), .out(n1[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV4_3 ( .in(n1[3]), .vss(vss), .out(n[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV4_2 ( .in(n1[2]), .vss(vss), .out(n[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV4_1 ( .in(n1[1]), .vss(vss), .out(n[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV4_0 ( .in(n1[0]), .vss(vss), .out(n[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV6_4 ( .in(p1[4]), .vss(vss), .out(p[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV6_3 ( .in(p1[3]), .vss(vss), .out(p[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV6_2 ( .in(p1[2]), .vss(vss), .out(p[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV6_1 ( .in(p1[1]), .vss(vss), .out(p[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV6_0 ( .in(p1[0]), .vss(vss), .out(p[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_5 ( .in(net023[5]), .vss(vss), .out(calp[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_4 ( .in(net023[4]), .vss(vss), .out(calp[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_3 ( .in(net023[3]), .vss(vss), .out(calp[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_2 ( .in(net023[2]), .vss(vss), .out(calp[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_1 ( .in(net023[1]), .vss(vss), .out(calp[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV15_0 ( .in(net023[0]), .vss(vss), .out(calp[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV16_4 ( .in(net022[4]), .vss(vss), .out(caln[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV16_3 ( .in(net022[3]), .vss(vss), .out(caln[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV16_2 ( .in(net022[2]), .vss(vss), .out(caln[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV16_1 ( .in(net022[1]), .vss(vss), .out(caln[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV16_0 ( .in(net022[0]), .vss(vss), .out(caln[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT INV14 ( .in(en_up), .vss(vss), .out(enup_b), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_6 ( .y(pb[6]), .vss(vss), .vdd(vddq), 
    .b(enup_b), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_5 ( .y(pb[5]), .vss(vss), .vdd(vddq), 
    .b(calp[5]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_4 ( .y(pb[4]), .vss(vss), .vdd(vddq), 
    .b(calp[4]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_3 ( .y(pb[3]), .vss(vss), .vdd(vddq), 
    .b(calp[3]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_2 ( .y(pb[2]), .vss(vss), .vdd(vddq), 
    .b(calp[2]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_1 ( .y(pb[1]), .vss(vss), .vdd(vddq), 
    .b(calp[1]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt NOR1_0 ( .y(pb[0]), .vss(vss), .vdd(vddq), 
    .b(calp[0]), .a(inb_p));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_7 ( .in(n[5]), .vss(vss), .out(n_fix), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_6 ( .in(n[5]), .vss(vss), .out(n_fix), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_5 ( .in(n[4]), .vss(vss), .out(dn_code[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_4 ( .in(n[4]), .vss(vss), .out(dn_code[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_3 ( .in(n[3]), .vss(vss), .out(dn_code[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_2 ( .in(n[2]), .vss(vss), .out(dn_code[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_1 ( .in(n[1]), .vss(vss), .out(dn_code[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV13_0 ( .in(n[0]), .vss(vss), .out(dn_code[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV17_1 ( .in(n1[5]), .vss(vss), .out(n[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV17_0 ( .in(n1[4]), .vss(vss), .out(n[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_8 ( .in(p[6]), .vss(vss), .out(p_fix), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_7 ( .in(p[6]), .vss(vss), .out(p_fix), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_6 ( .in(p[5]), .vss(vss), .out(up_code[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_5 ( .in(p[5]), .vss(vss), .out(up_code[5]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_4 ( .in(p[4]), .vss(vss), .out(up_code[4]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_3 ( .in(p[3]), .vss(vss), .out(up_code[3]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_2 ( .in(p[2]), .vss(vss), .out(up_code[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_1 ( .in(p[1]), .vss(vss), .out(up_code[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT INV9_0 ( .in(p[0]), .vss(vss), .out(up_code[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240p I8 ( .vddq(vddq), .vss(vss), .out(drv_out), 
    .up_code(up_code), .up_fix(p_fix));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT NAND_4 ( .tiehi(vddq), .vdd(vddq), .y(net022[4]), 
    .vss(vss), .tielo(vss), .b(ncal[4]), .a(en_dn));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT NAND_3 ( .tiehi(vddq), .vdd(vddq), .y(net022[3]), 
    .vss(vss), .tielo(vss), .b(ncal[3]), .a(en_dn));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT NAND_2 ( .tiehi(vddq), .vdd(vddq), .y(net022[2]), 
    .vss(vss), .tielo(vss), .b(ncal[2]), .a(en_dn));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT NAND_1 ( .tiehi(vddq), .vdd(vddq), .y(net022[1]), 
    .vss(vss), .tielo(vss), .b(ncal[1]), .a(en_dn));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT NAND_0 ( .tiehi(vddq), .vdd(vddq), .y(net022[0]), 
    .vss(vss), .tielo(vss), .b(ncal[0]), .a(en_dn));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_5 ( .vdd(vddq), .y(nbb[5]), .vss(vss), 
    .b(en_dn), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_4 ( .vdd(vddq), .y(nbb[4]), .vss(vss), 
    .b(caln[4]), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_3 ( .vdd(vddq), .y(nbb[3]), .vss(vss), 
    .b(caln[3]), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_2 ( .vdd(vddq), .y(nbb[2]), .vss(vss), 
    .b(caln[2]), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_1 ( .vdd(vddq), .y(nbb[1]), .vss(vss), 
    .b(caln[1]), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt NAND0_0 ( .vdd(vddq), .y(nbb[0]), .vss(vss), 
    .b(caln[0]), .a(inb_n));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_5 ( .tiehi(vddq), .tielo(vss), .y(net023[5]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[5]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_4 ( .tiehi(vddq), .tielo(vss), .y(net023[4]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[4]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_3 ( .tiehi(vddq), .tielo(vss), .y(net023[3]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[3]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_2 ( .tiehi(vddq), .tielo(vss), .y(net023[2]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_1 ( .tiehi(vddq), .tielo(vss), .y(net023[1]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT NOR_0 ( .tiehi(vddq), .tielo(vss), .y(net023[0]), 
    .vss(vss), .vdd(vddq), .b(enup_b), .a(pcal[0]));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice,
//View - schematic
// LAST TIME SAVED: Dec  2 23:33:43 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice (out_t, vddq, vss, impd, in_t, ncal, 
    ovrd, ovrd_b, ovrd_n_b, ovrd_p_b, pcal);

output  out_t;

inout  vddq, vss;

input  impd, in_t, ovrd, ovrd_b, ovrd_n_b, ovrd_p_b;

input [4:0]  ncal;
input [5:0]  pcal;


wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240 I0 ( .pcal(pcal[5:0]), .vddq(vddq), .vss(vss), 
    .drv_out(out_t), .inb_n(data_b), .inb_p(data_b), .ncal(ncal[4:0]), 
    .en_dn(impd), .en_up(impd));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_predrv INVT0 ( .pd(ovrd_n_b), .pu(ovrd_p_b), .out(data_b), 
    .en(ovrd_b), .enb(ovrd), .vss(vss), .in(in_t), .vdd(vddq));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core, View -
//schematic
// LAST TIME SAVED: Dec  2 23:34:10 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core (out_t, vddq, vss, impd, impd_b, in_t, ncal, 
    ovrd, ovrd_b, ovrd_n_b, ovrd_p_b, pcal);

output  out_t;

inout  vddq, vss;

input  in_t;

input [4:0]  ncal;
input [2:0]  ovrd_p_b;
input [2:0]  ovrd_n_b;
input [2:0]  ovrd_b;
input [2:0]  impd_b;
input [5:0]  pcal;
input [2:0]  ovrd;
input [2:0]  impd;


wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE0 ( .out_t(out_t), .impd(impd[0]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[0]), .ovrd_b(ovrd_b[0]), 
    .ovrd_n_b(ovrd_n_b[0]), .ovrd_p_b(ovrd_p_b[0]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE1_1 ( .out_t(out_t), .impd(impd[1]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[1]), .ovrd_b(ovrd_b[1]), 
    .ovrd_n_b(ovrd_n_b[1]), .ovrd_p_b(ovrd_p_b[1]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE1_0 ( .out_t(out_t), .impd(impd[1]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[1]), .ovrd_b(ovrd_b[1]), 
    .ovrd_n_b(ovrd_n_b[1]), .ovrd_p_b(ovrd_p_b[1]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE2_3 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE2_2 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE2_1 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core_slice DRV_SLICE2_0 ( .out_t(out_t), .impd(impd[2]), 
    .in_t(in_t), .ncal(ncal[4:0]), .ovrd(ovrd[2]), .ovrd_b(ovrd_b[2]), 
    .ovrd_n_b(ovrd_n_b[2]), .ovrd_p_b(ovrd_p_b[2]), .pcal(pcal[5:0]), 
    .vss(vss), .vddq(vddq));

endmodule
// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_dqs_drvr_w_lpbk_SE2DIHS_D2_GL16_RVT, View
//- schematic
// LAST TIME SAVED: Dec  3 11:26:50 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_drvr_w_lpbk_SE2DIHS_D2_GL16_RVT (outn, outp, vdd, vss, in, tiehi, tielo);

output  outn, outp;

inout  vdd, vss;

input  in, tiehi, tielo;


wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV4_1 ( .in(p1), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV4_0 ( .in(p1), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV6 ( .in(inb), .vss(vss), .out(p1), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV8 ( .in(in), .vss(vss), .out(inb), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV7 ( .in(in), .vss(vss), .out(inb), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV5_1 ( .in(n1), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV5_0 ( .in(n1), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_PU_D1_GL16_RVT PU0 ( .vdd(vdd), .en(tiehi), .y(inb));

wphy_lp4x5_dqs_drvr_w_lpbk_PU_D1_GL16_RVT PU1 ( .vdd(vdd), .en(tiehi), .y(n1));

wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT XGATE0_4 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT XGATE0_3 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT XGATE0_2 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT XGATE0_1 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT XGATE0_0 ( .y(n1), .a(inb), .en(tiehi), .enb(tielo), 
    .vdd(vdd), .vss(vss));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel INV10 ( .tiehi(tiehi), .tielo(tielo), 
    .in(outp), .vss(vss), .out(outn), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel INV3 ( .tiehi(tiehi), .tielo(tielo), 
    .in(n1), .vss(vss), .out(p1), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel INV2 ( .tiehi(tiehi), .tielo(tielo), 
    .in(p1), .vss(vss), .out(n1), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel INV9 ( .tiehi(tiehi), .tielo(tielo), 
    .in(outn), .vss(vss), .out(outp), .vdd(vdd));

wphy_lp4x5_dqs_drvr_w_lpbk_PD_D1_GL16_RVT PD0 ( .vss(vss), .enb(tielo), .y(inb));

wphy_lp4x5_dqs_drvr_w_lpbk_PD_D1_GL16_RVT PD1 ( .vss(vss), .enb(tielo), .y(n1));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_drvr_w_lpbk,
//View - schematic
// LAST TIME SAVED: Dec 14 16:24:59 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_dqs_drvr_w_lpbk (dqs_rx_in_c, dqs_rx_in_t, 
    lpbk_out_c, lpbk_out_t, pad_c, pad_t,     
    d_bs_din_c, d_bs_din_t, d_bs_ena, d_drv_impd, d_in_c, d_lpbk_ena, 
    d_ncal, d_ovrd, d_ovrd_val_c, d_ovrd_val_t, d_pcal, d_se_mode, 
    freeze_n
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vddq  
 ,vdd_aon  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vddq;
assign vddq=1'b1;
wire vdd_aon;
assign vdd_aon=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vddq;
inout vdd_aon;
inout vss;
`endif


output  dqs_rx_in_c, dqs_rx_in_t, lpbk_out_c, lpbk_out_t;

inout  pad_c, pad_t;

input  d_bs_din_c, d_bs_din_t, d_bs_ena, d_in_c, d_lpbk_ena, 
    d_ovrd_val_c, d_ovrd_val_t, d_se_mode, freeze_n;

input [2:0]  d_drv_impd;
input [5:0]  d_pcal;
input [4:0]  d_ncal;
input [2:0]  d_ovrd;

// Buses in the design 
`ifdef SYNTHESIS 
`else

wire  [2:0]  ovrd_c;

wire  [2:0]  ovrd_n_b;

wire  [2:0]  impd;

wire  [2:0]  ovrd_c_b;

wire  [2:0]  impd_b;

wire  [2:0]  ovrd_buf;

wire  [2:0]  ovrd_b;

wire  [2:0]  ovrd_p_b;

wire  [2:0]  impd_b_frz;

wire  [2:0]  net038;

wire  [2:0]  ovrd_p_c_b;

wire  [2:0]  net061;

wire  [2:0]  ovrd_b_frz;

wire  [2:0]  ovrd_n_c_b;


wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NAND2 ( .tielo(vss), .tiehi(vddq), .y(impd_b_frz[0]), 
    .vss(vss), .vdd(vddq), .b(freeze_vq), .a(d_drv_impd[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR2 ( .tielo(vss), .tiehi(vddq), .y(ovrd_b_frz[0]), 
    .vss(vss), .vdd(vddq), .b(freeze_vq), .a(d_ovrd[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR0_2 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[2]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR0_1 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[1]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR0_0 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_b[0]), 
    .vss(vss), .vdd(vddq), .b(ovrd_val_b), .a(ovrd_b[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR1_2 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_c_b[2]), 
    .vss(vss), .vdd(vddq), .b(ovrd_c_val_b), .a(ovrd_c_b[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR1_1 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_c_b[1]), 
    .vss(vss), .vdd(vddq), .b(ovrd_c_val_b), .a(ovrd_c_b[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR1_0 ( .tielo(vss), .tiehi(vddq), .y(ovrd_n_c_b[0]), 
    .vss(vss), .vdd(vddq), .b(ovrd_c_val_b), .a(ovrd_c_b[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR5_2 ( .tielo(vss), .tiehi(vddq), .y(ovrd_c_b[2]), 
    .vss(vss), .vdd(vddq), .b(d_se_mode), .a(net038[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR5_1 ( .tielo(vss), .tiehi(vddq), .y(ovrd_c_b[1]), 
    .vss(vss), .vdd(vddq), .b(d_se_mode), .a(net038[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR5_0 ( .tielo(vss), .tiehi(vddq), .y(ovrd_c_b[0]), 
    .vss(vss), .vdd(vddq), .b(d_se_mode), .a(net038[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT NOR6 ( .tielo(vss), .tiehi(vddq), .y(net041), 
    .vss(vss), .vdd(vddq), .b(net018), .a(d_se_mode));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_lvlsht_vq2va LS0 ( .d_ena(d_lpbk_ena), .vddq(vddq), 
    .out(lpbk_out_t), .outb(net023), .vss(vss), .vdda(vdda), 
    .in_vq(dqs_rx_in_t), .freeze_n(freeze_n));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_lvlsht_vq2va LS1 ( .d_ena(d_lpbk_ena), .vddq(vddq), 
    .out(lpbk_out_c), .outb(net022), .vss(vss), .vdda(vdda), 
    .in_vq(dqs_rx_in_c), .freeze_n(freeze_n));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV21_2 ( .in(impd_b_frz[2]), .vss(vss), 
    .out(net061[2]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV21_1 ( .in(impd_b_frz[1]), .vss(vss), 
    .out(net061[1]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV21_0 ( .in(impd_b_frz[0]), .vss(vss), 
    .out(net061[0]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV20 ( .in(net054), .vss(vss), .out(net053), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV16_2 ( .in(ovrd_b_frz[2]), .vss(vss), 
    .out(net038[2]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV16_1 ( .in(ovrd_b_frz[1]), .vss(vss), 
    .out(net038[1]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV16_0 ( .in(ovrd_b_frz[0]), .vss(vss), 
    .out(net038[0]), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT INV13 ( .in(freeze_n), .vss(vss), .out(freeze_vq), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_INVT_D2_GL16_RVT_withR INVT1 ( .out(pad_c), .en(bs_ena_vq), 
    .enb(bs_enb_vq), .vss(vss), .in(net028), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_INVT_D2_GL16_RVT_withR INVT0 ( .out(pad_t), .en(bs_ena_vq), 
    .enb(bs_enb_vq), .vss(vss), .in(net029), .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_hbm PRIM_ESD_C ( .vdd(vddq), .vss(vss), .pad(pad_c));

wphy_lp4x5_dqs_drvr_w_lpbk_hbm PRIM_ESD0_T ( .vdd(vddq), .vss(vss), .pad(pad_t));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND9 ( .tielo(vss), .vdd(vddq), .y(net018), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd_val_c));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND8 ( .tielo(vss), .vdd(vddq), .y(net054), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd_val_t));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND1_2 ( .tielo(vss), .vdd(vddq), .y(impd_b_frz[2]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_drv_impd[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND1_1 ( .tielo(vss), .vdd(vddq), .y(impd_b_frz[1]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_drv_impd[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND4_2 ( .tielo(vss), .vdd(vddq), .y(ovrd_b_frz[2]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND4_1 ( .tielo(vss), .vdd(vddq), .y(ovrd_b_frz[1]), 
    .vss(vss), .tiehi(vddq), .b(freeze_n_vq), .a(d_ovrd[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND7 ( .tielo(vss), .vdd(vddq), .y(bs_enb_vq), 
    .vss(vss), .tiehi(vddq), .b(freeze_n), .a(d_bs_ena));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND3_2 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_c_b[2]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_c_val_b), .a(ovrd_c[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND3_1 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_c_b[1]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_c_val_b), .a(ovrd_c[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND3_0 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_c_b[0]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_c_val_b), .a(ovrd_c[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND0_2 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[2]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[2]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND0_1 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[1]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[1]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND0_0 ( .tielo(vss), .vdd(vddq), .y(ovrd_p_b[0]), 
    .vss(vss), .tiehi(vddq), .b(ovrd_val_b), .a(ovrd_buf[0]));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND6 ( .tielo(vss), .vdd(vddq), .y(net028), 
    .vss(vss), .tiehi(vddq), .b(freeze_n), .a(d_bs_din_c));

wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT NAND5 ( .tielo(vss), .vdd(vddq), .y(net029), 
    .vss(vss), .tiehi(vddq), .b(freeze_n), .a(d_bs_din_t));

wphy_lp4x5_dqs_drvr_w_lpbk_cdm_50ohm CDM_C ( .pad(pad_c), .vdd(vddq), .vss(vss), 
    .out(dqs_rx_in_c));

wphy_lp4x5_dqs_drvr_w_lpbk_cdm_50ohm CDM_T ( .out(dqs_rx_in_t), .vss(vss), .vdd(vddq), 
    .pad(pad_t));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core DRV_T ( .ovrd(ovrd_buf[2:0]), .ovrd_b(ovrd_b[2:0]), 
    .vddq(vddq), .vss(vss), .out_t(pad_t), .impd(impd[2:0]), 
    .impd_b(impd_b[2:0]), .in_t(in_t), .ncal(d_ncal[4:0]), 
    .ovrd_n_b(ovrd_n_b[2:0]), .ovrd_p_b(ovrd_p_b[2:0]), 
    .pcal(d_pcal[5:0]));

wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_core DRV_C ( .ovrd(ovrd_c[2:0]), .ovrd_b(ovrd_c_b[2:0]), 
    .vddq(vddq), .vss(vss), .out_t(pad_c), .impd(impd[2:0]), 
    .impd_b(impd_b[2:0]), .in_t(in_c), .ncal(d_ncal[4:0]), 
    .ovrd_n_b(ovrd_n_c_b[2:0]), .ovrd_p_b(ovrd_p_c_b[2:0]), 
    .pcal(d_pcal[5:0]));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV23_2 ( .in(net061[2]), .vss(vss), .out(impd_b[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV23_1 ( .in(net061[1]), .vss(vss), .out(impd_b[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV23_0 ( .in(net061[0]), .vss(vss), .out(impd_b[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV19 ( .in(net041), .vss(vss), .out(ovrd_c_val_b), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV17 ( .in(net053), .vss(vss), .out(ovrd_val_b), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV15_2 ( .in(net038[2]), .vss(vss), .out(ovrd_b[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV15_1 ( .in(net038[1]), .vss(vss), .out(ovrd_b[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV15_0 ( .in(net038[0]), .vss(vss), .out(ovrd_b[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV14_2 ( .in(ovrd_b[2]), .vss(vss), .out(ovrd_buf[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV14_1 ( .in(ovrd_b[1]), .vss(vss), .out(ovrd_buf[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV14_0 ( .in(ovrd_b[0]), .vss(vss), .out(ovrd_buf[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV12 ( .in(freeze_vq), .vss(vss), .out(freeze_n_vq), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV25_2 ( .in(ovrd_c_b[2]), .vss(vss), .out(ovrd_c[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV25_1 ( .in(ovrd_c_b[1]), .vss(vss), .out(ovrd_c[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV25_0 ( .in(ovrd_c_b[0]), .vss(vss), .out(ovrd_c[0]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT INV24 ( .in(bs_enb_vq), .vss(vss), .out(bs_ena_vq), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_SE2DIHS_D2_GL16_RVT SE2DIFF0 ( .tiehi(vdda), .vdd(vdda), .vss(vss), 
    .tielo(vss), .outp(in_c), .outn(in_t), .in(d_in_c));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D8_GL16_RVT INV22_2 ( .in(impd_b[2]), .vss(vss), .out(impd[2]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D8_GL16_RVT INV22_1 ( .in(impd_b[1]), .vss(vss), .out(impd[1]), 
    .vdd(vddq));

wphy_lp4x5_dqs_drvr_w_lpbk_INV_D8_GL16_RVT INV22_0 ( .in(impd_b[0]), .vss(vss), .out(impd[0]), 
    .vdd(vddq));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell -
//wphy_lp4x5_dqs_drvr_w_lpbk_tb, View - schematic
// LAST TIME SAVED: Dec 17 16:38:34 2020
// NETLIST TIME: Dec 17 16:39:03 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D8_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D8_GL16_RVT ( in,  out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_PD_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_dqs_drvr_w_lpbk_PD_D1_GL16_RVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel"
//"systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_RVT_Mmod_nomodel ( in, out, tiehi, tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
  input tiehi;
  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_XG_D1_GL16_RVT ( y, en, enb, a
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input a;
  input en;
  output y;
  input enb;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign y = (en && ~enb) ? a:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_PU_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_PU_D1_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_predrv" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_predrv ( out, vdd, vss, en, enb, in, pd, pu );

  input in;
  input pu;
  output out;
  input en;
  inout vdd;
  input pd;
  input enb;
  inout vss;

wire power_ok;
assign power_ok = ~vss & vdd;

assign #(10) out= power_ok ? (en) ? ~in:1'bz : 1'bx;
assign #(10) out= (pu) ? 1'bz:1'b1;
assign #(10) out= (pd) ? 1'b0:1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_SLVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//Verilog HDL for "wavshared_tsmc14lpp_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nanad_d2_slvt ( y, a, b, vdd, vss );

  input b;
  input a;
  inout vdd;
  output y;
  inout vss;


assign y=~(a&b);


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "NAND2_D1_GL16_LVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_SLVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//Verilog HDL for "wmx_lpddr5_lib", "wmx_lpddr5_drv_240p" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240p ( out, vddq, vss, up_code, up_fix );

  input up_fix;
  output out;
  inout vddq;
  input  [5:0] up_code;
  inout vss;

  wire power_ok;
  assign power_ok = vddq & ~vss ;
  wire in_ok;
  assign in_ok = (up_code <63) == (~up_fix);
  wire  inb_pn ;
  assign inb_pn = (power_ok&in_ok) ?  ~up_fix   : 1'bx;
  

  assign (supply1, weak0) out = 	(inb_pn == 1'b1 ) ? 1'b1: 	
						 		(inb_pn == 1'b0 ) ? 1'bz : 1'bx ;
endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D4_GL16_SLVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//Verilog HDL for "wavshared_tsmc14lpp_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_nor_d2_slvt ( y, a, b, vdd, vss );

  input b;
  input a;
  inout vdd;
  output y;
  inout vss;

assign y=~(a|b);
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "INV_D2_GL16_LVT" "systemVerilog"

module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_SLVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT" "systemVerilog"

module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D1_GL16_SLVT( in, out
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign out = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out =  ~in;

endmodule
//Verilog HDL for "wmx_lpddr5_lib", "wmx_lpddr5_drv_240n" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_drv_240n ( out, dn_code, dn_fix, vss );

  input dn_fix;
  output out;
  input  [4:0] dn_code;
  inout vss;


  wire power_ok;
  assign power_ok =  ~vss ;
  wire in_ok;
  assign in_ok = (dn_code >0) == (dn_fix);
  wire  inb_pn ;
  assign inb_pn = (power_ok&in_ok) ?  dn_fix   : 1'bx;
  

  assign (supply1, weak0) out = 	(inb_pn == 1'b1 ) ? 1'b0: 	
						 		(inb_pn == 1'b0 ) ? 1'bz : 1'bx ;


endmodule
//systemVerilog HDL for "wavshared_gf12lp_ana_lib", "cdm" "systemVerilog"

module wphy_lp4x5_dqs_drvr_w_lpbk_cdm_50ohm ( out, pad, vdd, vss );

  input reg pad;
  inout vdd;
`ifdef WPIN_EN
  output integer out;
`else
  output reg out;
`endif
  inout vss;

initial begin
  if (pad === 1'bx) begin
    out = 1'bx;
  end else if (pad === 1'bz) begin
    out = 1'bz;
  end else if (pad == 1'b1) begin
`ifdef WPIN_EN
    out = 1000;
`else
    out = 1;
`endif
  end else if (pad == 1'b0) begin
    out = 0;
  end
end

always @(*) begin
  if (pad === 1'bx) begin
    out = 1'bx;
  end else if (pad === 1'bz) begin
    out = 1'bz;
  end else if (pad == 1'b1) begin
`ifdef WPIN_EN
    out = 1000;
`else
    out = 1;
`endif
  end else if (pad == 1'b0) begin
    out = 0;
  end 
end

endmodule



module wphy_lp4x5_dqs_drvr_w_lpbk_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//Verilog HDL for "wavshared_gf12lp_ana_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_hbm" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_hbm ( pad, vdd, vss );

  inout pad;
  inout vdd;
  inout vss;
endmodule
//Verilog HDL for "Serdes", "cmos_inv2_tst" "behavioral"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_INVT_D2_GL16_RVT_withR( in, vdd, vss, out, en, enb );

  inout vss;
  input in;
  inout vdd;
  input en, enb;
  output out;
  wire out;

assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//Verilog HDL for "wphy_lp4x5_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_lvlsht_vq2va" "functional"


module wphy_lp4x5_dqs_drvr_w_lpbk_wphy_lp4x5_lvlsht_vq2va ( out, outb, vdda, vddq, vss, d_ena, freeze_n, in_vq );

  inout vdda;
  output out;
  input in_vq;
  input d_ena;
  input freeze_n;
  output outb;
  inout vddq;
  inout vss;

  wire out_int;

  wire check_en;

`ifdef WANALOG_CHECK_VALID_OUT
  assign check_en=1'b1;
`else
  assign check_en=1'b0;
`endif

	wire pwr_ok;
	assign pwr_ok = vdda & freeze_n &vddq & ~vss;
   assign out_int = pwr_ok ? (in_vq &d_ena ):1'bx;
   assign out  = (check_en===1'b1 && out_int===1'bx) ? 1'b1 : out_int;    // FIXME: ADDED per Sushma's request, may remove it later
	assign outb = ~out;

//   wire pwr_ok;
//   assign pwr_ok = vdda & freeze_n &vddq & ~vss;
//   assign out = pwr_ok ? (in_vq &d_ena ):1'bx;
//   assign outb = ~out;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_drvr_w_lpbk_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
`endif //SYNTHESIS
