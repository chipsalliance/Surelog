module shift();
function logic [1-1:0] fshr_u;
  reg signed [2-1:0] signed_result;
  reg unsigned [3-1:0] unsigned_result;
  reg [4-1:0] nosign_result;
endfunction
endmodule // shift
