module alert_handler_reg_wrap;
 for (genvar i_word = 0; i_word < 8; ++i_word) begin : g_dmem_intg_check
  end
endmodule
