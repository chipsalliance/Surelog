/*
:name: class_member_test_20
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function void subr(ducktype #(3) x);
endclass