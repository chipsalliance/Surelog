/*
:name: iface_class_test_10
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic;
pure virtual function void pure_task1;
pure virtual function string concatenator(string arg);
endclass