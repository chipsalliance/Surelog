/*
:name: preproc_test_5
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`define INCEPTION(a, b, c)
