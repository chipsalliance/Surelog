/*
:name: initial
:description: initial check
:tags: 9.2.1
*/
module initial_tb ();
	reg a = 0;
	initial
		a = 1;
endmodule
