module top
(
	input x,
	input y,
	output o
);

assign o = x + y;
endmodule
