/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s001
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 15762
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_clk_div_2ph_4g_svt_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_clk_div_2ph_4g_svt_wphy_clk_div2_4g_core_svt,
//View - schematic
// LAST TIME SAVED: Sep 17 20:50:32 2020
// NETLIST TIME: Oct 27 01:15:37 2020
`timescale 1ps / 1ps 




 

module wphy_clk_div_2ph_4g_svt_wphy_clk_div2_4g_core_svt (o_clk0, o_clk90, o_clk180, o_clk270, 
    vdda, vss, i_byp, i_clk0, i_clk180, i_rst);

output  o_clk0, o_clk90, o_clk180, o_clk270;

inout  vdda, vss;

input  i_byp, i_clk0, i_clk180, i_rst;


wphy_clk_div_2ph_4g_svt_TIELO_D2_GL16_RVT I6 ( .tielo(tielo), .vss(vss), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_NOR2_D1_GL16_RVT NOR0 ( .tielo(tielo), .tiehi(tiehi), .y(rst_or_byp_n), 
    .vss(vss), .vdd(vdda), .b(i_byp), .a(i_rst));

wphy_clk_div_2ph_4g_svt_TIEHI_D2_GL16_RVT I5 ( .tiehi(tiehi), .vss(vss), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV16 ( .in(x90), .vss(vss), .out(x270), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV19 ( .in(net021), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV18 ( .in(net029), .vss(vss), .out(o_clk270), 
    .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV17 ( .in(net028), .vss(vss), .out(o_clk90), 
    .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV14 ( .in(x180), .vss(vss), .out(x0), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV20 ( .in(net030), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV1 ( .in(bypb), .vss(vss), .out(bypa), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV0 ( .in(i_byp), .vss(vss), .out(bypb), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV15 ( .in(net020), .vss(vss), .out(x90), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV2 ( .in(net015), .vss(vss), .out(x180), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT INV9 ( .in(rst_or_byp_n), .vss(vss), .out(rst_or_byp), 
    .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT I3 ( .out(net028), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk180), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT3 ( .out(net021), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk0), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT2 ( .out(net021), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x0), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT8 ( .out(net028), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x90), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT1 ( .out(net030), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x180), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT7 ( .out(net029), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x270), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT INVT0 ( .out(net030), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk180), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT I4 ( .out(net029), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk0), .vdd(vdda));

wphy_clk_div_2ph_4g_svt_LATRES_D1_GL16_RVT LAT0 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(net020), .clkb(i_clk0), 
    .clk(i_clk180), .q(net015));

wphy_clk_div_2ph_4g_svt_LATRES_D1_GL16_RVT LAT1 ( .tiehi(tiehi), .tielo(tielo), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(x180), .clkb(i_clk180), 
    .clk(i_clk0), .q(net020));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_clk_div_2ph_4g_svt, View
//- schematic
// LAST TIME SAVED: Sep 17 20:51:35 2020
// NETLIST TIME: Oct 27 01:15:38 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_clk_div_2ph_4g_svt (o_clk0, o_clk180,   i_byp, 
    i_clk0, i_clk180, i_rst
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  o_clk0, o_clk180;



input  i_byp, i_clk0, i_clk180, i_rst;

`ifdef SYNTHESIS
`else 

wphy_clk_div_2ph_4g_svt_wphy_clk_div2_4g_core_svt IDIV2 ( .o_clk90(o_clk90), 
    .o_clk270(o_clk270), .o_clk0(o_clk0), .o_clk180(o_clk180), 
    .i_byp(i_byp), .i_clk0(i_clk0), .i_clk180(i_clk180), .i_rst(i_rst), 
    .vdda(vdda), .vss(vss));

`ifdef WPHY_ANA_TIMING

specify

 if(i_byp===1'b0) 
  (i_clk0    => o_clk0)      = 136;
 if(i_byp===1'b0) 
  (i_clk180   => o_clk180)   = 136;

 if(i_byp===1'b1) 
  (i_clk0    => o_clk0)      = 62;
 if(i_byp===1'b1) 
  (i_clk180   => o_clk180)   = 62;
  //$setup(ena,posedge i_clk,45);
  //$hold(posedge i_clk,ena,30);

endspecify

`endif

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell -
//wphy_clk_div_2ph_4g_svt_tb, View - schematic
// LAST TIME SAVED: Oct 26 22:03:43 2020
// NETLIST TIME: Oct 27 01:15:38 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "LATRES_D1_GL16_LVT" "systemVerilog"


`timescale 1ps/1ps
module wphy_clk_div_2ph_4g_svt_LATRES_D1_GL16_RVT( q, clk, clkb, d, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo 
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  input clk;
  output q;
  input d;
  input clkb;
  input rstb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ? 
                           (~rstb) ? 
                                 1'b0 
                                 : (clkb) ? 
                                          (d===1'bx) ? $random : d&rstb
                                          : q 
                           : 1'bx;

endmodule

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT" "systemVerilog"


module wphy_clk_div_2ph_4g_svt_INVT_D2_GL16_RVT( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT" "systemVerilog"


module wphy_clk_div_2ph_4g_svt_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_clk_div_2ph_4g_svt_TIEHI_D2_GL16_RVT" "systemVerilog"


module wphy_clk_div_2ph_4g_svt_TIEHI_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);


  output tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tiehi = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tiehi =  1'b1 ;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clk_div_2ph_4g_svt_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_clk_div_2ph_4g_svt_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_clk_div_2ph_4g_svt_TIELO_D2_GL16_RVT" "systemVerilog"


module wphy_clk_div_2ph_4g_svt_TIELO_D2_GL16_RVT ( tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  output tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tielo = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tielo =  1'b0 ;


endmodule
`endif //SYNTHESIS
