/*
:name: class_member_test_16
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subroutine;
endclass
