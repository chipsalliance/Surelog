/*
:name: cover0_test
:description: cover #0 test
:tags: 16.4
*/
module top();

logic a = 1;

cover #0 (a != 0);

endmodule
