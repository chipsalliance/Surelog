module a(b);
input b;
reg c;parameter
signed b=b;
endmodule
