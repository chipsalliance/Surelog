/*
:name: parameter
:description: parameter tests
:tags: 6.20.2
*/
module top();
	parameter p = 123;
endmodule
