/*
:name: 22.11--pragma-invalid
:description: Test
:should_fail: 1
:tags: 22.11
:type: preprocessing
*/
`pragma
