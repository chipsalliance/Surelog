/*
:name: celldefine
:description: Celldefine check
:should_fail: 0
:tags: 5.6.4
*/

`celldefine
module cd();
endmodule
`endcelldefine

module ncd();
endmodule
