// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.11--pragma-basic
:description: Test
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_name "pragma_value"
