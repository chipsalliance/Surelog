/*
:name: class_member_test_5
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
pure virtual task pure_task1;
pure virtual task pure_task2(arg_type arg);
endclass