/*
:name: dummy_include
:description: Utility for testing `include directive
:type: preprocessing
:tags: 22.4
*/
