/*
:name: typedef_test_14
:description: Test
:tags: 6.18
*/
package some_package;
   typedef bit some_type;
endpackage

typedef some_package::some_type myalias;
