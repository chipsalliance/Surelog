module top(output int a);
   import "DPI-C" context task get_2(output int x);
endmodule // top
