/*
:name: dyn-arr-basic
:description: Test dynamic arrays support
:tags: 7.5
*/
module top ();

bit [7:0] arr[];

endmodule
