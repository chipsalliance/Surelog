/*
:name: class_member_test_36
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
virtual function virtual cmd_array_if subroutine();
endfunction
endclass