/******************************************************************************
 * (C) Copyright 2014 AMIQ Consulting
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * NAME:        amiq_eth_ve_top.sv
 * PROJECT:     amiq_eth
 * Description: This file declares the top module from which the UVM flow is run
 *******************************************************************************/

`ifndef __AMIQ_ETH_VE_TOP
	`define __AMIQ_ETH_VE_TOP
	
`timescale 10ns/10ns

`include "amiq_eth_ve_pkg.sv"

import uvm_pkg::*;
import amiq_eth_ve_pkg::*;

//top module for starting the UVM flow
module amiq_eth_ve_top;
	initial begin
		run_test();	
	end
endmodule

`endif
	