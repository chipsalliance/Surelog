module top();

	enum logic [2:0]  {
	  Global = 4'h2
	} myenum;

endmodule
