package pkg;
   typedef struct packed {
      logic 	  x;
   } a;
   typedef a[5:0] b;
endpackage // pkg
   
