/*
:name: typedef
:description: user types tests
:should_fail: 0
:tags: 6.18
*/
module top();
	typedef logic logic_t;

	logic_t a;
endmodule
