/*
:name: iface_class_test_4
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic extends base1, base2, base3;
endclass