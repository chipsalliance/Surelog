/*
:name: class_member_test_42
:description: Test
:should_fail: 0
:tags: 8.3
*/
class constructible;
function new (string name, virtual time_if vif);
  this.name = name;
endfunction
endclass