/*
:name: type_op
:description: type operator tests
:tags: 6.23
*/
module top();
	real a = 4.76;
	real b = 0.74;
	var type(a+b) c;
endmodule
