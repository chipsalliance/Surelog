/*
:name: 22.3--resetall_multiple
:description: Test
:tags: 22.3
:type: preprocessing parsing
*/
`resetall
`resetall
`resetall

module top ();
endmodule

