// Fist very simple test of the Surelog regression

module top(input logic a);

  bottom b (a);

endmodule
