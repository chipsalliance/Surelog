/*
:name: typedef
:description: user types tests
:should_fail: 0
:tags: 6.18
*/
module top();
	typedef wire wire_t;

	wire_t a;
endmodule
