// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: parameter_range
:description: parameter with implied range tests
:tags: 6.20.2
*/
module top();
	parameter p = 16'h1234;
endmodule
