module m1(input clk, output out);
  initial begin
    $display("%d", clk);
  end
endmodule
