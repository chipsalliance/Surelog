module DUT (input wire i, output reg o);
  assign o = i;
endmodule
