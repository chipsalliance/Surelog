`define DDR_ANA_SA_2PH_CAL_CODE_0_RANGE              3:0
`define DDR_ANA_SA_2PH_CAL_CODE_180_RANGE           11:8
`define DDR_ANA_SA_2PH_CAL_DIR_0_RANGE                 16
`define DDR_ANA_SA_2PH_CAL_DIR_180_RANGE               18
