module a(b);
input b;
reg c;
task a(b);

endmodule
