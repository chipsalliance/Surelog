/*
:name: celldefine
:description: Celldefine check
:tags: 5.6.4
*/

`celldefine
module cd();
endmodule
`endcelldefine

module ncd();
endmodule
