// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: typedef
:description: user types tests
:tags: 6.18
*/
module top();
	typedef logic logic_t;

	logic_t a;
endmodule
