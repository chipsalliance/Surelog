/*
:name: exit_task
:description: $exit test
:tags: 20.2
*/
module top();

initial
	$exit;

endmodule
