/*
:name: enum_typedef
:description: typedef enum tests
:tags: 6.19.1
*/
module top();
	typedef enum {a, b, c} e;
	e val;
endmodule
