/*
:name: real
:description: real type tests
:tags: 6.12
*/
module top();
	real a = 0.5;
endmodule
