/*
:name: 22.8--default_nettype
:description: Test
:tags: 22.8
:type: preprocessing
*/
`default_nettype wire
