/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 11499
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_cmn_clks_svt_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wavshared_gf12lp_dig_lib, Cell - wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT,
//View - schematic
// LAST TIME SAVED: Nov 10 10:24:09 2020
// NETLIST TIME: May 26 14:59:42 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT (q, vdd, vss, clk, clkb, d, rst, rstb, 
    tiehi, tielo);

output  q;

inout  vdd, vss;

input  clk, clkb, d, rst, rstb, tiehi, tielo;


wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF0 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd), .rstb(rstb), .d(d), .clkb(clkb), .clk(clk), 
    .q(q_mid));

wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF1 ( .tielo(tielo), .tiehi(tiehi), .rst(rst), 
    .vss(vss), .vdd(vdd), .rstb(rstb), .d(q_mid), .clkb(clkb), 
    .clk(clk), .q(q));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt, View -
//schematic
// LAST TIME SAVED: Dec 29 15:13:54 2020
// NETLIST TIME: May 26 14:59:43 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt (o_clk, o_clk_b, vdd, vss, ena, i_clk, 
    i_clk_b);

output  o_clk, o_clk_b;

inout  vdd, vss;

input  ena, i_clk, i_clk_b;


wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(ckb), .en(en), .enb(enb), .vss(vss), 
    .in(i_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT1 ( .out(ckbb), .en(en), .enb(enb), .vss(vss), 
    .in(i_clk_b), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_PU_D2_GL16_RVT PU0 ( .vdd(vdd), .en(en), .y(ckb));

wphy_lp4x5_cmn_clks_svt_PD_D2_GL16_RVT PD0 ( .vss(vss), .enb(enb), .y(ckbb));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(ena), .vss(vss), .out(net012), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1_1 ( .in(ckb), .vss(vss), .out(o_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1_0 ( .in(ckb), .vss(vss), .out(o_clk), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(enb), .vss(vss), .out(en), .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2_1 ( .in(ckbb), .vss(vss), .out(o_clk_b), 
    .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2_0 ( .in(ckbb), .vss(vss), .out(o_clk_b), 
    .vdd(vdd));

wphy_lp4x5_cmn_clks_svt_PUDUM_D2_GL16_RVT PUDUM ( .vdd(vdd), .tiehi(vdd));

wphy_lp4x5_cmn_clks_svt_PDDUM_D2_GL16_RVT PDDUM ( .vss(vss), .tielo(vss));

wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT LA0 ( .tielo(vss), .vss(vss), .vdd(vdd), .tiehi(vdd), 
    .d(net012), .clkb(i_clk_b), .clk(i_clk), .q(enb));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt,
//View - schematic
// LAST TIME SAVED: Jan 21 22:52:59 2021
// NETLIST TIME: May 26 14:59:43 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt (o_clk0, o_clk90, o_clk180, o_clk270, 
    vdda, vss, i_byp, i_clk0, i_clk180, i_rst);

output  o_clk0, o_clk90, o_clk180, o_clk270;

inout  vdda, vss;

input  i_byp, i_clk0, i_clk180, i_rst;


wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_0 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_1 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_2 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_3 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_4 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_5 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_6 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_7 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_8 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_9 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_10 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_11 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_12 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_13 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_14 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_15 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_16 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_17 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_18 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_19 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_20 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_21 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_22 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_23 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_24 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_25 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_26 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_27 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_28 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_29 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_30 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_31 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_32 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_33 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_34 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_35 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_36 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_37 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_38 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_39 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM0_40 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR0 ( .tielo(vss), .tiehi(vdda), .y(rst_or_byp_n), 
    .vss(vss), .vdd(vdda), .b(i_byp), .a(i_rst));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV16 ( .in(x90), .vss(vss), .out(x270), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV19 ( .in(net021), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV18 ( .in(net029), .vss(vss), .out(o_clk270), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV17 ( .in(net028), .vss(vss), .out(o_clk90), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14 ( .in(x180), .vss(vss), .out(x0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV20 ( .in(net030), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(bypb), .vss(vss), .out(bypa), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(i_byp), .vss(vss), .out(bypb), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15 ( .in(net020), .vss(vss), .out(x90), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2 ( .in(net015), .vss(vss), .out(x180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9 ( .in(rst_or_byp_n), .vss(vss), .out(rst_or_byp), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT I3 ( .out(net028), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT3 ( .out(net021), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT2 ( .out(net021), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT8 ( .out(net028), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x90), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT1 ( .out(net030), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT7 ( .out(net029), .en(bypb), .enb(bypa), 
    .vss(vss), .in(x270), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(net030), .en(bypa), .enb(bypb), 
    .vss(vss), .in(i_clk180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT I4 ( .out(net029), .en(bypa), .enb(bypb), .vss(vss), 
    .in(i_clk0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT0 ( .tiehi(vdda), .tielo(vss), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(net020), .clkb(i_clk0), 
    .clk(i_clk180), .q(net015));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT1 ( .tiehi(vdda), .tielo(vss), .vss(vss), 
    .vdd(vdda), .rstb(rst_or_byp_n), .d(x180), .clkb(i_clk180), 
    .clk(i_clk0), .q(net020));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt, View -
//schematic
// LAST TIME SAVED: May 26 13:50:27 2021
// NETLIST TIME: May 26 14:59:43 2021
`timescale 1ps / 1ps 




 

module wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt (clka_sel, clkb_sel, o_clk0, o_clk180, vdda, vss, 
    clk_sel, ena, i_clka0, i_clka180, i_clkb0, i_clkb180);

output  clka_sel, clkb_sel, o_clk0, o_clk180;

inout  vdda, vss;

input  clk_sel, ena, i_clka0, i_clka180, i_clkb0, i_clkb180;


wphy_lp4x5_cmn_clks_svt_PUDUM_D2_GL16_RVT PUDUM ( .vdd(vdda), .tiehi(vdda));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA1 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net6), .clkb(clka180), .clk(clka0), .q(net023));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA4 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net3), .clkb(clkb180), .clk(clkb0), .q(net022));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA2 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net023), .clkb(clka0), .clk(clka180), .q(net5));

wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT LA3 ( .tielo(vss), .set(enb), .vss(vss), .vdd(vdda), 
    .tiehi(vdda), .d(net022), .clkb(clkb0), .clk(clkb180), .q(net2));

wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT LA02 ( .prst(enb), .prstb(en), .tielo(vss), 
    .vss(vss), .vdd(vdda), .tiehi(vdda), .d(y), .clkb(clkb180), 
    .clk(clkb0), .q(net3));

wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT LA01 ( .prst(enb), .prstb(en), .tielo(vss), 
    .vss(vss), .vdd(vdda), .tiehi(vdda), .d(net4), .clkb(clka180), 
    .clk(clka0), .q(net6));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND2 ( .tielo(vss), .vdd(vdda), .y(pu_en), 
    .vss(vss), .tiehi(vdda), .b(enb_b), .a(enb_a));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND1 ( .tielo(vss), .vdd(vdda), .y(y), .vss(vss), 
    .tiehi(vdda), .b(enb_a), .a(sel_clkb));

wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT NAND0 ( .tielo(vss), .vdd(vdda), .y(net4), .vss(vss), 
    .tiehi(vdda), .b(enb_b), .a(sel_cala));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT0 ( .out(net036), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT5 ( .out(net035), .en(en_a), .enb(enb_a), 
    .vss(vss), .in(clka180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT4 ( .out(net035), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb180), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT INVT3 ( .out(net036), .en(en_b), .enb(enb_b), 
    .vss(vss), .in(clkb0), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LA0 ( .tiehi(vdda), .tielo(vss), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net09), .clkb(clkb180), .clk(clkb0), 
    .q(en_b));

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LA00 ( .tiehi(vdda), .tielo(vss), .vss(vss), 
    .vdd(vdda), .rstb(en), .d(net038), .clkb(clka180), .clk(clka0), 
    .q(en_a));

wphy_lp4x5_cmn_clks_svt_PD_D2_GL16_RVT PD0 ( .vss(vss), .enb(pd_enb), .y(net035));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR0 ( .tielo(vss), .tiehi(vdda), .y(sel_clkb), 
    .vss(vss), .vdd(vdda), .b(enb), .a(clk_selb));

wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT NOR1 ( .tielo(vss), .tiehi(vdda), .y(sel_cala), 
    .vss(vss), .vdd(vdda), .b(enb), .a(sel_clkb));

wphy_lp4x5_cmn_clks_svt_PDDUM_D2_GL16_RVT PDDUM ( .vss(vss), .tielo(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_0 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_1 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_2 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_3 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_4 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_5 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_6 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_7 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_8 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_9 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_10 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_11 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_12 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_13 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_14 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_15 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_16 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_17 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_18 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_19 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_20 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_21 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_22 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_23 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_24 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_25 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_26 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_27 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_28 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_29 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_30 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_31 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_32 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_33 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_34 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_35 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_36 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_37 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_38 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_39 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_40 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_41 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_42 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_43 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_44 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_45 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_46 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_47 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_48 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_49 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_50 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_51 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_52 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_53 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_54 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_55 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_56 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_57 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_58 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_59 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_60 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_61 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_62 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_63 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_64 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_65 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_66 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_67 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_68 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_69 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_70 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_71 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_72 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_73 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_74 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_75 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_76 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_77 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_78 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_79 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_80 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_81 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_82 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_83 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_84 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_85 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_86 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_87 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_88 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_89 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_90 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_91 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_92 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_93 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_94 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_95 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_96 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_97 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_98 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_99 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_100 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_101 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_102 ( .tiehi(vdda), .tielo(vss), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV5 ( .in(enb_b), .vss(vss), .out(clkb_sel), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV4 ( .in(enb_a), .vss(vss), .out(clka_sel), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2 ( .in(enb), .vss(vss), .out(en), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV19 ( .in(pu_en), .vss(vss), .out(pd_enb), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(clk_sel), .vss(vss), .out(clk_selb), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV16 ( .in(en_b), .vss(vss), .out(enb_b), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15_1 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV15_0 ( .in(net050), .vss(vss), .out(clkb180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14_1 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV14_0 ( .in(net034), .vss(vss), .out(clkb0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV13 ( .in(i_clkb0), .vss(vss), .out(net034), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV12 ( .in(i_clkb180), .vss(vss), .out(net050), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV11_1 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV11_0 ( .in(net049), .vss(vss), .out(clka180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV8 ( .in(i_clka0), .vss(vss), .out(net019), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT I1 ( .in(net5), .vss(vss), .out(net038), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(net2), .vss(vss), .out(net09), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(en_a), .vss(vss), .out(enb_a), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7 ( .in(net035), .vss(vss), .out(o_clk180), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV6 ( .in(net036), .vss(vss), .out(o_clk0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV20 ( .in(ena), .vss(vss), .out(enb), .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9_1 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV9_0 ( .in(net019), .vss(vss), .out(clka0), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV10 ( .in(i_clka180), .vss(vss), .out(net049), 
    .vdd(vdda));

wphy_lp4x5_cmn_clks_svt_PU_D2_GL16_RVT PU0 ( .vdd(vdda), .en(pu_en), .y(net036));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cmn_clks_svt,
//View - schematic
// LAST TIME SAVED: Apr  8 15:10:04 2021
// NETLIST TIME: May 26 14:59:43 2021
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_cmn_clks_svt (gfcm0_clka_sel, gfcm0_clkb_sel, 
    gfcm1_clka_sel, gfcm1_clkb_sel, phy_clk0, phy_clk90, phy_clk180, 
    phy_clk270, pll0_div_clk,   gfcm_clksel, gfcm_ena, 
    phy_clk_ena, pll0_div_clk_byp, pll0_div_clk_ena, pll0_div_clk_rst, 
    vco1_clk0, vco1_clk90, vco1_clk180, vco1_clk270, vco2_clk0, 
    vco2_clk90, vco2_clk180, vco2_clk270
`ifdef WLOGIC_NO_PG 
`else  
 ,vdd_phy  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdd_phy;
assign vdd_phy=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdd_phy;
inout vss;
`endif


output  gfcm0_clka_sel, gfcm0_clkb_sel, gfcm1_clka_sel, gfcm1_clkb_sel, 
    phy_clk0, phy_clk90, phy_clk180, phy_clk270, pll0_div_clk;



input  gfcm_clksel, gfcm_ena, phy_clk_ena, pll0_div_clk_byp, 
    pll0_div_clk_ena, pll0_div_clk_rst, vco1_clk0, vco1_clk90, 
    vco1_clk180, vco1_clk270, vco2_clk0, vco2_clk90, vco2_clk180, 
    vco2_clk270;

`ifdef SYNTHESIS
`else 

wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT LAT0 ( .tiehi(vdd_phy), .tielo(vss), .vss(vss), 
    .vdd(vdd_phy), .rstb(rst_n), .d(clk_ena_ff), .clkb(div_clk90), 
    .clk(div_clk270), .q(clk_ena_ff1p5));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV12 ( .in(net6), .vss(vss), .out(net20), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV11 ( .in(net5), .vss(vss), .out(net14), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV6 ( .in(net2), .vss(vss), .out(net9), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV13 ( .in(net3), .vss(vss), .out(net10), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV14 ( .in(net8), .vss(vss), .out(net7), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT INV5 ( .in(net1), .vss(vss), .out(net4), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT FF1 ( .tielo(vss), .tiehi(vdd_phy), .rst(rst), 
    .vss(vss), .vdd(vdd_phy), .rstb(rst_n), .d(phy_clk_ena), 
    .clkb(div_clk180), .clk(div_clk0), .q(net136));

wphy_lp4x5_cmn_clks_svt_FFRES_DEMET_D1_GL16_RVT FF0 ( .tielo(vss), .tiehi(vdd_phy), .rst(rst), 
    .vss(vss), .vdd(vdd_phy), .rstb(rst_n), .d(pll0_div_clk_ena), 
    .clkb(net9), .clk(net4), .q(div_clk_ena_ff));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC2 ( .o_clk(net133), .o_clk_b(net134), 
    .ena(div_clk_ena_ff), .i_clk(net4), .i_clk_b(net9), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC0 ( .o_clk(net6), .o_clk_b(net5), 
    .ena(clk_ena_ff), .i_clk(gfm_clk0), .i_clk_b(gfm_clk180), 
    .vdd(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_cgc_diff_svt CGC1 ( .o_clk(net8), .o_clk_b(net3), 
    .ena(clk_ena_ff1p5), .i_clk(gfm_clk90), .i_clk_b(gfm_clk270), 
    .vdd(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_clk_div2_4g_core_svt IDIV2 ( .o_clk90(div_clk90), 
    .o_clk270(div_clk270), .o_clk0(div_clk0), .o_clk180(div_clk180), 
    .i_byp(pll0_div_clk_byp), .i_clk0(net133), .i_clk180(net134), 
    .i_rst(rst), .vdda(vdd_phy), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt GFCM0 ( .clka_sel(gfcm0_clka_sel), 
    .clkb_sel(gfcm0_clkb_sel), .vdda(vdd_phy), .i_clka0(vco1_clk0), 
    .o_clk0(gfm_clk0), .o_clk180(gfm_clk180), .clk_sel(gfcm_clksel), 
    .i_clka180(vco1_clk180), .i_clkb0(vco2_clk0), 
    .i_clkb180(vco2_clk180), .ena(gfcm_ena), .vss(vss));

wphy_lp4x5_cmn_clks_svt_wphy_gfcm_svt GFCM1 ( .clka_sel(gfcm1_clka_sel), 
    .clkb_sel(gfcm1_clkb_sel), .vdda(vdd_phy), .i_clka0(vco1_clk90), 
    .o_clk0(gfm_clk90), .o_clk180(gfm_clk270), .clk_sel(gfcm_clksel), 
    .i_clka180(vco1_clk270), .i_clkb0(vco2_clk90), 
    .i_clkb180(vco2_clk270), .ena(gfcm_ena), .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUMLOAD_D2_GL16_RVT I9 ( .vdd(vdd_phy), .inn(gfm_clk90), .vss(vss), 
    .inp(gfm_clk90));

wphy_lp4x5_cmn_clks_svt_DUMLOAD_D2_GL16_RVT I8 ( .vdd(vdd_phy), .inn(gfm_clk270), .vss(vss), 
    .inp(gfm_clk270));

wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT I5 ( .in(net20), .vss(vss), .out(phy_clk0), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT I4 ( .in(net14), .vss(vss), .out(phy_clk180), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT I6 ( .in(net10), .vss(vss), .out(phy_clk270), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT I7 ( .in(net7), .vss(vss), .out(phy_clk90), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV8 ( .in(gfm_clk180), .vss(vss), .out(net2), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7_1 ( .in(div_clk180), .vss(vss), 
    .out(pll0_div_clk), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV7_0 ( .in(div_clk180), .vss(vss), 
    .out(pll0_div_clk), .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV3 ( .in(net136), .vss(vss), .out(net135), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV4 ( .in(net135), .vss(vss), .out(clk_ena_ff), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV2 ( .in(gfm_clk0), .vss(vss), .out(net1), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV1 ( .in(rst_n), .vss(vss), .out(rst), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT INV0 ( .in(pll0_div_clk_rst), .vss(vss), .out(rst_n), 
    .vdd(vdd_phy));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_0 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_1 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_2 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_3 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_4 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_5 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_6 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_7 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_8 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_9 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_10 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_11 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_12 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_13 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_14 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_15 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_16 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_17 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_18 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_19 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_20 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_21 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_22 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_23 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_24 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_25 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_26 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_27 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_28 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_29 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_30 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_31 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_32 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_33 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_34 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_35 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_36 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_37 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_38 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_39 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_40 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_41 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_42 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_43 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_44 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_45 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_46 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_47 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_48 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_49 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_50 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_51 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_52 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_53 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_54 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_55 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_56 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_57 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_58 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_59 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_60 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_61 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_62 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_63 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_64 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_65 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_66 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_67 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_68 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_69 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_70 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_71 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_72 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_73 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_74 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_75 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_76 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_77 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_78 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_79 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_80 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_81 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_82 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_83 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_84 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_85 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_86 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_87 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_88 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_89 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_90 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_91 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_92 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_93 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_94 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_95 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_96 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_97 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_98 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_99 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_100 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_101 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_102 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_103 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_104 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_105 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_106 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_107 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_108 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_109 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_110 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_111 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_112 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_113 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_114 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_115 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_116 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_117 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_118 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_119 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_120 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_121 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_122 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_123 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_124 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_125 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_126 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_127 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_128 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_129 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_130 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_131 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_132 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_133 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_134 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_135 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_136 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_137 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_138 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_139 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_140 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_141 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_142 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_143 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_144 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_145 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_146 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_147 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_148 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_149 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_150 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_151 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_152 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_153 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_154 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT DUM_155 ( .tiehi(vdd_phy), .tielo(vss), .vdd(vdd_phy), 
    .vss(vss));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell -
//wphy_lp4x5_cmn_clks_svt_tb, View - schematic
// LAST TIME SAVED: Dec  7 22:24:21 2020
// NETLIST TIME: May 26 14:59:43 2021
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INV_D8_GL16_RVT ( in,  out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "DUMLOAD_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_DUMLOAD_D2_GL16_RVT ( inp, inn
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input inp;
  input inn;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule



module wphy_lp4x5_cmn_clks_svt_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_clks_svt_FFSET_D1_GL16_RVT( q, clk, clkb, d, prst, prstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input clk;
  input prst;
  input prstb;
  output q;
  input d;
  input clkb;  
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  initial  begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  initial  begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  reg q;

  initial begin
    q = $random;
  end

  always @(posedge clk or posedge prst) begin
   if(prst) begin
       q <= 1'b1;
    end else begin
       q <= d;
    end
  end

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_cmn_clks_svt_LATSET_D1_GL16_RVT ( q, clk, clkb, d, set
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  output q;
  input set;
  input d;
  input clk;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ?
                           (set) ?
                                 1'b1
                                 : (clkb) ?
                                          (d===1'bx) ? $random : d
                                          : q
                           : 1'bx;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//systemVerilog HDL for "wavshared_gf12lp_dig_lib", "wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_DUM_D1_GL16_RVT ( tielo, tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG

 );

  input tiehi;
  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT" "systemVerilog"

`timescale 1ps/1ps
module wphy_lp4x5_cmn_clks_svt_LAT_D1_GL16_RVT( q, clk, clkb, d
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
);
 
  input clk;
  output q;  
  input d;
  input clkb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG


  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;

  assign q = (power_ok) ? 1'bz : 1'bx;
  
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ?
                           (clkb) ?
                                  (d===1'bx) ? $random : d
                                  : q
                           : 1'bx;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PDDUM_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_PDDUM_D2_GL16_RVT (  tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PUDUM_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_PUDUM_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PD_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_PD_D2_GL16_RVT ( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_PU_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_PU_D2_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INVT_D2_GL16_RVT( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT" "systemVerilog"

module wphy_lp4x5_cmn_clks_svt_FFRES_D1_GL16_RVT( q, clk, clkb, d, rst, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input clk;
  input rst;
  input rstb;
  output q;
  input d;
  input clkb;  
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  reg q;

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;

  initial  begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (signals_ok) ? 1'bz : 1'bx;
  end
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd ;
  
  initial  begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
  always @(*) begin
       q = (power_ok) ? 1'bz : 1'bx;
  end
`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  initial begin
    q = $random;
  end

  always @(posedge clk or posedge rst) begin
   if(rst) begin
       q <= 1'b0;
    end else begin
       q <= d;
    end
  end

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cmn_clks_svt_INV_D4_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;


endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "LATRES_D1_GL16_LVT" "systemVerilog"


`timescale 1ps/1ps
module wphy_lp4x5_cmn_clks_svt_LATRES_D1_GL16_RVT( q, clk, clkb, d, rstb
`ifdef WLOGIC_MODEL_NO_TIE
`else
, tiehi, tielo 
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PGL
);

  input clk;
  output q;
  input d;
  input clkb;
  input rstb;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire #0 polarity_ok = clk^clkb;

`ifdef WLOGIC_MODEL_NO_TIE
`else
  wire signals_ok;
  assign signals_ok = tiehi & ~tielo ;

  assign q = (signals_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign q = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


assign #1  q = polarity_ok ? 
                           (~rstb) ? 
                                 1'b0 
                                 : (clkb) ? 
                                          (d===1'bx) ? $random : d&rstb
                                          : q 
                           : 1'bx;

endmodule

`endif //SYNTHESIS
