/*
:name: preproc_test_2
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`include "preproc_test_2.svh"
`ifndef SUCCESS
Didn't successfully include preproc_test_2.svh!
`endif
`ifndef SANITY
`define SANITY
`endif
