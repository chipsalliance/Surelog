/*
:name: class_member_test_43
:description: Test
:tags: 8.3
*/
class constructible;
function new (foo::bar name,
    virtual interface time_if vif,
    baz#(M,N)::foo bar, bit [K:0] b);
  this.name = name;
endfunction
endclass