/*
:name: preproc_test_11
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`define LONG_MACRO(\
    a,\
    b\
, c\
) \
more text c, b, a \
blah blah macro ends here
