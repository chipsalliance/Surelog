/*
:name: typedef_test_4
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef enum { RED, GREEN, BLUE } colors;