

module mod3();


NO_DEF_6 nodef6();

endmodule
