module top;
   localparam int P [2] = '{11, 12};
endmodule // top
