/*
:name: class_test_54
:description: Test
:tags: 6.15 8.3
*/
class event_calendar;
  event birthday;
  event first_date, anniversary;
  event revolution[4:0], independence[2:0];
endclass