`ifdef SURELOG

module top();

endmodule

`endif
