package pkg1;

  typedef enum {
    HERE
  } enum1;

endpackage
