/*
:name: 22.5.1--define_expansion_19
:description: Test
:should_fail: 0
:tags: 22.5.1
:type: preprocessing
*/
`define wordsize 8
module top ();
logic [1:`wordsize] data;
endmodule
