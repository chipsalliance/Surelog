
module def ();
parameter SIZE1 = 2;

defparam small_top.u1.SIZE = SIZE1;

defparam small_top.u1.dummy = 4;
endmodule
