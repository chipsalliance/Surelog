/*
:name: final
:description: final check
:tags: 9.2.3
*/
module initial_tb ();
	reg a = 0;
	final
		a = 1;
endmodule
