/*
:name: class_member_test_1
:description: Test
:tags: 8.3
*/
class c;
  task intf.task1();
  endtask
endclass