/*
:name: class_member_test_4
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern virtual task subtask(arg_type arg);
endclass