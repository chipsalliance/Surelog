module DUT (input wire i, output wire o);
  assign o = i;
endmodule
