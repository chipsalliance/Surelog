/*
:name: enum_anon
:description: anonymous enum tests
:tags: 6.19
*/
module top();
	enum {a, b, c} val;
endmodule
