/*
:name: 22.12--line-illegal-2
:description: The filename parameter shall be a string literal
:should_fail: 1
:tags: 22.12
:type: preprocessing
*/
`line 1 somefile 2
