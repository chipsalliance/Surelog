/*
:name: cont_assignment
:description: continuous assignment test
:tags: 10.3.2
*/
module top(input a, input b);

wire w;
assign w = a & b;

endmodule
