/*
:name: 22.8--default_nettype
:description: Test
:should_fail: 0
:tags: 22.8
:type: preprocessing
*/
`default_nettype wire
