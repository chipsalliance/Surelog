/*
:name: 22.9--unconnected_drive-invalid-1
:description: Test
:should_fail: 1
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive
`nounconnected_drive
