package top1_1;








`include "middle.v"












`include "middle.v"









endpackage


`include "mod.v"


/*
top1
*/

module top_43 ();
endmodule

`include "middle.v"


module bottom_49 ();
endmodule

/*
top2
*/