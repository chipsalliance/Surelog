module dut ;
 logic [63:0]
        o06;
       assign o06 = 3'('1);                                                                   
endmodule
