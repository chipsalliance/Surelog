module dut;

  function automatic int get_expected_command (int slave_id);
     int write_command_queue_slave [10];
  
     foreach (write_command_queue_slave[slave_id,i]) begin
     end
 endfunction

endmodule


