 module test_wand_wor(); 

   wand a;
   wor  b;
   reg c, d; 

   assign a = c;
   assign b = d;   

 endmodule
