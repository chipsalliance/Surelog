/*
:name: 22.12--line-basic
:description: Test
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 2
