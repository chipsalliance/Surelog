/*
:name: info_task
:description: $info test
:tags: 20.10
:type: simulation parsing
*/

module top();

initial begin
	$info("info");
end

endmodule
