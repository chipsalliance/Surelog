// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: arrays-key-index
:description: Basic arrays test
:tags: 5.11
*/
module top();
  typedef int triple [1:3];
  triple b = '{1:1, default:0};
endmodule
