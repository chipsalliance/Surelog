/*
:name: stop_task
:description: $stop test
:tags: 20.2
*/
module top();

initial
	$stop;

endmodule
