module top( input   type_scr1_mem_resp_e                dmem2exu_resp_i);

type_scr1_mem_resp_e                dmem2exu_resp_ii;

endmodule
