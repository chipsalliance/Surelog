/*
:name: class_member_test_38
:description: Test
:tags: 8.3
*/
class myclass;
virtual function virtual array_if.modport_x subroutine();
endfunction
endclass