`define DDR_ANA_PI_MATCH_RSV_RANGE             5:0
`define DDR_ANA_PI_MATCH_GEAR_RANGE            9:6
`define DDR_ANA_PI_MATCH_XCPL_RANGE            13:10
`define DDR_ANA_PI_MATCH_EN_RANGE              14

`define DDR_ANA_PI_MATCH_RANGE                 14:0
