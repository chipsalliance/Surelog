`ifndef TNOC_BFM_STATUS_SVH
`define TNOC_BFM_STATUS_SVH
typedef tue_status_dummy  tnoc_bfm_status;
`endif
