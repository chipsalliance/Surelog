/*
:name: preproc_test_1
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`define FOO BAR-1
