module dut (/*output logic[80:0] a, output logic[80:0] b*/);
   assign a =    147573952589676412928;
   assign b = 'sd147573952589676412928;
   assign c =     18446744073709551615; // 2^64
   assign d =     18446744073709551616; // 2^64 + 1
   assign e =    -18446744073709551616; // 2^64 + 1

endmodule
