// $Id: base_compatibility.svh,v 1.3 2007/12/21 12:49:44 jlrose Exp $
//----------------------------------------------------------------------
//   Copyright 2007-2009 Mentor Graphics Corporation
//   Copyright 2007-2009 Cadence Design Systems, Inc.
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------
`ifndef BASE_COMPATIBILITY_SVH
`define BASE_COMPATIBILITY_SVH

`include "compatibility/urm_macro_compatibility.svh"
`include "compatibility/urm_message_defines.svh"
`include "compatibility/urm_type_compatibility.svh"

`endif //BASE_COMPATIBILITY_SVH

