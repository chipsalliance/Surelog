nettype real my_real;

module dut ();

    my_real my_real_net;

endmodule
