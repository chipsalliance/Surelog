/*
:name: class_test_49
:description: Test
:tags: 6.15 8.3
*/
class params_as_class_item;
  parameter N = 2;
  parameter reg P = '1;
  localparam M = f(glb::arr[N]) + 1;
endclass