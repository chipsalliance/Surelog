/*
:name: finish_task
:description: $finish test
:tags: 20.2
*/
module top();

initial
	$finish;

endmodule
