/*
:name: desc_test_13
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
package foo_pkg;
endpackage
`ifdef F00
`MACRO(stuff)
`endif
