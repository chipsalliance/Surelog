/*
:name: include-directive
:description: Include empty file
:should_fail: 0
:tags: 5.6.4
*/

`include "/dev/null"

module empty();
endmodule
