/*
:name: var_protected
:description: class with protected variable
:tags: 8.18
*/
module class_tb ();
	class a_cls;
		protected int a_prot = 2;
	endclass
endmodule
