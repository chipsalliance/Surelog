 module top;
   logic [31:0] a = 'Z;
   logic [31:0] b = 'X;
   logic [31:0] c = '0;
   logic [31:0] d = '1;
endmodule // top

