// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: attributes-module
:description: Assing attributes to a module
:tags: 5.12
*/

(* optimize_power *)
module topa();
endmodule

(* optimize_power=0 *)
module topb();
endmodule

(* optimize_power=1 *)
module topc();
endmodule
