/*
:name: 22.5.2--undef-nonexisting
:description: Test
:tags: 22.5.2
:type: preprocessing
*/
`undef FOO
`undef BAR
