// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: basic-packed
:description: Test packed arrays support
:tags: 7.4.1 7.4
*/
module top ();

bit [7:0] _bit;
logic [7:0] _logic;
reg [7:0] _reg;

endmodule
