`define DDR_ANA_SA_4PH_CAL_CODE_0_RANGE            3:0
`define DDR_ANA_SA_4PH_CAL_CODE_90_RANGE           7:4
`define DDR_ANA_SA_4PH_CAL_CODE_180_RANGE         11:8
`define DDR_ANA_SA_4PH_CAL_CODE_270_RANGE         15:12
`define DDR_ANA_SA_4PH_CAL_DIR_0_RANGE               16
`define DDR_ANA_SA_4PH_CAL_DIR_90_RANGE              17
`define DDR_ANA_SA_4PH_CAL_DIR_180_RANGE             18
`define DDR_ANA_SA_4PH_CAL_DIR_270_RANGE             19
