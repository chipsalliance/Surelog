/*
:name: class_test_40
:description: Test
:tags: 6.15 8.3
*/
class macros_as_class_item;
 `uvm_object_registry(myclass, "class_name")
endclass