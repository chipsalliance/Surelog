/*
:name: class_test_14
:description: Test
:tags: 6.15 8.3
*/
class Foo #(T=int);
endclass