/*
:name: class_member_test_47
:description: Test
:tags: 8.3
*/
class fun_with_typedef_members;
typedef struct { int i; bool b; } mystruct;
typedef enum { RED, GREEN, BLUE } colors;
typedef virtual blah_if harness_if;
typedef virtual interface blah_if harness_if;
typedef virtual blah_if#(N) foo_if;
typedef virtual blah_if#(N).modport_id foo_if;
endclass