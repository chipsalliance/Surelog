/*
:name: integers-token
:description: Testing the integer variable type
:tags: 5.7.1
*/
module top();
  integer a;
endmodule
