
module top;
   if (1) begin
    assign a = b;
   end
   else begin
    assign c = d;
   end
endmodule