/*
:name: basic-unpacked
:description: Test unpacked arrays support
:tags: 7.4.2 7.4
*/
module top ();

bit _bit [7:0];
logic _logic [7:0];
reg _reg [7:0];

endmodule
