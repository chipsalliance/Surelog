/*
:name: typedef_test_2
:description: Test
:tags: 6.18
*/
typedef reg quartet[3:0];