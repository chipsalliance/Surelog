//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_arbitrator (
                                          // inputs:
                                           clk,
                                           cpu_jtag_debug_module_readdata,
                                           cpu_jtag_debug_module_resetrequest,
                                           pipeline_bridge_m1_address_to_slave,
                                           pipeline_bridge_m1_burstcount,
                                           pipeline_bridge_m1_byteenable,
                                           pipeline_bridge_m1_chipselect,
                                           pipeline_bridge_m1_debugaccess,
                                           pipeline_bridge_m1_latency_counter,
                                           pipeline_bridge_m1_read,
                                           pipeline_bridge_m1_write,
                                           pipeline_bridge_m1_writedata,
                                           reset_n,

                                          // outputs:
                                           cpu_jtag_debug_module_address,
                                           cpu_jtag_debug_module_begintransfer,
                                           cpu_jtag_debug_module_byteenable,
                                           cpu_jtag_debug_module_chipselect,
                                           cpu_jtag_debug_module_debugaccess,
                                           cpu_jtag_debug_module_readdata_from_sa,
                                           cpu_jtag_debug_module_reset_n,
                                           cpu_jtag_debug_module_resetrequest_from_sa,
                                           cpu_jtag_debug_module_write,
                                           cpu_jtag_debug_module_writedata,
                                           d1_cpu_jtag_debug_module_end_xfer,
                                           pipeline_bridge_m1_granted_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
                                           pipeline_bridge_m1_requests_cpu_jtag_debug_module
                                        )
;

  output  [  8: 0] cpu_jtag_debug_module_address;
  output           cpu_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_jtag_debug_module_byteenable;
  output           cpu_jtag_debug_module_chipselect;
  output           cpu_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  output           cpu_jtag_debug_module_reset_n;
  output           cpu_jtag_debug_module_resetrequest_from_sa;
  output           cpu_jtag_debug_module_write;
  output  [ 31: 0] cpu_jtag_debug_module_writedata;
  output           d1_cpu_jtag_debug_module_end_xfer;
  output           pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  output           pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata;
  input            cpu_jtag_debug_module_resetrequest;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_debugaccess;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_allgrants;
  wire             cpu_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_jtag_debug_module_any_continuerequest;
  wire             cpu_jtag_debug_module_arb_counter_enable;
  reg              cpu_jtag_debug_module_arb_share_counter;
  wire             cpu_jtag_debug_module_arb_share_counter_next_value;
  wire             cpu_jtag_debug_module_arb_share_set_values;
  wire             cpu_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_jtag_debug_module_begins_xfer;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire             cpu_jtag_debug_module_end_xfer;
  wire             cpu_jtag_debug_module_firsttransfer;
  wire             cpu_jtag_debug_module_grant_vector;
  wire             cpu_jtag_debug_module_in_a_read_cycle;
  wire             cpu_jtag_debug_module_in_a_write_cycle;
  wire             cpu_jtag_debug_module_master_qreq_vector;
  wire             cpu_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  reg              cpu_jtag_debug_module_reg_firsttransfer;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  reg              cpu_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_jtag_debug_module_waits_for_read;
  wire             cpu_jtag_debug_module_waits_for_write;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  reg              d1_cpu_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module;
  wire    [ 11: 0] shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1;
  wire             wait_for_cpu_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_jtag_debug_module_end_xfer;
    end


  assign cpu_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module));
  //assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata;

  assign pipeline_bridge_m1_requests_cpu_jtag_debug_module = ({pipeline_bridge_m1_address_to_slave[11] , 11'b0} == 12'h0) & pipeline_bridge_m1_chipselect;
  //cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_jtag_debug_module_arb_share_set_values = 1;

  //cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_jtag_debug_module_non_bursting_master_requests = pipeline_bridge_m1_requests_cpu_jtag_debug_module;

  //cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_jtag_debug_module_arb_share_counter_next_value = cpu_jtag_debug_module_firsttransfer ? (cpu_jtag_debug_module_arb_share_set_values - 1) : |cpu_jtag_debug_module_arb_share_counter ? (cpu_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_jtag_debug_module_allgrants = |cpu_jtag_debug_module_grant_vector;

  //cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_jtag_debug_module_end_xfer = ~(cpu_jtag_debug_module_waits_for_read | cpu_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_jtag_debug_module = cpu_jtag_debug_module_end_xfer & (~cpu_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & cpu_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests);

  //cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_jtag_debug_module_arb_counter_enable)
          cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_jtag_debug_module & ~cpu_jtag_debug_module_non_bursting_master_requests))
          cpu_jtag_debug_module_slavearbiterlockenable <= |cpu_jtag_debug_module_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = cpu_jtag_debug_module_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_jtag_debug_module_slavearbiterlockenable2 = |cpu_jtag_debug_module_arb_share_counter_next_value;

  //pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = cpu_jtag_debug_module_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_assign
  assign cpu_jtag_debug_module_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module = pipeline_bridge_m1_requests_cpu_jtag_debug_module & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~cpu_jtag_debug_module_waits_for_read;

  //cpu_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_jtag_debug_module_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_cpu_jtag_debug_module = pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;

  //pipeline_bridge/m1 saved-grant cpu/jtag_debug_module, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module = pipeline_bridge_m1_requests_cpu_jtag_debug_module;

  //allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  assign cpu_jtag_debug_module_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign cpu_jtag_debug_module_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign cpu_jtag_debug_module_master_qreq_vector = 1;

  assign cpu_jtag_debug_module_begintransfer = cpu_jtag_debug_module_begins_xfer;
  //cpu_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_jtag_debug_module_reset_n = reset_n;

  //assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest;

  assign cpu_jtag_debug_module_chipselect = pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  //cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_firsttransfer = cpu_jtag_debug_module_begins_xfer ? cpu_jtag_debug_module_unreg_firsttransfer : cpu_jtag_debug_module_reg_firsttransfer;

  //cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_jtag_debug_module_unreg_firsttransfer = ~(cpu_jtag_debug_module_slavearbiterlockenable & cpu_jtag_debug_module_any_continuerequest);

  //cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_jtag_debug_module_begins_xfer)
          cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_jtag_debug_module_beginbursttransfer_internal = cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_jtag_debug_module_write = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //cpu_jtag_debug_module_address mux, which is an e_mux
  assign cpu_jtag_debug_module_address = shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 >> 2;

  //d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end


  //cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_read = cpu_jtag_debug_module_in_a_read_cycle & cpu_jtag_debug_module_begins_xfer;

  //cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_read_cycle = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_jtag_debug_module_in_a_read_cycle;

  //cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_jtag_debug_module_waits_for_write = cpu_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_jtag_debug_module_in_a_write_cycle = pipeline_bridge_m1_granted_cpu_jtag_debug_module & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_jtag_debug_module_counter = 0;
  //cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_jtag_debug_module_byteenable = (pipeline_bridge_m1_granted_cpu_jtag_debug_module)? pipeline_bridge_m1_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_jtag_debug_module_debugaccess = (pipeline_bridge_m1_granted_cpu_jtag_debug_module)? pipeline_bridge_m1_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_cpu_jtag_debug_module && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_data_master_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_data_master_address,
                                     cpu_data_master_burstcount,
                                     cpu_data_master_byteenable,
                                     cpu_data_master_granted_custom_dma_burst_0_upstream,
                                     cpu_data_master_granted_custom_dma_burst_2_upstream,
                                     cpu_data_master_granted_custom_dma_burst_4_upstream,
                                     cpu_data_master_qualified_request_custom_dma_burst_0_upstream,
                                     cpu_data_master_qualified_request_custom_dma_burst_2_upstream,
                                     cpu_data_master_qualified_request_custom_dma_burst_4_upstream,
                                     cpu_data_master_read,
                                     cpu_data_master_read_data_valid_custom_dma_burst_0_upstream,
                                     cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register,
                                     cpu_data_master_read_data_valid_custom_dma_burst_2_upstream,
                                     cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register,
                                     cpu_data_master_read_data_valid_custom_dma_burst_4_upstream,
                                     cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register,
                                     cpu_data_master_requests_custom_dma_burst_0_upstream,
                                     cpu_data_master_requests_custom_dma_burst_2_upstream,
                                     cpu_data_master_requests_custom_dma_burst_4_upstream,
                                     cpu_data_master_write,
                                     cpu_data_master_writedata,
                                     custom_dma_burst_0_upstream_readdata_from_sa,
                                     custom_dma_burst_0_upstream_waitrequest_from_sa,
                                     custom_dma_burst_2_upstream_readdata_from_sa,
                                     custom_dma_burst_2_upstream_waitrequest_from_sa,
                                     custom_dma_burst_4_upstream_readdata_from_sa,
                                     custom_dma_burst_4_upstream_waitrequest_from_sa,
                                     d1_custom_dma_burst_0_upstream_end_xfer,
                                     d1_custom_dma_burst_2_upstream_end_xfer,
                                     d1_custom_dma_burst_4_upstream_end_xfer,
                                     fir_dma_control_irq_from_sa,
                                     jtag_uart_avalon_jtag_slave_irq_from_sa,
                                     reset_n,
                                     timestamp_timer_s1_irq_from_sa,

                                    // outputs:
                                     cpu_data_master_address_to_slave,
                                     cpu_data_master_irq,
                                     cpu_data_master_latency_counter,
                                     cpu_data_master_readdata,
                                     cpu_data_master_readdatavalid,
                                     cpu_data_master_waitrequest
                                  )
;

  output  [ 26: 0] cpu_data_master_address_to_slave;
  output  [ 31: 0] cpu_data_master_irq;
  output           cpu_data_master_latency_counter;
  output  [ 31: 0] cpu_data_master_readdata;
  output           cpu_data_master_readdatavalid;
  output           cpu_data_master_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_data_master_address;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_granted_custom_dma_burst_0_upstream;
  input            cpu_data_master_granted_custom_dma_burst_2_upstream;
  input            cpu_data_master_granted_custom_dma_burst_4_upstream;
  input            cpu_data_master_qualified_request_custom_dma_burst_0_upstream;
  input            cpu_data_master_qualified_request_custom_dma_burst_2_upstream;
  input            cpu_data_master_qualified_request_custom_dma_burst_4_upstream;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_custom_dma_burst_0_upstream;
  input            cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  input            cpu_data_master_read_data_valid_custom_dma_burst_2_upstream;
  input            cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  input            cpu_data_master_read_data_valid_custom_dma_burst_4_upstream;
  input            cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  input            cpu_data_master_requests_custom_dma_burst_0_upstream;
  input            cpu_data_master_requests_custom_dma_burst_2_upstream;
  input            cpu_data_master_requests_custom_dma_burst_4_upstream;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] custom_dma_burst_0_upstream_readdata_from_sa;
  input            custom_dma_burst_0_upstream_waitrequest_from_sa;
  input   [ 31: 0] custom_dma_burst_2_upstream_readdata_from_sa;
  input            custom_dma_burst_2_upstream_waitrequest_from_sa;
  input   [ 31: 0] custom_dma_burst_4_upstream_readdata_from_sa;
  input            custom_dma_burst_4_upstream_waitrequest_from_sa;
  input            d1_custom_dma_burst_0_upstream_end_xfer;
  input            d1_custom_dma_burst_2_upstream_end_xfer;
  input            d1_custom_dma_burst_4_upstream_end_xfer;
  input            fir_dma_control_irq_from_sa;
  input            jtag_uart_avalon_jtag_slave_irq_from_sa;
  input            reset_n;
  input            timestamp_timer_s1_irq_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_data_master_address_last_time;
  wire    [ 26: 0] cpu_data_master_address_to_slave;
  reg     [  3: 0] cpu_data_master_burstcount_last_time;
  reg     [  3: 0] cpu_data_master_byteenable_last_time;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_is_granted_some_slave;
  reg              cpu_data_master_latency_counter;
  reg              cpu_data_master_read_but_no_slave_selected;
  reg              cpu_data_master_read_last_time;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_run;
  wire             cpu_data_master_waitrequest;
  reg              cpu_data_master_write_last_time;
  reg     [ 31: 0] cpu_data_master_writedata_last_time;
  wire             latency_load_value;
  wire             p1_cpu_data_master_latency_counter;
  wire             pre_flush_cpu_data_master_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_data_master_qualified_request_custom_dma_burst_0_upstream | ~cpu_data_master_requests_custom_dma_burst_0_upstream) & ((~cpu_data_master_qualified_request_custom_dma_burst_0_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_0_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_custom_dma_burst_0_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_0_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_custom_dma_burst_2_upstream | ~cpu_data_master_requests_custom_dma_burst_2_upstream) & ((~cpu_data_master_qualified_request_custom_dma_burst_2_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_2_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_custom_dma_burst_2_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_2_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & 1 & (cpu_data_master_qualified_request_custom_dma_burst_4_upstream | ~cpu_data_master_requests_custom_dma_burst_4_upstream) & ((~cpu_data_master_qualified_request_custom_dma_burst_4_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_4_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write)))) & ((~cpu_data_master_qualified_request_custom_dma_burst_4_upstream | ~(cpu_data_master_read | cpu_data_master_write) | (1 & ~custom_dma_burst_4_upstream_waitrequest_from_sa & (cpu_data_master_read | cpu_data_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_data_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_data_master_address_to_slave = cpu_data_master_address[26 : 0];

  //cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_data_master_read_but_no_slave_selected <= cpu_data_master_read & cpu_data_master_run & ~cpu_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_data_master_is_granted_some_slave = cpu_data_master_granted_custom_dma_burst_0_upstream |
    cpu_data_master_granted_custom_dma_burst_2_upstream |
    cpu_data_master_granted_custom_dma_burst_4_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_data_master_readdatavalid = cpu_data_master_read_data_valid_custom_dma_burst_0_upstream |
    cpu_data_master_read_data_valid_custom_dma_burst_2_upstream |
    cpu_data_master_read_data_valid_custom_dma_burst_4_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_data_master_readdatavalid = cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid |
    cpu_data_master_read_but_no_slave_selected |
    pre_flush_cpu_data_master_readdatavalid;

  //cpu/data_master readdata mux, which is an e_mux
  assign cpu_data_master_readdata = ({32 {~cpu_data_master_read_data_valid_custom_dma_burst_0_upstream}} | custom_dma_burst_0_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_custom_dma_burst_2_upstream}} | custom_dma_burst_2_upstream_readdata_from_sa) &
    ({32 {~cpu_data_master_read_data_valid_custom_dma_burst_4_upstream}} | custom_dma_burst_4_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_data_master_waitrequest = ~cpu_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_latency_counter <= 0;
      else 
        cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_data_master_latency_counter = ((cpu_data_master_run & cpu_data_master_read))? latency_load_value :
    (cpu_data_master_latency_counter)? cpu_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //irq assign, which is an e_assign
  assign cpu_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    fir_dma_control_irq_from_sa,
    jtag_uart_avalon_jtag_slave_irq_from_sa,
    timestamp_timer_s1_irq_from_sa};


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_address_last_time <= 0;
      else 
        cpu_data_master_address_last_time <= cpu_data_master_address;
    end


  //cpu/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_data_master_waitrequest & (cpu_data_master_read | cpu_data_master_write);
    end


  //cpu_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_address != cpu_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_burstcount_last_time <= 0;
      else 
        cpu_data_master_burstcount_last_time <= cpu_data_master_burstcount;
    end


  //cpu_data_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_burstcount != cpu_data_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_data_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_byteenable_last_time <= 0;
      else 
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
    end


  //cpu_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_byteenable != cpu_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_read_last_time <= 0;
      else 
        cpu_data_master_read_last_time <= cpu_data_master_read;
    end


  //cpu_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_read != cpu_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_write_last_time <= 0;
      else 
        cpu_data_master_write_last_time <= cpu_data_master_write;
    end


  //cpu_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_write != cpu_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_data_master_writedata_last_time <= 0;
      else 
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
    end


  //cpu_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_data_master_writedata != cpu_data_master_writedata_last_time) & cpu_data_master_write)
        begin
          $write("%0d ns: cpu_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_instruction_master_arbitrator (
                                           // inputs:
                                            clk,
                                            cpu_instruction_master_address,
                                            cpu_instruction_master_burstcount,
                                            cpu_instruction_master_granted_custom_dma_burst_1_upstream,
                                            cpu_instruction_master_granted_custom_dma_burst_3_upstream,
                                            cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream,
                                            cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream,
                                            cpu_instruction_master_read,
                                            cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream,
                                            cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register,
                                            cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream,
                                            cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register,
                                            cpu_instruction_master_requests_custom_dma_burst_1_upstream,
                                            cpu_instruction_master_requests_custom_dma_burst_3_upstream,
                                            custom_dma_burst_1_upstream_readdata_from_sa,
                                            custom_dma_burst_1_upstream_waitrequest_from_sa,
                                            custom_dma_burst_3_upstream_readdata_from_sa,
                                            custom_dma_burst_3_upstream_waitrequest_from_sa,
                                            d1_custom_dma_burst_1_upstream_end_xfer,
                                            d1_custom_dma_burst_3_upstream_end_xfer,
                                            reset_n,

                                           // outputs:
                                            cpu_instruction_master_address_to_slave,
                                            cpu_instruction_master_latency_counter,
                                            cpu_instruction_master_readdata,
                                            cpu_instruction_master_readdatavalid,
                                            cpu_instruction_master_waitrequest
                                         )
;

  output  [ 26: 0] cpu_instruction_master_address_to_slave;
  output           cpu_instruction_master_latency_counter;
  output  [ 31: 0] cpu_instruction_master_readdata;
  output           cpu_instruction_master_readdatavalid;
  output           cpu_instruction_master_waitrequest;
  input            clk;
  input   [ 26: 0] cpu_instruction_master_address;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_granted_custom_dma_burst_1_upstream;
  input            cpu_instruction_master_granted_custom_dma_burst_3_upstream;
  input            cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream;
  input            cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register;
  input            cpu_instruction_master_requests_custom_dma_burst_1_upstream;
  input            cpu_instruction_master_requests_custom_dma_burst_3_upstream;
  input   [ 31: 0] custom_dma_burst_1_upstream_readdata_from_sa;
  input            custom_dma_burst_1_upstream_waitrequest_from_sa;
  input   [ 31: 0] custom_dma_burst_3_upstream_readdata_from_sa;
  input            custom_dma_burst_3_upstream_waitrequest_from_sa;
  input            d1_custom_dma_burst_1_upstream_end_xfer;
  input            d1_custom_dma_burst_3_upstream_end_xfer;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 26: 0] cpu_instruction_master_address_last_time;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  reg     [  3: 0] cpu_instruction_master_burstcount_last_time;
  wire             cpu_instruction_master_is_granted_some_slave;
  reg              cpu_instruction_master_latency_counter;
  reg              cpu_instruction_master_read_but_no_slave_selected;
  reg              cpu_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_run;
  wire             cpu_instruction_master_waitrequest;
  wire             latency_load_value;
  wire             p1_cpu_instruction_master_latency_counter;
  wire             pre_flush_cpu_instruction_master_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream | ~cpu_instruction_master_requests_custom_dma_burst_1_upstream) & ((~cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream | ~(cpu_instruction_master_read) | (1 & ~custom_dma_burst_1_upstream_waitrequest_from_sa & (cpu_instruction_master_read)))) & 1 & (cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream | ~cpu_instruction_master_requests_custom_dma_burst_3_upstream) & ((~cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream | ~(cpu_instruction_master_read) | (1 & ~custom_dma_burst_3_upstream_waitrequest_from_sa & (cpu_instruction_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign cpu_instruction_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_instruction_master_address_to_slave = cpu_instruction_master_address[26 : 0];

  //cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_instruction_master_read_but_no_slave_selected <= cpu_instruction_master_read & cpu_instruction_master_run & ~cpu_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_instruction_master_is_granted_some_slave = cpu_instruction_master_granted_custom_dma_burst_1_upstream |
    cpu_instruction_master_granted_custom_dma_burst_3_upstream;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_instruction_master_readdatavalid = cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream |
    cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_instruction_master_readdatavalid = cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid |
    cpu_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_instruction_master_readdatavalid;

  //cpu/instruction_master readdata mux, which is an e_mux
  assign cpu_instruction_master_readdata = ({32 {~cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream}} | custom_dma_burst_1_upstream_readdata_from_sa) &
    ({32 {~cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream}} | custom_dma_burst_3_upstream_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign cpu_instruction_master_waitrequest = ~cpu_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_latency_counter <= 0;
      else 
        cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_instruction_master_latency_counter = ((cpu_instruction_master_run & cpu_instruction_master_read))? latency_load_value :
    (cpu_instruction_master_latency_counter)? cpu_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_address_last_time <= 0;
      else 
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
    end


  //cpu/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_instruction_master_waitrequest & (cpu_instruction_master_read);
    end


  //cpu_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_address != cpu_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_burstcount_last_time <= 0;
      else 
        cpu_instruction_master_burstcount_last_time <= cpu_instruction_master_burstcount;
    end


  //cpu_instruction_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_burstcount != cpu_instruction_master_burstcount_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_instruction_master_read_last_time <= 0;
      else 
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
    end


  //cpu_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_instruction_master_read != cpu_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_custom_dma_burst_0_upstream_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_0_upstream_module (
                                                                            // inputs:
                                                                             clear_fifo,
                                                                             clk,
                                                                             data_in,
                                                                             read,
                                                                             reset_n,
                                                                             sync_reset,
                                                                             write,

                                                                            // outputs:
                                                                             data_out,
                                                                             empty,
                                                                             fifo_contains_ones_n,
                                                                             full
                                                                          )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_0_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_data_master_address_to_slave,
                                                 cpu_data_master_burstcount,
                                                 cpu_data_master_byteenable,
                                                 cpu_data_master_debugaccess,
                                                 cpu_data_master_latency_counter,
                                                 cpu_data_master_read,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register,
                                                 cpu_data_master_write,
                                                 cpu_data_master_writedata,
                                                 custom_dma_burst_0_upstream_readdata,
                                                 custom_dma_burst_0_upstream_readdatavalid,
                                                 custom_dma_burst_0_upstream_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_data_master_granted_custom_dma_burst_0_upstream,
                                                 cpu_data_master_qualified_request_custom_dma_burst_0_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_0_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register,
                                                 cpu_data_master_requests_custom_dma_burst_0_upstream,
                                                 custom_dma_burst_0_upstream_address,
                                                 custom_dma_burst_0_upstream_burstcount,
                                                 custom_dma_burst_0_upstream_byteaddress,
                                                 custom_dma_burst_0_upstream_byteenable,
                                                 custom_dma_burst_0_upstream_debugaccess,
                                                 custom_dma_burst_0_upstream_read,
                                                 custom_dma_burst_0_upstream_readdata_from_sa,
                                                 custom_dma_burst_0_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_0_upstream_write,
                                                 custom_dma_burst_0_upstream_writedata,
                                                 d1_custom_dma_burst_0_upstream_end_xfer
                                              )
;

  output           cpu_data_master_granted_custom_dma_burst_0_upstream;
  output           cpu_data_master_qualified_request_custom_dma_burst_0_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_0_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  output           cpu_data_master_requests_custom_dma_burst_0_upstream;
  output  [ 20: 0] custom_dma_burst_0_upstream_address;
  output  [  3: 0] custom_dma_burst_0_upstream_burstcount;
  output  [ 22: 0] custom_dma_burst_0_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_0_upstream_byteenable;
  output           custom_dma_burst_0_upstream_debugaccess;
  output           custom_dma_burst_0_upstream_read;
  output  [ 31: 0] custom_dma_burst_0_upstream_readdata_from_sa;
  output           custom_dma_burst_0_upstream_waitrequest_from_sa;
  output           custom_dma_burst_0_upstream_write;
  output  [ 31: 0] custom_dma_burst_0_upstream_writedata;
  output           d1_custom_dma_burst_0_upstream_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  input            cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] custom_dma_burst_0_upstream_readdata;
  input            custom_dma_burst_0_upstream_readdatavalid;
  input            custom_dma_burst_0_upstream_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_custom_dma_burst_0_upstream;
  wire             cpu_data_master_qualified_request_custom_dma_burst_0_upstream;
  wire             cpu_data_master_rdv_fifo_empty_custom_dma_burst_0_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_custom_dma_burst_0_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_0_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  wire             cpu_data_master_requests_custom_dma_burst_0_upstream;
  wire             cpu_data_master_saved_grant_custom_dma_burst_0_upstream;
  wire    [ 20: 0] custom_dma_burst_0_upstream_address;
  wire             custom_dma_burst_0_upstream_allgrants;
  wire             custom_dma_burst_0_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_0_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_0_upstream_any_continuerequest;
  wire             custom_dma_burst_0_upstream_arb_counter_enable;
  reg     [  3: 0] custom_dma_burst_0_upstream_arb_share_counter;
  wire    [  3: 0] custom_dma_burst_0_upstream_arb_share_counter_next_value;
  wire    [  3: 0] custom_dma_burst_0_upstream_arb_share_set_values;
  reg     [  2: 0] custom_dma_burst_0_upstream_bbt_burstcounter;
  wire             custom_dma_burst_0_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_0_upstream_begins_xfer;
  wire    [  3: 0] custom_dma_burst_0_upstream_burstcount;
  wire             custom_dma_burst_0_upstream_burstcount_fifo_empty;
  wire    [ 22: 0] custom_dma_burst_0_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_0_upstream_byteenable;
  reg     [  3: 0] custom_dma_burst_0_upstream_current_burst;
  wire    [  3: 0] custom_dma_burst_0_upstream_current_burst_minus_one;
  wire             custom_dma_burst_0_upstream_debugaccess;
  wire             custom_dma_burst_0_upstream_end_xfer;
  wire             custom_dma_burst_0_upstream_firsttransfer;
  wire             custom_dma_burst_0_upstream_grant_vector;
  wire             custom_dma_burst_0_upstream_in_a_read_cycle;
  wire             custom_dma_burst_0_upstream_in_a_write_cycle;
  reg              custom_dma_burst_0_upstream_load_fifo;
  wire             custom_dma_burst_0_upstream_master_qreq_vector;
  wire             custom_dma_burst_0_upstream_move_on_to_next_transaction;
  wire    [  2: 0] custom_dma_burst_0_upstream_next_bbt_burstcount;
  wire    [  3: 0] custom_dma_burst_0_upstream_next_burst_count;
  wire             custom_dma_burst_0_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_0_upstream_read;
  wire    [ 31: 0] custom_dma_burst_0_upstream_readdata_from_sa;
  wire             custom_dma_burst_0_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_0_upstream_reg_firsttransfer;
  wire    [  3: 0] custom_dma_burst_0_upstream_selected_burstcount;
  reg              custom_dma_burst_0_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_0_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_0_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] custom_dma_burst_0_upstream_transaction_burst_count;
  wire             custom_dma_burst_0_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_0_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_0_upstream_waits_for_read;
  wire             custom_dma_burst_0_upstream_waits_for_write;
  wire             custom_dma_burst_0_upstream_write;
  wire    [ 31: 0] custom_dma_burst_0_upstream_writedata;
  reg              d1_custom_dma_burst_0_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_custom_dma_burst_0_upstream_load_fifo;
  wire             wait_for_custom_dma_burst_0_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_0_upstream_end_xfer;
    end


  assign custom_dma_burst_0_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_custom_dma_burst_0_upstream));
  //assign custom_dma_burst_0_upstream_readdata_from_sa = custom_dma_burst_0_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_0_upstream_readdata_from_sa = custom_dma_burst_0_upstream_readdata;

  assign cpu_data_master_requests_custom_dma_burst_0_upstream = ({cpu_data_master_address_to_slave[26 : 21] , 21'b0} == 27'h6000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign custom_dma_burst_0_upstream_waitrequest_from_sa = custom_dma_burst_0_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_0_upstream_waitrequest_from_sa = custom_dma_burst_0_upstream_waitrequest;

  //assign custom_dma_burst_0_upstream_readdatavalid_from_sa = custom_dma_burst_0_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_0_upstream_readdatavalid_from_sa = custom_dma_burst_0_upstream_readdatavalid;

  //custom_dma_burst_0_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_0_upstream_arb_share_set_values = (cpu_data_master_granted_custom_dma_burst_0_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //custom_dma_burst_0_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_0_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_0_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_0_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_custom_dma_burst_0_upstream;

  //custom_dma_burst_0_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_0_upstream_arb_share_counter_next_value = custom_dma_burst_0_upstream_firsttransfer ? (custom_dma_burst_0_upstream_arb_share_set_values - 1) : |custom_dma_burst_0_upstream_arb_share_counter ? (custom_dma_burst_0_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_0_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_0_upstream_allgrants = |custom_dma_burst_0_upstream_grant_vector;

  //custom_dma_burst_0_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_0_upstream_end_xfer = ~(custom_dma_burst_0_upstream_waits_for_read | custom_dma_burst_0_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream = custom_dma_burst_0_upstream_end_xfer & (~custom_dma_burst_0_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_0_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_0_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream & custom_dma_burst_0_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream & ~custom_dma_burst_0_upstream_non_bursting_master_requests);

  //custom_dma_burst_0_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_0_upstream_arb_counter_enable)
          custom_dma_burst_0_upstream_arb_share_counter <= custom_dma_burst_0_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_0_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_0_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_0_upstream & ~custom_dma_burst_0_upstream_non_bursting_master_requests))
          custom_dma_burst_0_upstream_slavearbiterlockenable <= |custom_dma_burst_0_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master custom_dma_burst_0/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = custom_dma_burst_0_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //custom_dma_burst_0_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_0_upstream_slavearbiterlockenable2 = |custom_dma_burst_0_upstream_arb_share_counter_next_value;

  //cpu/data_master custom_dma_burst_0/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = custom_dma_burst_0_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //custom_dma_burst_0_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_0_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_custom_dma_burst_0_upstream = cpu_data_master_requests_custom_dma_burst_0_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register) | (|cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register))));
  //unique name for custom_dma_burst_0_upstream_move_on_to_next_transaction, which is an e_assign
  assign custom_dma_burst_0_upstream_move_on_to_next_transaction = custom_dma_burst_0_upstream_this_cycle_is_the_last_burst & custom_dma_burst_0_upstream_load_fifo;

  //the currently selected burstcount for custom_dma_burst_0_upstream, which is an e_mux
  assign custom_dma_burst_0_upstream_selected_burstcount = (cpu_data_master_granted_custom_dma_burst_0_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_custom_dma_burst_0_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_custom_dma_burst_0_upstream_module burstcount_fifo_for_custom_dma_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_0_upstream_selected_burstcount),
      .data_out             (custom_dma_burst_0_upstream_transaction_burst_count),
      .empty                (custom_dma_burst_0_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (custom_dma_burst_0_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read & custom_dma_burst_0_upstream_load_fifo & ~(custom_dma_burst_0_upstream_this_cycle_is_the_last_burst & custom_dma_burst_0_upstream_burstcount_fifo_empty))
    );

  //custom_dma_burst_0_upstream current burst minus one, which is an e_assign
  assign custom_dma_burst_0_upstream_current_burst_minus_one = custom_dma_burst_0_upstream_current_burst - 1;

  //what to load in current_burst, for custom_dma_burst_0_upstream, which is an e_mux
  assign custom_dma_burst_0_upstream_next_burst_count = (((in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read) & ~custom_dma_burst_0_upstream_load_fifo))? custom_dma_burst_0_upstream_selected_burstcount :
    ((in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read & custom_dma_burst_0_upstream_this_cycle_is_the_last_burst & custom_dma_burst_0_upstream_burstcount_fifo_empty))? custom_dma_burst_0_upstream_selected_burstcount :
    (custom_dma_burst_0_upstream_this_cycle_is_the_last_burst)? custom_dma_burst_0_upstream_transaction_burst_count :
    custom_dma_burst_0_upstream_current_burst_minus_one;

  //the current burst count for custom_dma_burst_0_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_current_burst <= 0;
      else if (custom_dma_burst_0_upstream_readdatavalid_from_sa | (~custom_dma_burst_0_upstream_load_fifo & (in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read)))
          custom_dma_burst_0_upstream_current_burst <= custom_dma_burst_0_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_custom_dma_burst_0_upstream_load_fifo = (~custom_dma_burst_0_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read) & custom_dma_burst_0_upstream_load_fifo))? 1 :
    ~custom_dma_burst_0_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read) & ~custom_dma_burst_0_upstream_load_fifo | custom_dma_burst_0_upstream_this_cycle_is_the_last_burst)
          custom_dma_burst_0_upstream_load_fifo <= p0_custom_dma_burst_0_upstream_load_fifo;
    end


  //the last cycle in the burst for custom_dma_burst_0_upstream, which is an e_assign
  assign custom_dma_burst_0_upstream_this_cycle_is_the_last_burst = ~(|custom_dma_burst_0_upstream_current_burst_minus_one) & custom_dma_burst_0_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_custom_dma_burst_0_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_custom_dma_burst_0_upstream_module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_0_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_custom_dma_burst_0_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_custom_dma_burst_0_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_custom_dma_burst_0_upstream),
      .full                 (),
      .read                 (custom_dma_burst_0_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_0_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_custom_dma_burst_0_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_custom_dma_burst_0_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_custom_dma_burst_0_upstream = custom_dma_burst_0_upstream_readdatavalid_from_sa;

  //custom_dma_burst_0_upstream_writedata mux, which is an e_mux
  assign custom_dma_burst_0_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for custom_dma_burst_0/upstream, which is an e_mux
  assign custom_dma_burst_0_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_custom_dma_burst_0_upstream = cpu_data_master_qualified_request_custom_dma_burst_0_upstream;

  //cpu/data_master saved-grant custom_dma_burst_0/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_custom_dma_burst_0_upstream = cpu_data_master_requests_custom_dma_burst_0_upstream;

  //allow new arb cycle for custom_dma_burst_0/upstream, which is an e_assign
  assign custom_dma_burst_0_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_0_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_0_upstream_master_qreq_vector = 1;

  //custom_dma_burst_0_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_0_upstream_firsttransfer = custom_dma_burst_0_upstream_begins_xfer ? custom_dma_burst_0_upstream_unreg_firsttransfer : custom_dma_burst_0_upstream_reg_firsttransfer;

  //custom_dma_burst_0_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_0_upstream_unreg_firsttransfer = ~(custom_dma_burst_0_upstream_slavearbiterlockenable & custom_dma_burst_0_upstream_any_continuerequest);

  //custom_dma_burst_0_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_0_upstream_begins_xfer)
          custom_dma_burst_0_upstream_reg_firsttransfer <= custom_dma_burst_0_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_0_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign custom_dma_burst_0_upstream_next_bbt_burstcount = ((((custom_dma_burst_0_upstream_write) && (custom_dma_burst_0_upstream_bbt_burstcounter == 0))))? (custom_dma_burst_0_upstream_burstcount - 1) :
    ((((custom_dma_burst_0_upstream_read) && (custom_dma_burst_0_upstream_bbt_burstcounter == 0))))? 0 :
    (custom_dma_burst_0_upstream_bbt_burstcounter - 1);

  //custom_dma_burst_0_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_upstream_bbt_burstcounter <= 0;
      else if (custom_dma_burst_0_upstream_begins_xfer)
          custom_dma_burst_0_upstream_bbt_burstcounter <= custom_dma_burst_0_upstream_next_bbt_burstcount;
    end


  //custom_dma_burst_0_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_0_upstream_beginbursttransfer_internal = custom_dma_burst_0_upstream_begins_xfer & (custom_dma_burst_0_upstream_bbt_burstcounter == 0);

  //custom_dma_burst_0_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_0_upstream_read = cpu_data_master_granted_custom_dma_burst_0_upstream & cpu_data_master_read;

  //custom_dma_burst_0_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_0_upstream_write = cpu_data_master_granted_custom_dma_burst_0_upstream & cpu_data_master_write;

  //custom_dma_burst_0_upstream_address mux, which is an e_mux
  assign custom_dma_burst_0_upstream_address = cpu_data_master_address_to_slave;

  //d1_custom_dma_burst_0_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_0_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_0_upstream_end_xfer <= custom_dma_burst_0_upstream_end_xfer;
    end


  //custom_dma_burst_0_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_0_upstream_waits_for_read = custom_dma_burst_0_upstream_in_a_read_cycle & custom_dma_burst_0_upstream_waitrequest_from_sa;

  //custom_dma_burst_0_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_0_upstream_in_a_read_cycle = cpu_data_master_granted_custom_dma_burst_0_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_0_upstream_in_a_read_cycle;

  //custom_dma_burst_0_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_0_upstream_waits_for_write = custom_dma_burst_0_upstream_in_a_write_cycle & custom_dma_burst_0_upstream_waitrequest_from_sa;

  //custom_dma_burst_0_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_0_upstream_in_a_write_cycle = cpu_data_master_granted_custom_dma_burst_0_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_0_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_0_upstream_counter = 0;
  //custom_dma_burst_0_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_0_upstream_byteenable = (cpu_data_master_granted_custom_dma_burst_0_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign custom_dma_burst_0_upstream_burstcount = (cpu_data_master_granted_custom_dma_burst_0_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_0_upstream_debugaccess = (cpu_data_master_granted_custom_dma_burst_0_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_0/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_custom_dma_burst_0_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_0/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_0_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_0_downstream_address,
                                                   custom_dma_burst_0_downstream_burstcount,
                                                   custom_dma_burst_0_downstream_byteenable,
                                                   custom_dma_burst_0_downstream_granted_ext_ssram_s1,
                                                   custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1,
                                                   custom_dma_burst_0_downstream_read,
                                                   custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1,
                                                   custom_dma_burst_0_downstream_requests_ext_ssram_s1,
                                                   custom_dma_burst_0_downstream_write,
                                                   custom_dma_burst_0_downstream_writedata,
                                                   d1_ext_ssram_bus_avalon_slave_end_xfer,
                                                   incoming_ext_ssram_bus_data,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_0_downstream_address_to_slave,
                                                   custom_dma_burst_0_downstream_latency_counter,
                                                   custom_dma_burst_0_downstream_readdata,
                                                   custom_dma_burst_0_downstream_readdatavalid,
                                                   custom_dma_burst_0_downstream_reset_n,
                                                   custom_dma_burst_0_downstream_waitrequest
                                                )
;

  output  [ 20: 0] custom_dma_burst_0_downstream_address_to_slave;
  output  [  2: 0] custom_dma_burst_0_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_0_downstream_readdata;
  output           custom_dma_burst_0_downstream_readdatavalid;
  output           custom_dma_burst_0_downstream_reset_n;
  output           custom_dma_burst_0_downstream_waitrequest;
  input            clk;
  input   [ 20: 0] custom_dma_burst_0_downstream_address;
  input            custom_dma_burst_0_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_0_downstream_byteenable;
  input            custom_dma_burst_0_downstream_granted_ext_ssram_s1;
  input            custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1;
  input            custom_dma_burst_0_downstream_read;
  input            custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1;
  input            custom_dma_burst_0_downstream_requests_ext_ssram_s1;
  input            custom_dma_burst_0_downstream_write;
  input   [ 31: 0] custom_dma_burst_0_downstream_writedata;
  input            d1_ext_ssram_bus_avalon_slave_end_xfer;
  input   [ 31: 0] incoming_ext_ssram_bus_data;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 20: 0] custom_dma_burst_0_downstream_address_last_time;
  wire    [ 20: 0] custom_dma_burst_0_downstream_address_to_slave;
  reg              custom_dma_burst_0_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_0_downstream_byteenable_last_time;
  wire             custom_dma_burst_0_downstream_is_granted_some_slave;
  reg     [  2: 0] custom_dma_burst_0_downstream_latency_counter;
  reg              custom_dma_burst_0_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_0_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_0_downstream_readdata;
  wire             custom_dma_burst_0_downstream_readdatavalid;
  wire             custom_dma_burst_0_downstream_reset_n;
  wire             custom_dma_burst_0_downstream_run;
  wire             custom_dma_burst_0_downstream_waitrequest;
  reg              custom_dma_burst_0_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_0_downstream_writedata_last_time;
  wire    [  2: 0] latency_load_value;
  wire    [  2: 0] p1_custom_dma_burst_0_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_0_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 | ~custom_dma_burst_0_downstream_requests_ext_ssram_s1) & (custom_dma_burst_0_downstream_granted_ext_ssram_s1 | ~custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1) & ((~custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 | ~(custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write) | (1 & (custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write)))) & ((~custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 | ~(custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write) | (1 & (custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_0_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_0_downstream_address_to_slave = custom_dma_burst_0_downstream_address;

  //custom_dma_burst_0_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_0_downstream_read_but_no_slave_selected <= custom_dma_burst_0_downstream_read & custom_dma_burst_0_downstream_run & ~custom_dma_burst_0_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_0_downstream_is_granted_some_slave = custom_dma_burst_0_downstream_granted_ext_ssram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_0_downstream_readdatavalid = custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_0_downstream_readdatavalid = custom_dma_burst_0_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_0_downstream_readdatavalid;

  //custom_dma_burst_0/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_0_downstream_readdata = incoming_ext_ssram_bus_data;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_0_downstream_waitrequest = ~custom_dma_burst_0_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_0_downstream_latency_counter <= p1_custom_dma_burst_0_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_0_downstream_latency_counter = ((custom_dma_burst_0_downstream_run & custom_dma_burst_0_downstream_read))? latency_load_value :
    (custom_dma_burst_0_downstream_latency_counter)? custom_dma_burst_0_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {3 {custom_dma_burst_0_downstream_requests_ext_ssram_s1}} & 4;

  //custom_dma_burst_0_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_0_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_0_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_address_last_time <= custom_dma_burst_0_downstream_address;
    end


  //custom_dma_burst_0/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_0_downstream_waitrequest & (custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write);
    end


  //custom_dma_burst_0_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_address != custom_dma_burst_0_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_0_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_burstcount_last_time <= custom_dma_burst_0_downstream_burstcount;
    end


  //custom_dma_burst_0_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_burstcount != custom_dma_burst_0_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_0_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_byteenable_last_time <= custom_dma_burst_0_downstream_byteenable;
    end


  //custom_dma_burst_0_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_byteenable != custom_dma_burst_0_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_0_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_read_last_time <= custom_dma_burst_0_downstream_read;
    end


  //custom_dma_burst_0_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_read != custom_dma_burst_0_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_0_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_write_last_time <= custom_dma_burst_0_downstream_write;
    end


  //custom_dma_burst_0_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_write != custom_dma_burst_0_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_0_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_0_downstream_writedata_last_time <= custom_dma_burst_0_downstream_writedata;
    end


  //custom_dma_burst_0_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_0_downstream_writedata != custom_dma_burst_0_downstream_writedata_last_time) & custom_dma_burst_0_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_0_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_custom_dma_burst_1_upstream_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_1_upstream_module (
                                                                                   // inputs:
                                                                                    clear_fifo,
                                                                                    clk,
                                                                                    data_in,
                                                                                    read,
                                                                                    reset_n,
                                                                                    sync_reset,
                                                                                    write,

                                                                                   // outputs:
                                                                                    data_out,
                                                                                    empty,
                                                                                    fifo_contains_ones_n,
                                                                                    full
                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_1_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_instruction_master_address_to_slave,
                                                 cpu_instruction_master_burstcount,
                                                 cpu_instruction_master_latency_counter,
                                                 cpu_instruction_master_read,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register,
                                                 custom_dma_burst_1_upstream_readdata,
                                                 custom_dma_burst_1_upstream_readdatavalid,
                                                 custom_dma_burst_1_upstream_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_instruction_master_granted_custom_dma_burst_1_upstream,
                                                 cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register,
                                                 cpu_instruction_master_requests_custom_dma_burst_1_upstream,
                                                 custom_dma_burst_1_upstream_address,
                                                 custom_dma_burst_1_upstream_byteaddress,
                                                 custom_dma_burst_1_upstream_byteenable,
                                                 custom_dma_burst_1_upstream_debugaccess,
                                                 custom_dma_burst_1_upstream_read,
                                                 custom_dma_burst_1_upstream_readdata_from_sa,
                                                 custom_dma_burst_1_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_1_upstream_write,
                                                 d1_custom_dma_burst_1_upstream_end_xfer
                                              )
;

  output           cpu_instruction_master_granted_custom_dma_burst_1_upstream;
  output           cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream;
  output           cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream;
  output           cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register;
  output           cpu_instruction_master_requests_custom_dma_burst_1_upstream;
  output  [ 11: 0] custom_dma_burst_1_upstream_address;
  output  [ 13: 0] custom_dma_burst_1_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_1_upstream_byteenable;
  output           custom_dma_burst_1_upstream_debugaccess;
  output           custom_dma_burst_1_upstream_read;
  output  [ 31: 0] custom_dma_burst_1_upstream_readdata_from_sa;
  output           custom_dma_burst_1_upstream_waitrequest_from_sa;
  output           custom_dma_burst_1_upstream_write;
  output           d1_custom_dma_burst_1_upstream_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register;
  input   [ 31: 0] custom_dma_burst_1_upstream_readdata;
  input            custom_dma_burst_1_upstream_readdatavalid;
  input            custom_dma_burst_1_upstream_waitrequest;
  input            reset_n;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register;
  wire             cpu_instruction_master_requests_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_saved_grant_custom_dma_burst_1_upstream;
  wire    [ 11: 0] custom_dma_burst_1_upstream_address;
  wire             custom_dma_burst_1_upstream_allgrants;
  wire             custom_dma_burst_1_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_1_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_1_upstream_any_continuerequest;
  wire             custom_dma_burst_1_upstream_arb_counter_enable;
  reg     [  3: 0] custom_dma_burst_1_upstream_arb_share_counter;
  wire    [  3: 0] custom_dma_burst_1_upstream_arb_share_counter_next_value;
  wire    [  3: 0] custom_dma_burst_1_upstream_arb_share_set_values;
  wire             custom_dma_burst_1_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_1_upstream_begins_xfer;
  wire             custom_dma_burst_1_upstream_burstcount_fifo_empty;
  wire    [ 13: 0] custom_dma_burst_1_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_1_upstream_byteenable;
  reg     [  3: 0] custom_dma_burst_1_upstream_current_burst;
  wire    [  3: 0] custom_dma_burst_1_upstream_current_burst_minus_one;
  wire             custom_dma_burst_1_upstream_debugaccess;
  wire             custom_dma_burst_1_upstream_end_xfer;
  wire             custom_dma_burst_1_upstream_firsttransfer;
  wire             custom_dma_burst_1_upstream_grant_vector;
  wire             custom_dma_burst_1_upstream_in_a_read_cycle;
  wire             custom_dma_burst_1_upstream_in_a_write_cycle;
  reg              custom_dma_burst_1_upstream_load_fifo;
  wire             custom_dma_burst_1_upstream_master_qreq_vector;
  wire             custom_dma_burst_1_upstream_move_on_to_next_transaction;
  wire    [  3: 0] custom_dma_burst_1_upstream_next_burst_count;
  wire             custom_dma_burst_1_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_1_upstream_read;
  wire    [ 31: 0] custom_dma_burst_1_upstream_readdata_from_sa;
  wire             custom_dma_burst_1_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_1_upstream_reg_firsttransfer;
  wire    [  3: 0] custom_dma_burst_1_upstream_selected_burstcount;
  reg              custom_dma_burst_1_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_1_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_1_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] custom_dma_burst_1_upstream_transaction_burst_count;
  wire             custom_dma_burst_1_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_1_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_1_upstream_waits_for_read;
  wire             custom_dma_burst_1_upstream_waits_for_write;
  wire             custom_dma_burst_1_upstream_write;
  reg              d1_custom_dma_burst_1_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_custom_dma_burst_1_upstream_load_fifo;
  wire             wait_for_custom_dma_burst_1_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_1_upstream_end_xfer;
    end


  assign custom_dma_burst_1_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream));
  //assign custom_dma_burst_1_upstream_readdata_from_sa = custom_dma_burst_1_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_1_upstream_readdata_from_sa = custom_dma_burst_1_upstream_readdata;

  assign cpu_instruction_master_requests_custom_dma_burst_1_upstream = (({cpu_instruction_master_address_to_slave[26 : 12] , 12'b0} == 27'h5000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign custom_dma_burst_1_upstream_waitrequest_from_sa = custom_dma_burst_1_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_1_upstream_waitrequest_from_sa = custom_dma_burst_1_upstream_waitrequest;

  //assign custom_dma_burst_1_upstream_readdatavalid_from_sa = custom_dma_burst_1_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_1_upstream_readdatavalid_from_sa = custom_dma_burst_1_upstream_readdatavalid;

  //custom_dma_burst_1_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_1_upstream_arb_share_set_values = 1;

  //custom_dma_burst_1_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_1_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_1_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_1_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_custom_dma_burst_1_upstream;

  //custom_dma_burst_1_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_1_upstream_arb_share_counter_next_value = custom_dma_burst_1_upstream_firsttransfer ? (custom_dma_burst_1_upstream_arb_share_set_values - 1) : |custom_dma_burst_1_upstream_arb_share_counter ? (custom_dma_burst_1_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_1_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_1_upstream_allgrants = |custom_dma_burst_1_upstream_grant_vector;

  //custom_dma_burst_1_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_1_upstream_end_xfer = ~(custom_dma_burst_1_upstream_waits_for_read | custom_dma_burst_1_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream = custom_dma_burst_1_upstream_end_xfer & (~custom_dma_burst_1_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_1_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_1_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream & custom_dma_burst_1_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream & ~custom_dma_burst_1_upstream_non_bursting_master_requests);

  //custom_dma_burst_1_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_1_upstream_arb_counter_enable)
          custom_dma_burst_1_upstream_arb_share_counter <= custom_dma_burst_1_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_1_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_1_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_1_upstream & ~custom_dma_burst_1_upstream_non_bursting_master_requests))
          custom_dma_burst_1_upstream_slavearbiterlockenable <= |custom_dma_burst_1_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master custom_dma_burst_1/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = custom_dma_burst_1_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //custom_dma_burst_1_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_1_upstream_slavearbiterlockenable2 = |custom_dma_burst_1_upstream_arb_share_counter_next_value;

  //cpu/instruction_master custom_dma_burst_1/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = custom_dma_burst_1_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //custom_dma_burst_1_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_1_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream = cpu_instruction_master_requests_custom_dma_burst_1_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register))));
  //unique name for custom_dma_burst_1_upstream_move_on_to_next_transaction, which is an e_assign
  assign custom_dma_burst_1_upstream_move_on_to_next_transaction = custom_dma_burst_1_upstream_this_cycle_is_the_last_burst & custom_dma_burst_1_upstream_load_fifo;

  //the currently selected burstcount for custom_dma_burst_1_upstream, which is an e_mux
  assign custom_dma_burst_1_upstream_selected_burstcount = (cpu_instruction_master_granted_custom_dma_burst_1_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_custom_dma_burst_1_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_custom_dma_burst_1_upstream_module burstcount_fifo_for_custom_dma_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_1_upstream_selected_burstcount),
      .data_out             (custom_dma_burst_1_upstream_transaction_burst_count),
      .empty                (custom_dma_burst_1_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (custom_dma_burst_1_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read & custom_dma_burst_1_upstream_load_fifo & ~(custom_dma_burst_1_upstream_this_cycle_is_the_last_burst & custom_dma_burst_1_upstream_burstcount_fifo_empty))
    );

  //custom_dma_burst_1_upstream current burst minus one, which is an e_assign
  assign custom_dma_burst_1_upstream_current_burst_minus_one = custom_dma_burst_1_upstream_current_burst - 1;

  //what to load in current_burst, for custom_dma_burst_1_upstream, which is an e_mux
  assign custom_dma_burst_1_upstream_next_burst_count = (((in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read) & ~custom_dma_burst_1_upstream_load_fifo))? custom_dma_burst_1_upstream_selected_burstcount :
    ((in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read & custom_dma_burst_1_upstream_this_cycle_is_the_last_burst & custom_dma_burst_1_upstream_burstcount_fifo_empty))? custom_dma_burst_1_upstream_selected_burstcount :
    (custom_dma_burst_1_upstream_this_cycle_is_the_last_burst)? custom_dma_burst_1_upstream_transaction_burst_count :
    custom_dma_burst_1_upstream_current_burst_minus_one;

  //the current burst count for custom_dma_burst_1_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_upstream_current_burst <= 0;
      else if (custom_dma_burst_1_upstream_readdatavalid_from_sa | (~custom_dma_burst_1_upstream_load_fifo & (in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read)))
          custom_dma_burst_1_upstream_current_burst <= custom_dma_burst_1_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_custom_dma_burst_1_upstream_load_fifo = (~custom_dma_burst_1_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read) & custom_dma_burst_1_upstream_load_fifo))? 1 :
    ~custom_dma_burst_1_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read) & ~custom_dma_burst_1_upstream_load_fifo | custom_dma_burst_1_upstream_this_cycle_is_the_last_burst)
          custom_dma_burst_1_upstream_load_fifo <= p0_custom_dma_burst_1_upstream_load_fifo;
    end


  //the last cycle in the burst for custom_dma_burst_1_upstream, which is an e_assign
  assign custom_dma_burst_1_upstream_this_cycle_is_the_last_burst = ~(|custom_dma_burst_1_upstream_current_burst_minus_one) & custom_dma_burst_1_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_1_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_1_upstream_module rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_1_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_custom_dma_burst_1_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_custom_dma_burst_1_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_1_upstream),
      .full                 (),
      .read                 (custom_dma_burst_1_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_1_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_1_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream = custom_dma_burst_1_upstream_readdatavalid_from_sa;

  //byteaddress mux for custom_dma_burst_1/upstream, which is an e_mux
  assign custom_dma_burst_1_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_custom_dma_burst_1_upstream = cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream;

  //cpu/instruction_master saved-grant custom_dma_burst_1/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_custom_dma_burst_1_upstream = cpu_instruction_master_requests_custom_dma_burst_1_upstream;

  //allow new arb cycle for custom_dma_burst_1/upstream, which is an e_assign
  assign custom_dma_burst_1_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_1_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_1_upstream_master_qreq_vector = 1;

  //custom_dma_burst_1_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_1_upstream_firsttransfer = custom_dma_burst_1_upstream_begins_xfer ? custom_dma_burst_1_upstream_unreg_firsttransfer : custom_dma_burst_1_upstream_reg_firsttransfer;

  //custom_dma_burst_1_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_1_upstream_unreg_firsttransfer = ~(custom_dma_burst_1_upstream_slavearbiterlockenable & custom_dma_burst_1_upstream_any_continuerequest);

  //custom_dma_burst_1_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_1_upstream_begins_xfer)
          custom_dma_burst_1_upstream_reg_firsttransfer <= custom_dma_burst_1_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_1_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_1_upstream_beginbursttransfer_internal = custom_dma_burst_1_upstream_begins_xfer;

  //custom_dma_burst_1_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_1_upstream_read = cpu_instruction_master_granted_custom_dma_burst_1_upstream & cpu_instruction_master_read;

  //custom_dma_burst_1_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_1_upstream_write = 0;

  //custom_dma_burst_1_upstream_address mux, which is an e_mux
  assign custom_dma_burst_1_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_custom_dma_burst_1_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_1_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_1_upstream_end_xfer <= custom_dma_burst_1_upstream_end_xfer;
    end


  //custom_dma_burst_1_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_1_upstream_waits_for_read = custom_dma_burst_1_upstream_in_a_read_cycle & custom_dma_burst_1_upstream_waitrequest_from_sa;

  //custom_dma_burst_1_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_1_upstream_in_a_read_cycle = cpu_instruction_master_granted_custom_dma_burst_1_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_1_upstream_in_a_read_cycle;

  //custom_dma_burst_1_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_1_upstream_waits_for_write = custom_dma_burst_1_upstream_in_a_write_cycle & custom_dma_burst_1_upstream_waitrequest_from_sa;

  //custom_dma_burst_1_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_1_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_1_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_1_upstream_counter = 0;
  //custom_dma_burst_1_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_1_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_1_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_1/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_custom_dma_burst_1_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_1/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_1_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_1_downstream_address,
                                                   custom_dma_burst_1_downstream_burstcount,
                                                   custom_dma_burst_1_downstream_byteenable,
                                                   custom_dma_burst_1_downstream_granted_pipeline_bridge_s1,
                                                   custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1,
                                                   custom_dma_burst_1_downstream_read,
                                                   custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1,
                                                   custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register,
                                                   custom_dma_burst_1_downstream_requests_pipeline_bridge_s1,
                                                   custom_dma_burst_1_downstream_write,
                                                   custom_dma_burst_1_downstream_writedata,
                                                   d1_pipeline_bridge_s1_end_xfer,
                                                   pipeline_bridge_s1_readdata_from_sa,
                                                   pipeline_bridge_s1_waitrequest_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_1_downstream_address_to_slave,
                                                   custom_dma_burst_1_downstream_latency_counter,
                                                   custom_dma_burst_1_downstream_readdata,
                                                   custom_dma_burst_1_downstream_readdatavalid,
                                                   custom_dma_burst_1_downstream_reset_n,
                                                   custom_dma_burst_1_downstream_waitrequest
                                                )
;

  output  [ 11: 0] custom_dma_burst_1_downstream_address_to_slave;
  output           custom_dma_burst_1_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_1_downstream_readdata;
  output           custom_dma_burst_1_downstream_readdatavalid;
  output           custom_dma_burst_1_downstream_reset_n;
  output           custom_dma_burst_1_downstream_waitrequest;
  input            clk;
  input   [ 11: 0] custom_dma_burst_1_downstream_address;
  input            custom_dma_burst_1_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_1_downstream_byteenable;
  input            custom_dma_burst_1_downstream_granted_pipeline_bridge_s1;
  input            custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1;
  input            custom_dma_burst_1_downstream_read;
  input            custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1;
  input            custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  input            custom_dma_burst_1_downstream_requests_pipeline_bridge_s1;
  input            custom_dma_burst_1_downstream_write;
  input   [ 31: 0] custom_dma_burst_1_downstream_writedata;
  input            d1_pipeline_bridge_s1_end_xfer;
  input   [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 11: 0] custom_dma_burst_1_downstream_address_last_time;
  wire    [ 11: 0] custom_dma_burst_1_downstream_address_to_slave;
  reg              custom_dma_burst_1_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_1_downstream_byteenable_last_time;
  wire             custom_dma_burst_1_downstream_is_granted_some_slave;
  reg              custom_dma_burst_1_downstream_latency_counter;
  reg              custom_dma_burst_1_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_1_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_1_downstream_readdata;
  wire             custom_dma_burst_1_downstream_readdatavalid;
  wire             custom_dma_burst_1_downstream_reset_n;
  wire             custom_dma_burst_1_downstream_run;
  wire             custom_dma_burst_1_downstream_waitrequest;
  reg              custom_dma_burst_1_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_1_downstream_writedata_last_time;
  wire             latency_load_value;
  wire             p1_custom_dma_burst_1_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_1_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1 | ~custom_dma_burst_1_downstream_requests_pipeline_bridge_s1) & (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 | ~custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1) & ((~custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1 | ~(custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write)))) & ((~custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1 | ~(custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_1_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_1_downstream_address_to_slave = custom_dma_burst_1_downstream_address;

  //custom_dma_burst_1_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_1_downstream_read_but_no_slave_selected <= custom_dma_burst_1_downstream_read & custom_dma_burst_1_downstream_run & ~custom_dma_burst_1_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_1_downstream_is_granted_some_slave = custom_dma_burst_1_downstream_granted_pipeline_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_1_downstream_readdatavalid = custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_1_downstream_readdatavalid = custom_dma_burst_1_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_1_downstream_readdatavalid;

  //custom_dma_burst_1/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_1_downstream_readdata = pipeline_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_1_downstream_waitrequest = ~custom_dma_burst_1_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_1_downstream_latency_counter <= p1_custom_dma_burst_1_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_1_downstream_latency_counter = ((custom_dma_burst_1_downstream_run & custom_dma_burst_1_downstream_read))? latency_load_value :
    (custom_dma_burst_1_downstream_latency_counter)? custom_dma_burst_1_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //custom_dma_burst_1_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_1_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_1_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_address_last_time <= custom_dma_burst_1_downstream_address;
    end


  //custom_dma_burst_1/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_1_downstream_waitrequest & (custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write);
    end


  //custom_dma_burst_1_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_address != custom_dma_burst_1_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_1_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_burstcount_last_time <= custom_dma_burst_1_downstream_burstcount;
    end


  //custom_dma_burst_1_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_burstcount != custom_dma_burst_1_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_1_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_byteenable_last_time <= custom_dma_burst_1_downstream_byteenable;
    end


  //custom_dma_burst_1_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_byteenable != custom_dma_burst_1_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_1_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_read_last_time <= custom_dma_burst_1_downstream_read;
    end


  //custom_dma_burst_1_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_read != custom_dma_burst_1_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_1_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_write_last_time <= custom_dma_burst_1_downstream_write;
    end


  //custom_dma_burst_1_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_write != custom_dma_burst_1_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_1_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_1_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_1_downstream_writedata_last_time <= custom_dma_burst_1_downstream_writedata;
    end


  //custom_dma_burst_1_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_1_downstream_writedata != custom_dma_burst_1_downstream_writedata_last_time) & custom_dma_burst_1_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_1_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_custom_dma_burst_2_upstream_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_2_upstream_module (
                                                                            // inputs:
                                                                             clear_fifo,
                                                                             clk,
                                                                             data_in,
                                                                             read,
                                                                             reset_n,
                                                                             sync_reset,
                                                                             write,

                                                                            // outputs:
                                                                             data_out,
                                                                             empty,
                                                                             fifo_contains_ones_n,
                                                                             full
                                                                          )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  wire             full_6;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_5;
  assign empty = !full_0;
  assign full_6 = 0;
  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    0;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_2_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_data_master_address_to_slave,
                                                 cpu_data_master_burstcount,
                                                 cpu_data_master_byteenable,
                                                 cpu_data_master_debugaccess,
                                                 cpu_data_master_latency_counter,
                                                 cpu_data_master_read,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register,
                                                 cpu_data_master_write,
                                                 cpu_data_master_writedata,
                                                 custom_dma_burst_2_upstream_readdata,
                                                 custom_dma_burst_2_upstream_readdatavalid,
                                                 custom_dma_burst_2_upstream_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_data_master_granted_custom_dma_burst_2_upstream,
                                                 cpu_data_master_qualified_request_custom_dma_burst_2_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_2_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register,
                                                 cpu_data_master_requests_custom_dma_burst_2_upstream,
                                                 custom_dma_burst_2_upstream_address,
                                                 custom_dma_burst_2_upstream_burstcount,
                                                 custom_dma_burst_2_upstream_byteaddress,
                                                 custom_dma_burst_2_upstream_byteenable,
                                                 custom_dma_burst_2_upstream_debugaccess,
                                                 custom_dma_burst_2_upstream_read,
                                                 custom_dma_burst_2_upstream_readdata_from_sa,
                                                 custom_dma_burst_2_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_2_upstream_write,
                                                 custom_dma_burst_2_upstream_writedata,
                                                 d1_custom_dma_burst_2_upstream_end_xfer
                                              )
;

  output           cpu_data_master_granted_custom_dma_burst_2_upstream;
  output           cpu_data_master_qualified_request_custom_dma_burst_2_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_2_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  output           cpu_data_master_requests_custom_dma_burst_2_upstream;
  output  [ 11: 0] custom_dma_burst_2_upstream_address;
  output  [  3: 0] custom_dma_burst_2_upstream_burstcount;
  output  [ 13: 0] custom_dma_burst_2_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_2_upstream_byteenable;
  output           custom_dma_burst_2_upstream_debugaccess;
  output           custom_dma_burst_2_upstream_read;
  output  [ 31: 0] custom_dma_burst_2_upstream_readdata_from_sa;
  output           custom_dma_burst_2_upstream_waitrequest_from_sa;
  output           custom_dma_burst_2_upstream_write;
  output  [ 31: 0] custom_dma_burst_2_upstream_writedata;
  output           d1_custom_dma_burst_2_upstream_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  input            cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] custom_dma_burst_2_upstream_readdata;
  input            custom_dma_burst_2_upstream_readdatavalid;
  input            custom_dma_burst_2_upstream_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_custom_dma_burst_2_upstream;
  wire             cpu_data_master_qualified_request_custom_dma_burst_2_upstream;
  wire             cpu_data_master_rdv_fifo_empty_custom_dma_burst_2_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_custom_dma_burst_2_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_2_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  wire             cpu_data_master_requests_custom_dma_burst_2_upstream;
  wire             cpu_data_master_saved_grant_custom_dma_burst_2_upstream;
  wire    [ 11: 0] custom_dma_burst_2_upstream_address;
  wire             custom_dma_burst_2_upstream_allgrants;
  wire             custom_dma_burst_2_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_2_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_2_upstream_any_continuerequest;
  wire             custom_dma_burst_2_upstream_arb_counter_enable;
  reg     [  3: 0] custom_dma_burst_2_upstream_arb_share_counter;
  wire    [  3: 0] custom_dma_burst_2_upstream_arb_share_counter_next_value;
  wire    [  3: 0] custom_dma_burst_2_upstream_arb_share_set_values;
  reg     [  2: 0] custom_dma_burst_2_upstream_bbt_burstcounter;
  wire             custom_dma_burst_2_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_2_upstream_begins_xfer;
  wire    [  3: 0] custom_dma_burst_2_upstream_burstcount;
  wire             custom_dma_burst_2_upstream_burstcount_fifo_empty;
  wire    [ 13: 0] custom_dma_burst_2_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_2_upstream_byteenable;
  reg     [  3: 0] custom_dma_burst_2_upstream_current_burst;
  wire    [  3: 0] custom_dma_burst_2_upstream_current_burst_minus_one;
  wire             custom_dma_burst_2_upstream_debugaccess;
  wire             custom_dma_burst_2_upstream_end_xfer;
  wire             custom_dma_burst_2_upstream_firsttransfer;
  wire             custom_dma_burst_2_upstream_grant_vector;
  wire             custom_dma_burst_2_upstream_in_a_read_cycle;
  wire             custom_dma_burst_2_upstream_in_a_write_cycle;
  reg              custom_dma_burst_2_upstream_load_fifo;
  wire             custom_dma_burst_2_upstream_master_qreq_vector;
  wire             custom_dma_burst_2_upstream_move_on_to_next_transaction;
  wire    [  2: 0] custom_dma_burst_2_upstream_next_bbt_burstcount;
  wire    [  3: 0] custom_dma_burst_2_upstream_next_burst_count;
  wire             custom_dma_burst_2_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_2_upstream_read;
  wire    [ 31: 0] custom_dma_burst_2_upstream_readdata_from_sa;
  wire             custom_dma_burst_2_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_2_upstream_reg_firsttransfer;
  wire    [  3: 0] custom_dma_burst_2_upstream_selected_burstcount;
  reg              custom_dma_burst_2_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_2_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_2_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] custom_dma_burst_2_upstream_transaction_burst_count;
  wire             custom_dma_burst_2_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_2_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_2_upstream_waits_for_read;
  wire             custom_dma_burst_2_upstream_waits_for_write;
  wire             custom_dma_burst_2_upstream_write;
  wire    [ 31: 0] custom_dma_burst_2_upstream_writedata;
  reg              d1_custom_dma_burst_2_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_custom_dma_burst_2_upstream_load_fifo;
  wire             wait_for_custom_dma_burst_2_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_2_upstream_end_xfer;
    end


  assign custom_dma_burst_2_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_custom_dma_burst_2_upstream));
  //assign custom_dma_burst_2_upstream_readdatavalid_from_sa = custom_dma_burst_2_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_2_upstream_readdatavalid_from_sa = custom_dma_burst_2_upstream_readdatavalid;

  //assign custom_dma_burst_2_upstream_readdata_from_sa = custom_dma_burst_2_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_2_upstream_readdata_from_sa = custom_dma_burst_2_upstream_readdata;

  assign cpu_data_master_requests_custom_dma_burst_2_upstream = ({cpu_data_master_address_to_slave[26 : 12] , 12'b0} == 27'h5000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign custom_dma_burst_2_upstream_waitrequest_from_sa = custom_dma_burst_2_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_2_upstream_waitrequest_from_sa = custom_dma_burst_2_upstream_waitrequest;

  //custom_dma_burst_2_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_2_upstream_arb_share_set_values = (cpu_data_master_granted_custom_dma_burst_2_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //custom_dma_burst_2_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_2_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_2_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_2_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_custom_dma_burst_2_upstream;

  //custom_dma_burst_2_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_2_upstream_arb_share_counter_next_value = custom_dma_burst_2_upstream_firsttransfer ? (custom_dma_burst_2_upstream_arb_share_set_values - 1) : |custom_dma_burst_2_upstream_arb_share_counter ? (custom_dma_burst_2_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_2_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_2_upstream_allgrants = |custom_dma_burst_2_upstream_grant_vector;

  //custom_dma_burst_2_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_2_upstream_end_xfer = ~(custom_dma_burst_2_upstream_waits_for_read | custom_dma_burst_2_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream = custom_dma_burst_2_upstream_end_xfer & (~custom_dma_burst_2_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_2_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_2_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream & custom_dma_burst_2_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream & ~custom_dma_burst_2_upstream_non_bursting_master_requests);

  //custom_dma_burst_2_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_2_upstream_arb_counter_enable)
          custom_dma_burst_2_upstream_arb_share_counter <= custom_dma_burst_2_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_2_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_2_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_2_upstream & ~custom_dma_burst_2_upstream_non_bursting_master_requests))
          custom_dma_burst_2_upstream_slavearbiterlockenable <= |custom_dma_burst_2_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master custom_dma_burst_2/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = custom_dma_burst_2_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //custom_dma_burst_2_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_2_upstream_slavearbiterlockenable2 = |custom_dma_burst_2_upstream_arb_share_counter_next_value;

  //cpu/data_master custom_dma_burst_2/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = custom_dma_burst_2_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //custom_dma_burst_2_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_2_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_custom_dma_burst_2_upstream = cpu_data_master_requests_custom_dma_burst_2_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register) | (|cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register))));
  //unique name for custom_dma_burst_2_upstream_move_on_to_next_transaction, which is an e_assign
  assign custom_dma_burst_2_upstream_move_on_to_next_transaction = custom_dma_burst_2_upstream_this_cycle_is_the_last_burst & custom_dma_burst_2_upstream_load_fifo;

  //the currently selected burstcount for custom_dma_burst_2_upstream, which is an e_mux
  assign custom_dma_burst_2_upstream_selected_burstcount = (cpu_data_master_granted_custom_dma_burst_2_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_custom_dma_burst_2_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_custom_dma_burst_2_upstream_module burstcount_fifo_for_custom_dma_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_2_upstream_selected_burstcount),
      .data_out             (custom_dma_burst_2_upstream_transaction_burst_count),
      .empty                (custom_dma_burst_2_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (custom_dma_burst_2_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read & custom_dma_burst_2_upstream_load_fifo & ~(custom_dma_burst_2_upstream_this_cycle_is_the_last_burst & custom_dma_burst_2_upstream_burstcount_fifo_empty))
    );

  //custom_dma_burst_2_upstream current burst minus one, which is an e_assign
  assign custom_dma_burst_2_upstream_current_burst_minus_one = custom_dma_burst_2_upstream_current_burst - 1;

  //what to load in current_burst, for custom_dma_burst_2_upstream, which is an e_mux
  assign custom_dma_burst_2_upstream_next_burst_count = (((in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read) & ~custom_dma_burst_2_upstream_load_fifo))? custom_dma_burst_2_upstream_selected_burstcount :
    ((in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read & custom_dma_burst_2_upstream_this_cycle_is_the_last_burst & custom_dma_burst_2_upstream_burstcount_fifo_empty))? custom_dma_burst_2_upstream_selected_burstcount :
    (custom_dma_burst_2_upstream_this_cycle_is_the_last_burst)? custom_dma_burst_2_upstream_transaction_burst_count :
    custom_dma_burst_2_upstream_current_burst_minus_one;

  //the current burst count for custom_dma_burst_2_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_current_burst <= 0;
      else if (custom_dma_burst_2_upstream_readdatavalid_from_sa | (~custom_dma_burst_2_upstream_load_fifo & (in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read)))
          custom_dma_burst_2_upstream_current_burst <= custom_dma_burst_2_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_custom_dma_burst_2_upstream_load_fifo = (~custom_dma_burst_2_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read) & custom_dma_burst_2_upstream_load_fifo))? 1 :
    ~custom_dma_burst_2_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read) & ~custom_dma_burst_2_upstream_load_fifo | custom_dma_burst_2_upstream_this_cycle_is_the_last_burst)
          custom_dma_burst_2_upstream_load_fifo <= p0_custom_dma_burst_2_upstream_load_fifo;
    end


  //the last cycle in the burst for custom_dma_burst_2_upstream, which is an e_assign
  assign custom_dma_burst_2_upstream_this_cycle_is_the_last_burst = ~(|custom_dma_burst_2_upstream_current_burst_minus_one) & custom_dma_burst_2_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_custom_dma_burst_2_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_custom_dma_burst_2_upstream_module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_2_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_custom_dma_burst_2_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_custom_dma_burst_2_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_custom_dma_burst_2_upstream),
      .full                 (),
      .read                 (custom_dma_burst_2_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_2_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_custom_dma_burst_2_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_custom_dma_burst_2_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_custom_dma_burst_2_upstream = custom_dma_burst_2_upstream_readdatavalid_from_sa;

  //custom_dma_burst_2_upstream_writedata mux, which is an e_mux
  assign custom_dma_burst_2_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for custom_dma_burst_2/upstream, which is an e_mux
  assign custom_dma_burst_2_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_custom_dma_burst_2_upstream = cpu_data_master_qualified_request_custom_dma_burst_2_upstream;

  //cpu/data_master saved-grant custom_dma_burst_2/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_custom_dma_burst_2_upstream = cpu_data_master_requests_custom_dma_burst_2_upstream;

  //allow new arb cycle for custom_dma_burst_2/upstream, which is an e_assign
  assign custom_dma_burst_2_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_2_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_2_upstream_master_qreq_vector = 1;

  //custom_dma_burst_2_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_2_upstream_firsttransfer = custom_dma_burst_2_upstream_begins_xfer ? custom_dma_burst_2_upstream_unreg_firsttransfer : custom_dma_burst_2_upstream_reg_firsttransfer;

  //custom_dma_burst_2_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_2_upstream_unreg_firsttransfer = ~(custom_dma_burst_2_upstream_slavearbiterlockenable & custom_dma_burst_2_upstream_any_continuerequest);

  //custom_dma_burst_2_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_2_upstream_begins_xfer)
          custom_dma_burst_2_upstream_reg_firsttransfer <= custom_dma_burst_2_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_2_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign custom_dma_burst_2_upstream_next_bbt_burstcount = ((((custom_dma_burst_2_upstream_write) && (custom_dma_burst_2_upstream_bbt_burstcounter == 0))))? (custom_dma_burst_2_upstream_burstcount - 1) :
    ((((custom_dma_burst_2_upstream_read) && (custom_dma_burst_2_upstream_bbt_burstcounter == 0))))? 0 :
    (custom_dma_burst_2_upstream_bbt_burstcounter - 1);

  //custom_dma_burst_2_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_upstream_bbt_burstcounter <= 0;
      else if (custom_dma_burst_2_upstream_begins_xfer)
          custom_dma_burst_2_upstream_bbt_burstcounter <= custom_dma_burst_2_upstream_next_bbt_burstcount;
    end


  //custom_dma_burst_2_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_2_upstream_beginbursttransfer_internal = custom_dma_burst_2_upstream_begins_xfer & (custom_dma_burst_2_upstream_bbt_burstcounter == 0);

  //custom_dma_burst_2_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_2_upstream_read = cpu_data_master_granted_custom_dma_burst_2_upstream & cpu_data_master_read;

  //custom_dma_burst_2_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_2_upstream_write = cpu_data_master_granted_custom_dma_burst_2_upstream & cpu_data_master_write;

  //custom_dma_burst_2_upstream_address mux, which is an e_mux
  assign custom_dma_burst_2_upstream_address = cpu_data_master_address_to_slave;

  //d1_custom_dma_burst_2_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_2_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_2_upstream_end_xfer <= custom_dma_burst_2_upstream_end_xfer;
    end


  //custom_dma_burst_2_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_2_upstream_waits_for_read = custom_dma_burst_2_upstream_in_a_read_cycle & custom_dma_burst_2_upstream_waitrequest_from_sa;

  //custom_dma_burst_2_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_2_upstream_in_a_read_cycle = cpu_data_master_granted_custom_dma_burst_2_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_2_upstream_in_a_read_cycle;

  //custom_dma_burst_2_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_2_upstream_waits_for_write = custom_dma_burst_2_upstream_in_a_write_cycle & custom_dma_burst_2_upstream_waitrequest_from_sa;

  //custom_dma_burst_2_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_2_upstream_in_a_write_cycle = cpu_data_master_granted_custom_dma_burst_2_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_2_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_2_upstream_counter = 0;
  //custom_dma_burst_2_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_2_upstream_byteenable = (cpu_data_master_granted_custom_dma_burst_2_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign custom_dma_burst_2_upstream_burstcount = (cpu_data_master_granted_custom_dma_burst_2_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_2_upstream_debugaccess = (cpu_data_master_granted_custom_dma_burst_2_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_2/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_custom_dma_burst_2_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_2/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_2_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_2_downstream_address,
                                                   custom_dma_burst_2_downstream_burstcount,
                                                   custom_dma_burst_2_downstream_byteenable,
                                                   custom_dma_burst_2_downstream_granted_pipeline_bridge_s1,
                                                   custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1,
                                                   custom_dma_burst_2_downstream_read,
                                                   custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1,
                                                   custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register,
                                                   custom_dma_burst_2_downstream_requests_pipeline_bridge_s1,
                                                   custom_dma_burst_2_downstream_write,
                                                   custom_dma_burst_2_downstream_writedata,
                                                   d1_pipeline_bridge_s1_end_xfer,
                                                   pipeline_bridge_s1_readdata_from_sa,
                                                   pipeline_bridge_s1_waitrequest_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_2_downstream_address_to_slave,
                                                   custom_dma_burst_2_downstream_latency_counter,
                                                   custom_dma_burst_2_downstream_readdata,
                                                   custom_dma_burst_2_downstream_readdatavalid,
                                                   custom_dma_burst_2_downstream_reset_n,
                                                   custom_dma_burst_2_downstream_waitrequest
                                                )
;

  output  [ 11: 0] custom_dma_burst_2_downstream_address_to_slave;
  output           custom_dma_burst_2_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_2_downstream_readdata;
  output           custom_dma_burst_2_downstream_readdatavalid;
  output           custom_dma_burst_2_downstream_reset_n;
  output           custom_dma_burst_2_downstream_waitrequest;
  input            clk;
  input   [ 11: 0] custom_dma_burst_2_downstream_address;
  input            custom_dma_burst_2_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_2_downstream_byteenable;
  input            custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;
  input            custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1;
  input            custom_dma_burst_2_downstream_read;
  input            custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1;
  input            custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  input            custom_dma_burst_2_downstream_requests_pipeline_bridge_s1;
  input            custom_dma_burst_2_downstream_write;
  input   [ 31: 0] custom_dma_burst_2_downstream_writedata;
  input            d1_pipeline_bridge_s1_end_xfer;
  input   [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  input            pipeline_bridge_s1_waitrequest_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 11: 0] custom_dma_burst_2_downstream_address_last_time;
  wire    [ 11: 0] custom_dma_burst_2_downstream_address_to_slave;
  reg              custom_dma_burst_2_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_2_downstream_byteenable_last_time;
  wire             custom_dma_burst_2_downstream_is_granted_some_slave;
  reg              custom_dma_burst_2_downstream_latency_counter;
  reg              custom_dma_burst_2_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_2_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_2_downstream_readdata;
  wire             custom_dma_burst_2_downstream_readdatavalid;
  wire             custom_dma_burst_2_downstream_reset_n;
  wire             custom_dma_burst_2_downstream_run;
  wire             custom_dma_burst_2_downstream_waitrequest;
  reg              custom_dma_burst_2_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_2_downstream_writedata_last_time;
  wire             latency_load_value;
  wire             p1_custom_dma_burst_2_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_2_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1 | ~custom_dma_burst_2_downstream_requests_pipeline_bridge_s1) & (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 | ~custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1) & ((~custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1 | ~(custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write)))) & ((~custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1 | ~(custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write) | (1 & ~pipeline_bridge_s1_waitrequest_from_sa & (custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_2_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_2_downstream_address_to_slave = custom_dma_burst_2_downstream_address;

  //custom_dma_burst_2_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_2_downstream_read_but_no_slave_selected <= custom_dma_burst_2_downstream_read & custom_dma_burst_2_downstream_run & ~custom_dma_burst_2_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_2_downstream_is_granted_some_slave = custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_2_downstream_readdatavalid = custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_2_downstream_readdatavalid = custom_dma_burst_2_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_2_downstream_readdatavalid;

  //custom_dma_burst_2/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_2_downstream_readdata = pipeline_bridge_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_2_downstream_waitrequest = ~custom_dma_burst_2_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_2_downstream_latency_counter <= p1_custom_dma_burst_2_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_2_downstream_latency_counter = ((custom_dma_burst_2_downstream_run & custom_dma_burst_2_downstream_read))? latency_load_value :
    (custom_dma_burst_2_downstream_latency_counter)? custom_dma_burst_2_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //custom_dma_burst_2_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_2_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_2_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_address_last_time <= custom_dma_burst_2_downstream_address;
    end


  //custom_dma_burst_2/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_2_downstream_waitrequest & (custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write);
    end


  //custom_dma_burst_2_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_address != custom_dma_burst_2_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_2_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_burstcount_last_time <= custom_dma_burst_2_downstream_burstcount;
    end


  //custom_dma_burst_2_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_burstcount != custom_dma_burst_2_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_2_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_byteenable_last_time <= custom_dma_burst_2_downstream_byteenable;
    end


  //custom_dma_burst_2_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_byteenable != custom_dma_burst_2_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_2_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_read_last_time <= custom_dma_burst_2_downstream_read;
    end


  //custom_dma_burst_2_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_read != custom_dma_burst_2_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_2_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_write_last_time <= custom_dma_burst_2_downstream_write;
    end


  //custom_dma_burst_2_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_write != custom_dma_burst_2_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_2_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_2_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_2_downstream_writedata_last_time <= custom_dma_burst_2_downstream_writedata;
    end


  //custom_dma_burst_2_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_2_downstream_writedata != custom_dma_burst_2_downstream_writedata_last_time) & custom_dma_burst_2_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_2_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_custom_dma_burst_3_upstream_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  wire             full_18;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_17;
  assign empty = !full_0;
  assign full_18 = 0;
  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    0;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_3_upstream_module (
                                                                                   // inputs:
                                                                                    clear_fifo,
                                                                                    clk,
                                                                                    data_in,
                                                                                    read,
                                                                                    reset_n,
                                                                                    sync_reset,
                                                                                    write,

                                                                                   // outputs:
                                                                                    data_out,
                                                                                    empty,
                                                                                    fifo_contains_ones_n,
                                                                                    full
                                                                                 )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  wire             full_18;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_17;
  assign empty = !full_0;
  assign full_18 = 0;
  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    0;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_3_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_instruction_master_address_to_slave,
                                                 cpu_instruction_master_burstcount,
                                                 cpu_instruction_master_latency_counter,
                                                 cpu_instruction_master_read,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register,
                                                 custom_dma_burst_3_upstream_readdata,
                                                 custom_dma_burst_3_upstream_readdatavalid,
                                                 custom_dma_burst_3_upstream_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_instruction_master_granted_custom_dma_burst_3_upstream,
                                                 cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream,
                                                 cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register,
                                                 cpu_instruction_master_requests_custom_dma_burst_3_upstream,
                                                 custom_dma_burst_3_upstream_address,
                                                 custom_dma_burst_3_upstream_byteaddress,
                                                 custom_dma_burst_3_upstream_byteenable,
                                                 custom_dma_burst_3_upstream_debugaccess,
                                                 custom_dma_burst_3_upstream_read,
                                                 custom_dma_burst_3_upstream_readdata_from_sa,
                                                 custom_dma_burst_3_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_3_upstream_write,
                                                 d1_custom_dma_burst_3_upstream_end_xfer
                                              )
;

  output           cpu_instruction_master_granted_custom_dma_burst_3_upstream;
  output           cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream;
  output           cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream;
  output           cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register;
  output           cpu_instruction_master_requests_custom_dma_burst_3_upstream;
  output  [ 24: 0] custom_dma_burst_3_upstream_address;
  output  [ 26: 0] custom_dma_burst_3_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_3_upstream_byteenable;
  output           custom_dma_burst_3_upstream_debugaccess;
  output           custom_dma_burst_3_upstream_read;
  output  [ 31: 0] custom_dma_burst_3_upstream_readdata_from_sa;
  output           custom_dma_burst_3_upstream_waitrequest_from_sa;
  output           custom_dma_burst_3_upstream_write;
  output           d1_custom_dma_burst_3_upstream_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_instruction_master_address_to_slave;
  input   [  3: 0] cpu_instruction_master_burstcount;
  input            cpu_instruction_master_latency_counter;
  input            cpu_instruction_master_read;
  input            cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register;
  input   [ 31: 0] custom_dma_burst_3_upstream_readdata;
  input            custom_dma_burst_3_upstream_readdatavalid;
  input            custom_dma_burst_3_upstream_waitrequest;
  input            reset_n;

  wire             cpu_instruction_master_arbiterlock;
  wire             cpu_instruction_master_arbiterlock2;
  wire             cpu_instruction_master_continuerequest;
  wire             cpu_instruction_master_granted_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_rdv_fifo_output_from_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register;
  wire             cpu_instruction_master_requests_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_saved_grant_custom_dma_burst_3_upstream;
  wire    [ 24: 0] custom_dma_burst_3_upstream_address;
  wire             custom_dma_burst_3_upstream_allgrants;
  wire             custom_dma_burst_3_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_3_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_3_upstream_any_continuerequest;
  wire             custom_dma_burst_3_upstream_arb_counter_enable;
  reg     [  3: 0] custom_dma_burst_3_upstream_arb_share_counter;
  wire    [  3: 0] custom_dma_burst_3_upstream_arb_share_counter_next_value;
  wire    [  3: 0] custom_dma_burst_3_upstream_arb_share_set_values;
  wire             custom_dma_burst_3_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_3_upstream_begins_xfer;
  wire             custom_dma_burst_3_upstream_burstcount_fifo_empty;
  wire    [ 26: 0] custom_dma_burst_3_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_3_upstream_byteenable;
  reg     [  3: 0] custom_dma_burst_3_upstream_current_burst;
  wire    [  3: 0] custom_dma_burst_3_upstream_current_burst_minus_one;
  wire             custom_dma_burst_3_upstream_debugaccess;
  wire             custom_dma_burst_3_upstream_end_xfer;
  wire             custom_dma_burst_3_upstream_firsttransfer;
  wire             custom_dma_burst_3_upstream_grant_vector;
  wire             custom_dma_burst_3_upstream_in_a_read_cycle;
  wire             custom_dma_burst_3_upstream_in_a_write_cycle;
  reg              custom_dma_burst_3_upstream_load_fifo;
  wire             custom_dma_burst_3_upstream_master_qreq_vector;
  wire             custom_dma_burst_3_upstream_move_on_to_next_transaction;
  wire    [  3: 0] custom_dma_burst_3_upstream_next_burst_count;
  wire             custom_dma_burst_3_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_3_upstream_read;
  wire    [ 31: 0] custom_dma_burst_3_upstream_readdata_from_sa;
  wire             custom_dma_burst_3_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_3_upstream_reg_firsttransfer;
  wire    [  3: 0] custom_dma_burst_3_upstream_selected_burstcount;
  reg              custom_dma_burst_3_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_3_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_3_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] custom_dma_burst_3_upstream_transaction_burst_count;
  wire             custom_dma_burst_3_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_3_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_3_upstream_waits_for_read;
  wire             custom_dma_burst_3_upstream_waits_for_write;
  wire             custom_dma_burst_3_upstream_write;
  reg              d1_custom_dma_burst_3_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_custom_dma_burst_3_upstream_load_fifo;
  wire             wait_for_custom_dma_burst_3_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_3_upstream_end_xfer;
    end


  assign custom_dma_burst_3_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream));
  //assign custom_dma_burst_3_upstream_readdatavalid_from_sa = custom_dma_burst_3_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_3_upstream_readdatavalid_from_sa = custom_dma_burst_3_upstream_readdatavalid;

  //assign custom_dma_burst_3_upstream_readdata_from_sa = custom_dma_burst_3_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_3_upstream_readdata_from_sa = custom_dma_burst_3_upstream_readdata;

  assign cpu_instruction_master_requests_custom_dma_burst_3_upstream = (({cpu_instruction_master_address_to_slave[26 : 25] , 25'b0} == 27'h2000000) & (cpu_instruction_master_read)) & cpu_instruction_master_read;
  //assign custom_dma_burst_3_upstream_waitrequest_from_sa = custom_dma_burst_3_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_3_upstream_waitrequest_from_sa = custom_dma_burst_3_upstream_waitrequest;

  //custom_dma_burst_3_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_3_upstream_arb_share_set_values = 1;

  //custom_dma_burst_3_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_3_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_3_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_3_upstream_any_bursting_master_saved_grant = cpu_instruction_master_saved_grant_custom_dma_burst_3_upstream;

  //custom_dma_burst_3_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_3_upstream_arb_share_counter_next_value = custom_dma_burst_3_upstream_firsttransfer ? (custom_dma_burst_3_upstream_arb_share_set_values - 1) : |custom_dma_burst_3_upstream_arb_share_counter ? (custom_dma_burst_3_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_3_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_3_upstream_allgrants = |custom_dma_burst_3_upstream_grant_vector;

  //custom_dma_burst_3_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_3_upstream_end_xfer = ~(custom_dma_burst_3_upstream_waits_for_read | custom_dma_burst_3_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream = custom_dma_burst_3_upstream_end_xfer & (~custom_dma_burst_3_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_3_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_3_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream & custom_dma_burst_3_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream & ~custom_dma_burst_3_upstream_non_bursting_master_requests);

  //custom_dma_burst_3_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_3_upstream_arb_counter_enable)
          custom_dma_burst_3_upstream_arb_share_counter <= custom_dma_burst_3_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_3_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_3_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_3_upstream & ~custom_dma_burst_3_upstream_non_bursting_master_requests))
          custom_dma_burst_3_upstream_slavearbiterlockenable <= |custom_dma_burst_3_upstream_arb_share_counter_next_value;
    end


  //cpu/instruction_master custom_dma_burst_3/upstream arbiterlock, which is an e_assign
  assign cpu_instruction_master_arbiterlock = custom_dma_burst_3_upstream_slavearbiterlockenable & cpu_instruction_master_continuerequest;

  //custom_dma_burst_3_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_3_upstream_slavearbiterlockenable2 = |custom_dma_burst_3_upstream_arb_share_counter_next_value;

  //cpu/instruction_master custom_dma_burst_3/upstream arbiterlock2, which is an e_assign
  assign cpu_instruction_master_arbiterlock2 = custom_dma_burst_3_upstream_slavearbiterlockenable2 & cpu_instruction_master_continuerequest;

  //custom_dma_burst_3_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_3_upstream_any_continuerequest = 1;

  //cpu_instruction_master_continuerequest continued request, which is an e_assign
  assign cpu_instruction_master_continuerequest = 1;

  assign cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream = cpu_instruction_master_requests_custom_dma_burst_3_upstream & ~((cpu_instruction_master_read & ((cpu_instruction_master_latency_counter != 0) | (1 < cpu_instruction_master_latency_counter) | (|cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register))));
  //unique name for custom_dma_burst_3_upstream_move_on_to_next_transaction, which is an e_assign
  assign custom_dma_burst_3_upstream_move_on_to_next_transaction = custom_dma_burst_3_upstream_this_cycle_is_the_last_burst & custom_dma_burst_3_upstream_load_fifo;

  //the currently selected burstcount for custom_dma_burst_3_upstream, which is an e_mux
  assign custom_dma_burst_3_upstream_selected_burstcount = (cpu_instruction_master_granted_custom_dma_burst_3_upstream)? cpu_instruction_master_burstcount :
    1;

  //burstcount_fifo_for_custom_dma_burst_3_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_custom_dma_burst_3_upstream_module burstcount_fifo_for_custom_dma_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_3_upstream_selected_burstcount),
      .data_out             (custom_dma_burst_3_upstream_transaction_burst_count),
      .empty                (custom_dma_burst_3_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (custom_dma_burst_3_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read & custom_dma_burst_3_upstream_load_fifo & ~(custom_dma_burst_3_upstream_this_cycle_is_the_last_burst & custom_dma_burst_3_upstream_burstcount_fifo_empty))
    );

  //custom_dma_burst_3_upstream current burst minus one, which is an e_assign
  assign custom_dma_burst_3_upstream_current_burst_minus_one = custom_dma_burst_3_upstream_current_burst - 1;

  //what to load in current_burst, for custom_dma_burst_3_upstream, which is an e_mux
  assign custom_dma_burst_3_upstream_next_burst_count = (((in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read) & ~custom_dma_burst_3_upstream_load_fifo))? custom_dma_burst_3_upstream_selected_burstcount :
    ((in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read & custom_dma_burst_3_upstream_this_cycle_is_the_last_burst & custom_dma_burst_3_upstream_burstcount_fifo_empty))? custom_dma_burst_3_upstream_selected_burstcount :
    (custom_dma_burst_3_upstream_this_cycle_is_the_last_burst)? custom_dma_burst_3_upstream_transaction_burst_count :
    custom_dma_burst_3_upstream_current_burst_minus_one;

  //the current burst count for custom_dma_burst_3_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_upstream_current_burst <= 0;
      else if (custom_dma_burst_3_upstream_readdatavalid_from_sa | (~custom_dma_burst_3_upstream_load_fifo & (in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read)))
          custom_dma_burst_3_upstream_current_burst <= custom_dma_burst_3_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_custom_dma_burst_3_upstream_load_fifo = (~custom_dma_burst_3_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read) & custom_dma_burst_3_upstream_load_fifo))? 1 :
    ~custom_dma_burst_3_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read) & ~custom_dma_burst_3_upstream_load_fifo | custom_dma_burst_3_upstream_this_cycle_is_the_last_burst)
          custom_dma_burst_3_upstream_load_fifo <= p0_custom_dma_burst_3_upstream_load_fifo;
    end


  //the last cycle in the burst for custom_dma_burst_3_upstream, which is an e_assign
  assign custom_dma_burst_3_upstream_this_cycle_is_the_last_burst = ~(|custom_dma_burst_3_upstream_current_burst_minus_one) & custom_dma_burst_3_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_3_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_3_upstream_module rdv_fifo_for_cpu_instruction_master_to_custom_dma_burst_3_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_instruction_master_granted_custom_dma_burst_3_upstream),
      .data_out             (cpu_instruction_master_rdv_fifo_output_from_custom_dma_burst_3_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_3_upstream),
      .full                 (),
      .read                 (custom_dma_burst_3_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_3_upstream_waits_for_read)
    );

  assign cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register = ~cpu_instruction_master_rdv_fifo_empty_custom_dma_burst_3_upstream;
  //local readdatavalid cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream, which is an e_mux
  assign cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream = custom_dma_burst_3_upstream_readdatavalid_from_sa;

  //byteaddress mux for custom_dma_burst_3/upstream, which is an e_mux
  assign custom_dma_burst_3_upstream_byteaddress = cpu_instruction_master_address_to_slave;

  //master is always granted when requested
  assign cpu_instruction_master_granted_custom_dma_burst_3_upstream = cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream;

  //cpu/instruction_master saved-grant custom_dma_burst_3/upstream, which is an e_assign
  assign cpu_instruction_master_saved_grant_custom_dma_burst_3_upstream = cpu_instruction_master_requests_custom_dma_burst_3_upstream;

  //allow new arb cycle for custom_dma_burst_3/upstream, which is an e_assign
  assign custom_dma_burst_3_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_3_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_3_upstream_master_qreq_vector = 1;

  //custom_dma_burst_3_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_3_upstream_firsttransfer = custom_dma_burst_3_upstream_begins_xfer ? custom_dma_burst_3_upstream_unreg_firsttransfer : custom_dma_burst_3_upstream_reg_firsttransfer;

  //custom_dma_burst_3_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_3_upstream_unreg_firsttransfer = ~(custom_dma_burst_3_upstream_slavearbiterlockenable & custom_dma_burst_3_upstream_any_continuerequest);

  //custom_dma_burst_3_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_3_upstream_begins_xfer)
          custom_dma_burst_3_upstream_reg_firsttransfer <= custom_dma_burst_3_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_3_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_3_upstream_beginbursttransfer_internal = custom_dma_burst_3_upstream_begins_xfer;

  //custom_dma_burst_3_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_3_upstream_read = cpu_instruction_master_granted_custom_dma_burst_3_upstream & cpu_instruction_master_read;

  //custom_dma_burst_3_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_3_upstream_write = 0;

  //custom_dma_burst_3_upstream_address mux, which is an e_mux
  assign custom_dma_burst_3_upstream_address = cpu_instruction_master_address_to_slave;

  //d1_custom_dma_burst_3_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_3_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_3_upstream_end_xfer <= custom_dma_burst_3_upstream_end_xfer;
    end


  //custom_dma_burst_3_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_3_upstream_waits_for_read = custom_dma_burst_3_upstream_in_a_read_cycle & custom_dma_burst_3_upstream_waitrequest_from_sa;

  //custom_dma_burst_3_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_3_upstream_in_a_read_cycle = cpu_instruction_master_granted_custom_dma_burst_3_upstream & cpu_instruction_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_3_upstream_in_a_read_cycle;

  //custom_dma_burst_3_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_3_upstream_waits_for_write = custom_dma_burst_3_upstream_in_a_write_cycle & custom_dma_burst_3_upstream_waitrequest_from_sa;

  //custom_dma_burst_3_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_3_upstream_in_a_write_cycle = 0;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_3_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_3_upstream_counter = 0;
  //custom_dma_burst_3_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_3_upstream_byteenable = -1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_3_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_3/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu/instruction_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_instruction_master_requests_custom_dma_burst_3_upstream && (cpu_instruction_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/instruction_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_3/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_3_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_3_downstream_address,
                                                   custom_dma_burst_3_downstream_burstcount,
                                                   custom_dma_burst_3_downstream_byteenable,
                                                   custom_dma_burst_3_downstream_granted_ddr_sdram_s1,
                                                   custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1,
                                                   custom_dma_burst_3_downstream_read,
                                                   custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1,
                                                   custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                                   custom_dma_burst_3_downstream_requests_ddr_sdram_s1,
                                                   custom_dma_burst_3_downstream_write,
                                                   custom_dma_burst_3_downstream_writedata,
                                                   d1_ddr_sdram_s1_end_xfer,
                                                   ddr_sdram_s1_readdata_from_sa,
                                                   ddr_sdram_s1_waitrequest_n_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_3_downstream_address_to_slave,
                                                   custom_dma_burst_3_downstream_latency_counter,
                                                   custom_dma_burst_3_downstream_readdata,
                                                   custom_dma_burst_3_downstream_readdatavalid,
                                                   custom_dma_burst_3_downstream_reset_n,
                                                   custom_dma_burst_3_downstream_waitrequest
                                                )
;

  output  [ 24: 0] custom_dma_burst_3_downstream_address_to_slave;
  output           custom_dma_burst_3_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_3_downstream_readdata;
  output           custom_dma_burst_3_downstream_readdatavalid;
  output           custom_dma_burst_3_downstream_reset_n;
  output           custom_dma_burst_3_downstream_waitrequest;
  input            clk;
  input   [ 24: 0] custom_dma_burst_3_downstream_address;
  input   [  2: 0] custom_dma_burst_3_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_3_downstream_byteenable;
  input            custom_dma_burst_3_downstream_granted_ddr_sdram_s1;
  input            custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1;
  input            custom_dma_burst_3_downstream_read;
  input            custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1;
  input            custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  input            custom_dma_burst_3_downstream_requests_ddr_sdram_s1;
  input            custom_dma_burst_3_downstream_write;
  input   [ 31: 0] custom_dma_burst_3_downstream_writedata;
  input            d1_ddr_sdram_s1_end_xfer;
  input   [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  input            ddr_sdram_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] custom_dma_burst_3_downstream_address_last_time;
  wire    [ 24: 0] custom_dma_burst_3_downstream_address_to_slave;
  reg     [  2: 0] custom_dma_burst_3_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_3_downstream_byteenable_last_time;
  wire             custom_dma_burst_3_downstream_is_granted_some_slave;
  reg              custom_dma_burst_3_downstream_latency_counter;
  reg              custom_dma_burst_3_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_3_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_3_downstream_readdata;
  wire             custom_dma_burst_3_downstream_readdatavalid;
  wire             custom_dma_burst_3_downstream_reset_n;
  wire             custom_dma_burst_3_downstream_run;
  wire             custom_dma_burst_3_downstream_waitrequest;
  reg              custom_dma_burst_3_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_3_downstream_writedata_last_time;
  wire             latency_load_value;
  wire             p1_custom_dma_burst_3_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_3_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1 | ~custom_dma_burst_3_downstream_requests_ddr_sdram_s1) & (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 | ~custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1) & ((~custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write)))) & ((~custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_3_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_3_downstream_address_to_slave = custom_dma_burst_3_downstream_address;

  //custom_dma_burst_3_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_3_downstream_read_but_no_slave_selected <= custom_dma_burst_3_downstream_read & custom_dma_burst_3_downstream_run & ~custom_dma_burst_3_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_3_downstream_is_granted_some_slave = custom_dma_burst_3_downstream_granted_ddr_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_3_downstream_readdatavalid = custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_3_downstream_readdatavalid = custom_dma_burst_3_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_3_downstream_readdatavalid;

  //custom_dma_burst_3/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_3_downstream_readdata = ddr_sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_3_downstream_waitrequest = ~custom_dma_burst_3_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_3_downstream_latency_counter <= p1_custom_dma_burst_3_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_3_downstream_latency_counter = ((custom_dma_burst_3_downstream_run & custom_dma_burst_3_downstream_read))? latency_load_value :
    (custom_dma_burst_3_downstream_latency_counter)? custom_dma_burst_3_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //custom_dma_burst_3_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_3_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_3_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_address_last_time <= custom_dma_burst_3_downstream_address;
    end


  //custom_dma_burst_3/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_3_downstream_waitrequest & (custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write);
    end


  //custom_dma_burst_3_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_address != custom_dma_burst_3_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_3_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_burstcount_last_time <= custom_dma_burst_3_downstream_burstcount;
    end


  //custom_dma_burst_3_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_burstcount != custom_dma_burst_3_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_3_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_byteenable_last_time <= custom_dma_burst_3_downstream_byteenable;
    end


  //custom_dma_burst_3_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_byteenable != custom_dma_burst_3_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_3_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_read_last_time <= custom_dma_burst_3_downstream_read;
    end


  //custom_dma_burst_3_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_read != custom_dma_burst_3_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_3_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_write_last_time <= custom_dma_burst_3_downstream_write;
    end


  //custom_dma_burst_3_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_write != custom_dma_burst_3_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_3_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_3_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_3_downstream_writedata_last_time <= custom_dma_burst_3_downstream_writedata;
    end


  //custom_dma_burst_3_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_3_downstream_writedata != custom_dma_burst_3_downstream_writedata_last_time) & custom_dma_burst_3_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_3_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_custom_dma_burst_4_upstream_module (
                                                                // inputs:
                                                                 clear_fifo,
                                                                 clk,
                                                                 data_in,
                                                                 read,
                                                                 reset_n,
                                                                 sync_reset,
                                                                 write,

                                                                // outputs:
                                                                 data_out,
                                                                 empty,
                                                                 fifo_contains_ones_n,
                                                                 full
                                                              )
;

  output  [  3: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  3: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  3: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  wire             full_18;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  3: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  3: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  3: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  3: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  3: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  3: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  3: 0] p15_stage_15;
  wire             p16_full_16;
  wire    [  3: 0] p16_stage_16;
  wire             p17_full_17;
  wire    [  3: 0] p17_stage_17;
  wire             p1_full_1;
  wire    [  3: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  3: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  3: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  3: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  3: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  3: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  3: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  3: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  3: 0] p9_stage_9;
  reg     [  3: 0] stage_0;
  reg     [  3: 0] stage_1;
  reg     [  3: 0] stage_10;
  reg     [  3: 0] stage_11;
  reg     [  3: 0] stage_12;
  reg     [  3: 0] stage_13;
  reg     [  3: 0] stage_14;
  reg     [  3: 0] stage_15;
  reg     [  3: 0] stage_16;
  reg     [  3: 0] stage_17;
  reg     [  3: 0] stage_2;
  reg     [  3: 0] stage_3;
  reg     [  3: 0] stage_4;
  reg     [  3: 0] stage_5;
  reg     [  3: 0] stage_6;
  reg     [  3: 0] stage_7;
  reg     [  3: 0] stage_8;
  reg     [  3: 0] stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_17;
  assign empty = !full_0;
  assign full_18 = 0;
  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    0;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_4_upstream_module (
                                                                            // inputs:
                                                                             clear_fifo,
                                                                             clk,
                                                                             data_in,
                                                                             read,
                                                                             reset_n,
                                                                             sync_reset,
                                                                             write,

                                                                            // outputs:
                                                                             data_out,
                                                                             empty,
                                                                             fifo_contains_ones_n,
                                                                             full
                                                                          )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  reg              full_16;
  reg              full_17;
  wire             full_18;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p16_full_16;
  wire             p16_stage_16;
  wire             p17_full_17;
  wire             p17_stage_17;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_16;
  reg              stage_17;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_17;
  assign empty = !full_0;
  assign full_18 = 0;
  //data_17, which is an e_mux
  assign p17_stage_17 = ((full_18 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_17 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_17))
          if (sync_reset & full_17 & !((full_18 == 0) & read & write))
              stage_17 <= 0;
          else 
            stage_17 <= p17_stage_17;
    end


  //control_17, which is an e_mux
  assign p17_full_17 = ((read & !write) == 0)? full_16 :
    0;

  //control_reg_17, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_17 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_17 <= 0;
          else 
            full_17 <= p17_full_17;
    end


  //data_16, which is an e_mux
  assign p16_stage_16 = ((full_17 & ~clear_fifo) == 0)? data_in :
    stage_17;

  //data_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_16 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_16))
          if (sync_reset & full_16 & !((full_17 == 0) & read & write))
              stage_16 <= 0;
          else 
            stage_16 <= p16_stage_16;
    end


  //control_16, which is an e_mux
  assign p16_full_16 = ((read & !write) == 0)? full_15 :
    full_17;

  //control_reg_16, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_16 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_16 <= 0;
          else 
            full_16 <= p16_full_16;
    end


  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    stage_16;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    full_16;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_4_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 cpu_data_master_address_to_slave,
                                                 cpu_data_master_burstcount,
                                                 cpu_data_master_byteenable,
                                                 cpu_data_master_debugaccess,
                                                 cpu_data_master_latency_counter,
                                                 cpu_data_master_read,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register,
                                                 cpu_data_master_write,
                                                 cpu_data_master_writedata,
                                                 custom_dma_burst_4_upstream_readdata,
                                                 custom_dma_burst_4_upstream_readdatavalid,
                                                 custom_dma_burst_4_upstream_waitrequest,
                                                 reset_n,

                                                // outputs:
                                                 cpu_data_master_granted_custom_dma_burst_4_upstream,
                                                 cpu_data_master_qualified_request_custom_dma_burst_4_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_4_upstream,
                                                 cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register,
                                                 cpu_data_master_requests_custom_dma_burst_4_upstream,
                                                 custom_dma_burst_4_upstream_address,
                                                 custom_dma_burst_4_upstream_burstcount,
                                                 custom_dma_burst_4_upstream_byteaddress,
                                                 custom_dma_burst_4_upstream_byteenable,
                                                 custom_dma_burst_4_upstream_debugaccess,
                                                 custom_dma_burst_4_upstream_read,
                                                 custom_dma_burst_4_upstream_readdata_from_sa,
                                                 custom_dma_burst_4_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_4_upstream_write,
                                                 custom_dma_burst_4_upstream_writedata,
                                                 d1_custom_dma_burst_4_upstream_end_xfer
                                              )
;

  output           cpu_data_master_granted_custom_dma_burst_4_upstream;
  output           cpu_data_master_qualified_request_custom_dma_burst_4_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_4_upstream;
  output           cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  output           cpu_data_master_requests_custom_dma_burst_4_upstream;
  output  [ 24: 0] custom_dma_burst_4_upstream_address;
  output  [  3: 0] custom_dma_burst_4_upstream_burstcount;
  output  [ 26: 0] custom_dma_burst_4_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_4_upstream_byteenable;
  output           custom_dma_burst_4_upstream_debugaccess;
  output           custom_dma_burst_4_upstream_read;
  output  [ 31: 0] custom_dma_burst_4_upstream_readdata_from_sa;
  output           custom_dma_burst_4_upstream_waitrequest_from_sa;
  output           custom_dma_burst_4_upstream_write;
  output  [ 31: 0] custom_dma_burst_4_upstream_writedata;
  output           d1_custom_dma_burst_4_upstream_end_xfer;
  input            clk;
  input   [ 26: 0] cpu_data_master_address_to_slave;
  input   [  3: 0] cpu_data_master_burstcount;
  input   [  3: 0] cpu_data_master_byteenable;
  input            cpu_data_master_debugaccess;
  input            cpu_data_master_latency_counter;
  input            cpu_data_master_read;
  input            cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  input            cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  input            cpu_data_master_write;
  input   [ 31: 0] cpu_data_master_writedata;
  input   [ 31: 0] custom_dma_burst_4_upstream_readdata;
  input            custom_dma_burst_4_upstream_readdatavalid;
  input            custom_dma_burst_4_upstream_waitrequest;
  input            reset_n;

  wire             cpu_data_master_arbiterlock;
  wire             cpu_data_master_arbiterlock2;
  wire             cpu_data_master_continuerequest;
  wire             cpu_data_master_granted_custom_dma_burst_4_upstream;
  wire             cpu_data_master_qualified_request_custom_dma_burst_4_upstream;
  wire             cpu_data_master_rdv_fifo_empty_custom_dma_burst_4_upstream;
  wire             cpu_data_master_rdv_fifo_output_from_custom_dma_burst_4_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_4_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  wire             cpu_data_master_requests_custom_dma_burst_4_upstream;
  wire             cpu_data_master_saved_grant_custom_dma_burst_4_upstream;
  wire    [ 24: 0] custom_dma_burst_4_upstream_address;
  wire             custom_dma_burst_4_upstream_allgrants;
  wire             custom_dma_burst_4_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_4_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_4_upstream_any_continuerequest;
  wire             custom_dma_burst_4_upstream_arb_counter_enable;
  reg     [  3: 0] custom_dma_burst_4_upstream_arb_share_counter;
  wire    [  3: 0] custom_dma_burst_4_upstream_arb_share_counter_next_value;
  wire    [  3: 0] custom_dma_burst_4_upstream_arb_share_set_values;
  reg     [  2: 0] custom_dma_burst_4_upstream_bbt_burstcounter;
  wire             custom_dma_burst_4_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_4_upstream_begins_xfer;
  wire    [  3: 0] custom_dma_burst_4_upstream_burstcount;
  wire             custom_dma_burst_4_upstream_burstcount_fifo_empty;
  wire    [ 26: 0] custom_dma_burst_4_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_4_upstream_byteenable;
  reg     [  3: 0] custom_dma_burst_4_upstream_current_burst;
  wire    [  3: 0] custom_dma_burst_4_upstream_current_burst_minus_one;
  wire             custom_dma_burst_4_upstream_debugaccess;
  wire             custom_dma_burst_4_upstream_end_xfer;
  wire             custom_dma_burst_4_upstream_firsttransfer;
  wire             custom_dma_burst_4_upstream_grant_vector;
  wire             custom_dma_burst_4_upstream_in_a_read_cycle;
  wire             custom_dma_burst_4_upstream_in_a_write_cycle;
  reg              custom_dma_burst_4_upstream_load_fifo;
  wire             custom_dma_burst_4_upstream_master_qreq_vector;
  wire             custom_dma_burst_4_upstream_move_on_to_next_transaction;
  wire    [  2: 0] custom_dma_burst_4_upstream_next_bbt_burstcount;
  wire    [  3: 0] custom_dma_burst_4_upstream_next_burst_count;
  wire             custom_dma_burst_4_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_4_upstream_read;
  wire    [ 31: 0] custom_dma_burst_4_upstream_readdata_from_sa;
  wire             custom_dma_burst_4_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_4_upstream_reg_firsttransfer;
  wire    [  3: 0] custom_dma_burst_4_upstream_selected_burstcount;
  reg              custom_dma_burst_4_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_4_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_4_upstream_this_cycle_is_the_last_burst;
  wire    [  3: 0] custom_dma_burst_4_upstream_transaction_burst_count;
  wire             custom_dma_burst_4_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_4_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_4_upstream_waits_for_read;
  wire             custom_dma_burst_4_upstream_waits_for_write;
  wire             custom_dma_burst_4_upstream_write;
  wire    [ 31: 0] custom_dma_burst_4_upstream_writedata;
  reg              d1_custom_dma_burst_4_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p0_custom_dma_burst_4_upstream_load_fifo;
  wire             wait_for_custom_dma_burst_4_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_4_upstream_end_xfer;
    end


  assign custom_dma_burst_4_upstream_begins_xfer = ~d1_reasons_to_wait & ((cpu_data_master_qualified_request_custom_dma_burst_4_upstream));
  //assign custom_dma_burst_4_upstream_readdatavalid_from_sa = custom_dma_burst_4_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_4_upstream_readdatavalid_from_sa = custom_dma_burst_4_upstream_readdatavalid;

  //assign custom_dma_burst_4_upstream_readdata_from_sa = custom_dma_burst_4_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_4_upstream_readdata_from_sa = custom_dma_burst_4_upstream_readdata;

  assign cpu_data_master_requests_custom_dma_burst_4_upstream = ({cpu_data_master_address_to_slave[26 : 25] , 25'b0} == 27'h2000000) & (cpu_data_master_read | cpu_data_master_write);
  //assign custom_dma_burst_4_upstream_waitrequest_from_sa = custom_dma_burst_4_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_4_upstream_waitrequest_from_sa = custom_dma_burst_4_upstream_waitrequest;

  //custom_dma_burst_4_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_4_upstream_arb_share_set_values = (cpu_data_master_granted_custom_dma_burst_4_upstream)? (((cpu_data_master_write) ? cpu_data_master_burstcount : 1)) :
    1;

  //custom_dma_burst_4_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_4_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_4_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_4_upstream_any_bursting_master_saved_grant = cpu_data_master_saved_grant_custom_dma_burst_4_upstream;

  //custom_dma_burst_4_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_4_upstream_arb_share_counter_next_value = custom_dma_burst_4_upstream_firsttransfer ? (custom_dma_burst_4_upstream_arb_share_set_values - 1) : |custom_dma_burst_4_upstream_arb_share_counter ? (custom_dma_burst_4_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_4_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_4_upstream_allgrants = |custom_dma_burst_4_upstream_grant_vector;

  //custom_dma_burst_4_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_4_upstream_end_xfer = ~(custom_dma_burst_4_upstream_waits_for_read | custom_dma_burst_4_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream = custom_dma_burst_4_upstream_end_xfer & (~custom_dma_burst_4_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_4_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_4_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream & custom_dma_burst_4_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream & ~custom_dma_burst_4_upstream_non_bursting_master_requests);

  //custom_dma_burst_4_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_4_upstream_arb_counter_enable)
          custom_dma_burst_4_upstream_arb_share_counter <= custom_dma_burst_4_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_4_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_4_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_4_upstream & ~custom_dma_burst_4_upstream_non_bursting_master_requests))
          custom_dma_burst_4_upstream_slavearbiterlockenable <= |custom_dma_burst_4_upstream_arb_share_counter_next_value;
    end


  //cpu/data_master custom_dma_burst_4/upstream arbiterlock, which is an e_assign
  assign cpu_data_master_arbiterlock = custom_dma_burst_4_upstream_slavearbiterlockenable & cpu_data_master_continuerequest;

  //custom_dma_burst_4_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_4_upstream_slavearbiterlockenable2 = |custom_dma_burst_4_upstream_arb_share_counter_next_value;

  //cpu/data_master custom_dma_burst_4/upstream arbiterlock2, which is an e_assign
  assign cpu_data_master_arbiterlock2 = custom_dma_burst_4_upstream_slavearbiterlockenable2 & cpu_data_master_continuerequest;

  //custom_dma_burst_4_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_4_upstream_any_continuerequest = 1;

  //cpu_data_master_continuerequest continued request, which is an e_assign
  assign cpu_data_master_continuerequest = 1;

  assign cpu_data_master_qualified_request_custom_dma_burst_4_upstream = cpu_data_master_requests_custom_dma_burst_4_upstream & ~((cpu_data_master_read & ((cpu_data_master_latency_counter != 0) | (1 < cpu_data_master_latency_counter) | (|cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register) | (|cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register))));
  //unique name for custom_dma_burst_4_upstream_move_on_to_next_transaction, which is an e_assign
  assign custom_dma_burst_4_upstream_move_on_to_next_transaction = custom_dma_burst_4_upstream_this_cycle_is_the_last_burst & custom_dma_burst_4_upstream_load_fifo;

  //the currently selected burstcount for custom_dma_burst_4_upstream, which is an e_mux
  assign custom_dma_burst_4_upstream_selected_burstcount = (cpu_data_master_granted_custom_dma_burst_4_upstream)? cpu_data_master_burstcount :
    1;

  //burstcount_fifo_for_custom_dma_burst_4_upstream, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_custom_dma_burst_4_upstream_module burstcount_fifo_for_custom_dma_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_4_upstream_selected_burstcount),
      .data_out             (custom_dma_burst_4_upstream_transaction_burst_count),
      .empty                (custom_dma_burst_4_upstream_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (custom_dma_burst_4_upstream_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read & custom_dma_burst_4_upstream_load_fifo & ~(custom_dma_burst_4_upstream_this_cycle_is_the_last_burst & custom_dma_burst_4_upstream_burstcount_fifo_empty))
    );

  //custom_dma_burst_4_upstream current burst minus one, which is an e_assign
  assign custom_dma_burst_4_upstream_current_burst_minus_one = custom_dma_burst_4_upstream_current_burst - 1;

  //what to load in current_burst, for custom_dma_burst_4_upstream, which is an e_mux
  assign custom_dma_burst_4_upstream_next_burst_count = (((in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read) & ~custom_dma_burst_4_upstream_load_fifo))? custom_dma_burst_4_upstream_selected_burstcount :
    ((in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read & custom_dma_burst_4_upstream_this_cycle_is_the_last_burst & custom_dma_burst_4_upstream_burstcount_fifo_empty))? custom_dma_burst_4_upstream_selected_burstcount :
    (custom_dma_burst_4_upstream_this_cycle_is_the_last_burst)? custom_dma_burst_4_upstream_transaction_burst_count :
    custom_dma_burst_4_upstream_current_burst_minus_one;

  //the current burst count for custom_dma_burst_4_upstream, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_current_burst <= 0;
      else if (custom_dma_burst_4_upstream_readdatavalid_from_sa | (~custom_dma_burst_4_upstream_load_fifo & (in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read)))
          custom_dma_burst_4_upstream_current_burst <= custom_dma_burst_4_upstream_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_custom_dma_burst_4_upstream_load_fifo = (~custom_dma_burst_4_upstream_load_fifo)? 1 :
    (((in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read) & custom_dma_burst_4_upstream_load_fifo))? 1 :
    ~custom_dma_burst_4_upstream_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_load_fifo <= 0;
      else if ((in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read) & ~custom_dma_burst_4_upstream_load_fifo | custom_dma_burst_4_upstream_this_cycle_is_the_last_burst)
          custom_dma_burst_4_upstream_load_fifo <= p0_custom_dma_burst_4_upstream_load_fifo;
    end


  //the last cycle in the burst for custom_dma_burst_4_upstream, which is an e_assign
  assign custom_dma_burst_4_upstream_this_cycle_is_the_last_burst = ~(|custom_dma_burst_4_upstream_current_burst_minus_one) & custom_dma_burst_4_upstream_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_data_master_to_custom_dma_burst_4_upstream, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_custom_dma_burst_4_upstream_module rdv_fifo_for_cpu_data_master_to_custom_dma_burst_4_upstream
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_data_master_granted_custom_dma_burst_4_upstream),
      .data_out             (cpu_data_master_rdv_fifo_output_from_custom_dma_burst_4_upstream),
      .empty                (),
      .fifo_contains_ones_n (cpu_data_master_rdv_fifo_empty_custom_dma_burst_4_upstream),
      .full                 (),
      .read                 (custom_dma_burst_4_upstream_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~custom_dma_burst_4_upstream_waits_for_read)
    );

  assign cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register = ~cpu_data_master_rdv_fifo_empty_custom_dma_burst_4_upstream;
  //local readdatavalid cpu_data_master_read_data_valid_custom_dma_burst_4_upstream, which is an e_mux
  assign cpu_data_master_read_data_valid_custom_dma_burst_4_upstream = custom_dma_burst_4_upstream_readdatavalid_from_sa;

  //custom_dma_burst_4_upstream_writedata mux, which is an e_mux
  assign custom_dma_burst_4_upstream_writedata = cpu_data_master_writedata;

  //byteaddress mux for custom_dma_burst_4/upstream, which is an e_mux
  assign custom_dma_burst_4_upstream_byteaddress = cpu_data_master_address_to_slave;

  //master is always granted when requested
  assign cpu_data_master_granted_custom_dma_burst_4_upstream = cpu_data_master_qualified_request_custom_dma_burst_4_upstream;

  //cpu/data_master saved-grant custom_dma_burst_4/upstream, which is an e_assign
  assign cpu_data_master_saved_grant_custom_dma_burst_4_upstream = cpu_data_master_requests_custom_dma_burst_4_upstream;

  //allow new arb cycle for custom_dma_burst_4/upstream, which is an e_assign
  assign custom_dma_burst_4_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_4_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_4_upstream_master_qreq_vector = 1;

  //custom_dma_burst_4_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_4_upstream_firsttransfer = custom_dma_burst_4_upstream_begins_xfer ? custom_dma_burst_4_upstream_unreg_firsttransfer : custom_dma_burst_4_upstream_reg_firsttransfer;

  //custom_dma_burst_4_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_4_upstream_unreg_firsttransfer = ~(custom_dma_burst_4_upstream_slavearbiterlockenable & custom_dma_burst_4_upstream_any_continuerequest);

  //custom_dma_burst_4_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_4_upstream_begins_xfer)
          custom_dma_burst_4_upstream_reg_firsttransfer <= custom_dma_burst_4_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_4_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign custom_dma_burst_4_upstream_next_bbt_burstcount = ((((custom_dma_burst_4_upstream_write) && (custom_dma_burst_4_upstream_bbt_burstcounter == 0))))? (custom_dma_burst_4_upstream_burstcount - 1) :
    ((((custom_dma_burst_4_upstream_read) && (custom_dma_burst_4_upstream_bbt_burstcounter == 0))))? 0 :
    (custom_dma_burst_4_upstream_bbt_burstcounter - 1);

  //custom_dma_burst_4_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_upstream_bbt_burstcounter <= 0;
      else if (custom_dma_burst_4_upstream_begins_xfer)
          custom_dma_burst_4_upstream_bbt_burstcounter <= custom_dma_burst_4_upstream_next_bbt_burstcount;
    end


  //custom_dma_burst_4_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_4_upstream_beginbursttransfer_internal = custom_dma_burst_4_upstream_begins_xfer & (custom_dma_burst_4_upstream_bbt_burstcounter == 0);

  //custom_dma_burst_4_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_4_upstream_read = cpu_data_master_granted_custom_dma_burst_4_upstream & cpu_data_master_read;

  //custom_dma_burst_4_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_4_upstream_write = cpu_data_master_granted_custom_dma_burst_4_upstream & cpu_data_master_write;

  //custom_dma_burst_4_upstream_address mux, which is an e_mux
  assign custom_dma_burst_4_upstream_address = cpu_data_master_address_to_slave;

  //d1_custom_dma_burst_4_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_4_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_4_upstream_end_xfer <= custom_dma_burst_4_upstream_end_xfer;
    end


  //custom_dma_burst_4_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_4_upstream_waits_for_read = custom_dma_burst_4_upstream_in_a_read_cycle & custom_dma_burst_4_upstream_waitrequest_from_sa;

  //custom_dma_burst_4_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_4_upstream_in_a_read_cycle = cpu_data_master_granted_custom_dma_burst_4_upstream & cpu_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_4_upstream_in_a_read_cycle;

  //custom_dma_burst_4_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_4_upstream_waits_for_write = custom_dma_burst_4_upstream_in_a_write_cycle & custom_dma_burst_4_upstream_waitrequest_from_sa;

  //custom_dma_burst_4_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_4_upstream_in_a_write_cycle = cpu_data_master_granted_custom_dma_burst_4_upstream & cpu_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_4_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_4_upstream_counter = 0;
  //custom_dma_burst_4_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_4_upstream_byteenable = (cpu_data_master_granted_custom_dma_burst_4_upstream)? cpu_data_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign custom_dma_burst_4_upstream_burstcount = (cpu_data_master_granted_custom_dma_burst_4_upstream)? cpu_data_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_4_upstream_debugaccess = (cpu_data_master_granted_custom_dma_burst_4_upstream)? cpu_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_4/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //cpu/data_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_data_master_requests_custom_dma_burst_4_upstream && (cpu_data_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: cpu/data_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_4/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_4_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_4_downstream_address,
                                                   custom_dma_burst_4_downstream_burstcount,
                                                   custom_dma_burst_4_downstream_byteenable,
                                                   custom_dma_burst_4_downstream_granted_ddr_sdram_s1,
                                                   custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1,
                                                   custom_dma_burst_4_downstream_read,
                                                   custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1,
                                                   custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                                   custom_dma_burst_4_downstream_requests_ddr_sdram_s1,
                                                   custom_dma_burst_4_downstream_write,
                                                   custom_dma_burst_4_downstream_writedata,
                                                   d1_ddr_sdram_s1_end_xfer,
                                                   ddr_sdram_s1_readdata_from_sa,
                                                   ddr_sdram_s1_waitrequest_n_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_4_downstream_address_to_slave,
                                                   custom_dma_burst_4_downstream_latency_counter,
                                                   custom_dma_burst_4_downstream_readdata,
                                                   custom_dma_burst_4_downstream_readdatavalid,
                                                   custom_dma_burst_4_downstream_reset_n,
                                                   custom_dma_burst_4_downstream_waitrequest
                                                )
;

  output  [ 24: 0] custom_dma_burst_4_downstream_address_to_slave;
  output           custom_dma_burst_4_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_4_downstream_readdata;
  output           custom_dma_burst_4_downstream_readdatavalid;
  output           custom_dma_burst_4_downstream_reset_n;
  output           custom_dma_burst_4_downstream_waitrequest;
  input            clk;
  input   [ 24: 0] custom_dma_burst_4_downstream_address;
  input   [  2: 0] custom_dma_burst_4_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_4_downstream_byteenable;
  input            custom_dma_burst_4_downstream_granted_ddr_sdram_s1;
  input            custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1;
  input            custom_dma_burst_4_downstream_read;
  input            custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1;
  input            custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  input            custom_dma_burst_4_downstream_requests_ddr_sdram_s1;
  input            custom_dma_burst_4_downstream_write;
  input   [ 31: 0] custom_dma_burst_4_downstream_writedata;
  input            d1_ddr_sdram_s1_end_xfer;
  input   [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  input            ddr_sdram_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] custom_dma_burst_4_downstream_address_last_time;
  wire    [ 24: 0] custom_dma_burst_4_downstream_address_to_slave;
  reg     [  2: 0] custom_dma_burst_4_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_4_downstream_byteenable_last_time;
  wire             custom_dma_burst_4_downstream_is_granted_some_slave;
  reg              custom_dma_burst_4_downstream_latency_counter;
  reg              custom_dma_burst_4_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_4_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_4_downstream_readdata;
  wire             custom_dma_burst_4_downstream_readdatavalid;
  wire             custom_dma_burst_4_downstream_reset_n;
  wire             custom_dma_burst_4_downstream_run;
  wire             custom_dma_burst_4_downstream_waitrequest;
  reg              custom_dma_burst_4_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_4_downstream_writedata_last_time;
  wire             latency_load_value;
  wire             p1_custom_dma_burst_4_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_4_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1 | ~custom_dma_burst_4_downstream_requests_ddr_sdram_s1) & (custom_dma_burst_4_downstream_granted_ddr_sdram_s1 | ~custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1) & ((~custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write)))) & ((~custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_4_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_4_downstream_address_to_slave = custom_dma_burst_4_downstream_address;

  //custom_dma_burst_4_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_4_downstream_read_but_no_slave_selected <= custom_dma_burst_4_downstream_read & custom_dma_burst_4_downstream_run & ~custom_dma_burst_4_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_4_downstream_is_granted_some_slave = custom_dma_burst_4_downstream_granted_ddr_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_4_downstream_readdatavalid = custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_4_downstream_readdatavalid = custom_dma_burst_4_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_4_downstream_readdatavalid;

  //custom_dma_burst_4/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_4_downstream_readdata = ddr_sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_4_downstream_waitrequest = ~custom_dma_burst_4_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_4_downstream_latency_counter <= p1_custom_dma_burst_4_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_4_downstream_latency_counter = ((custom_dma_burst_4_downstream_run & custom_dma_burst_4_downstream_read))? latency_load_value :
    (custom_dma_burst_4_downstream_latency_counter)? custom_dma_burst_4_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //custom_dma_burst_4_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_4_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_4_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_address_last_time <= custom_dma_burst_4_downstream_address;
    end


  //custom_dma_burst_4/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_4_downstream_waitrequest & (custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write);
    end


  //custom_dma_burst_4_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_address != custom_dma_burst_4_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_4_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_burstcount_last_time <= custom_dma_burst_4_downstream_burstcount;
    end


  //custom_dma_burst_4_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_burstcount != custom_dma_burst_4_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_4_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_byteenable_last_time <= custom_dma_burst_4_downstream_byteenable;
    end


  //custom_dma_burst_4_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_byteenable != custom_dma_burst_4_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_4_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_read_last_time <= custom_dma_burst_4_downstream_read;
    end


  //custom_dma_burst_4_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_read != custom_dma_burst_4_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_4_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_write_last_time <= custom_dma_burst_4_downstream_write;
    end


  //custom_dma_burst_4_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_write != custom_dma_burst_4_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_4_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_4_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_4_downstream_writedata_last_time <= custom_dma_burst_4_downstream_writedata;
    end


  //custom_dma_burst_4_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_4_downstream_writedata != custom_dma_burst_4_downstream_writedata_last_time) & custom_dma_burst_4_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_4_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_5_upstream_arbitrator (
                                                // inputs:
                                                 clk,
                                                 custom_dma_burst_5_upstream_readdata,
                                                 custom_dma_burst_5_upstream_readdatavalid,
                                                 custom_dma_burst_5_upstream_waitrequest,
                                                 fir_dma_write_master_address_to_slave,
                                                 fir_dma_write_master_burstcount,
                                                 fir_dma_write_master_byteenable,
                                                 fir_dma_write_master_write,
                                                 fir_dma_write_master_writedata,
                                                 reset_n,

                                                // outputs:
                                                 custom_dma_burst_5_upstream_address,
                                                 custom_dma_burst_5_upstream_burstcount,
                                                 custom_dma_burst_5_upstream_byteaddress,
                                                 custom_dma_burst_5_upstream_byteenable,
                                                 custom_dma_burst_5_upstream_debugaccess,
                                                 custom_dma_burst_5_upstream_read,
                                                 custom_dma_burst_5_upstream_readdata_from_sa,
                                                 custom_dma_burst_5_upstream_readdatavalid_from_sa,
                                                 custom_dma_burst_5_upstream_waitrequest_from_sa,
                                                 custom_dma_burst_5_upstream_write,
                                                 custom_dma_burst_5_upstream_writedata,
                                                 d1_custom_dma_burst_5_upstream_end_xfer,
                                                 fir_dma_write_master_granted_custom_dma_burst_5_upstream,
                                                 fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream,
                                                 fir_dma_write_master_requests_custom_dma_burst_5_upstream
                                              )
;

  output  [ 24: 0] custom_dma_burst_5_upstream_address;
  output  [  2: 0] custom_dma_burst_5_upstream_burstcount;
  output  [ 26: 0] custom_dma_burst_5_upstream_byteaddress;
  output  [  3: 0] custom_dma_burst_5_upstream_byteenable;
  output           custom_dma_burst_5_upstream_debugaccess;
  output           custom_dma_burst_5_upstream_read;
  output  [ 31: 0] custom_dma_burst_5_upstream_readdata_from_sa;
  output           custom_dma_burst_5_upstream_readdatavalid_from_sa;
  output           custom_dma_burst_5_upstream_waitrequest_from_sa;
  output           custom_dma_burst_5_upstream_write;
  output  [ 31: 0] custom_dma_burst_5_upstream_writedata;
  output           d1_custom_dma_burst_5_upstream_end_xfer;
  output           fir_dma_write_master_granted_custom_dma_burst_5_upstream;
  output           fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream;
  output           fir_dma_write_master_requests_custom_dma_burst_5_upstream;
  input            clk;
  input   [ 31: 0] custom_dma_burst_5_upstream_readdata;
  input            custom_dma_burst_5_upstream_readdatavalid;
  input            custom_dma_burst_5_upstream_waitrequest;
  input   [ 31: 0] fir_dma_write_master_address_to_slave;
  input   [  2: 0] fir_dma_write_master_burstcount;
  input   [  3: 0] fir_dma_write_master_byteenable;
  input            fir_dma_write_master_write;
  input   [ 31: 0] fir_dma_write_master_writedata;
  input            reset_n;

  wire    [ 24: 0] custom_dma_burst_5_upstream_address;
  wire             custom_dma_burst_5_upstream_allgrants;
  wire             custom_dma_burst_5_upstream_allow_new_arb_cycle;
  wire             custom_dma_burst_5_upstream_any_bursting_master_saved_grant;
  wire             custom_dma_burst_5_upstream_any_continuerequest;
  wire             custom_dma_burst_5_upstream_arb_counter_enable;
  reg     [  2: 0] custom_dma_burst_5_upstream_arb_share_counter;
  wire    [  2: 0] custom_dma_burst_5_upstream_arb_share_counter_next_value;
  wire    [  2: 0] custom_dma_burst_5_upstream_arb_share_set_values;
  reg     [  1: 0] custom_dma_burst_5_upstream_bbt_burstcounter;
  wire             custom_dma_burst_5_upstream_beginbursttransfer_internal;
  wire             custom_dma_burst_5_upstream_begins_xfer;
  wire    [  2: 0] custom_dma_burst_5_upstream_burstcount;
  wire    [ 26: 0] custom_dma_burst_5_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_5_upstream_byteenable;
  wire             custom_dma_burst_5_upstream_debugaccess;
  wire             custom_dma_burst_5_upstream_end_xfer;
  wire             custom_dma_burst_5_upstream_firsttransfer;
  wire             custom_dma_burst_5_upstream_grant_vector;
  wire             custom_dma_burst_5_upstream_in_a_read_cycle;
  wire             custom_dma_burst_5_upstream_in_a_write_cycle;
  wire             custom_dma_burst_5_upstream_master_qreq_vector;
  wire    [  1: 0] custom_dma_burst_5_upstream_next_bbt_burstcount;
  wire             custom_dma_burst_5_upstream_non_bursting_master_requests;
  wire             custom_dma_burst_5_upstream_read;
  wire    [ 31: 0] custom_dma_burst_5_upstream_readdata_from_sa;
  wire             custom_dma_burst_5_upstream_readdatavalid_from_sa;
  reg              custom_dma_burst_5_upstream_reg_firsttransfer;
  reg              custom_dma_burst_5_upstream_slavearbiterlockenable;
  wire             custom_dma_burst_5_upstream_slavearbiterlockenable2;
  wire             custom_dma_burst_5_upstream_unreg_firsttransfer;
  wire             custom_dma_burst_5_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_5_upstream_waits_for_read;
  wire             custom_dma_burst_5_upstream_waits_for_write;
  wire             custom_dma_burst_5_upstream_write;
  wire    [ 31: 0] custom_dma_burst_5_upstream_writedata;
  reg              d1_custom_dma_burst_5_upstream_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_arbiterlock;
  wire             fir_dma_write_master_arbiterlock2;
  wire             fir_dma_write_master_continuerequest;
  wire             fir_dma_write_master_granted_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_requests_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_saved_grant_custom_dma_burst_5_upstream;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             wait_for_custom_dma_burst_5_upstream_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_burst_5_upstream_end_xfer;
    end


  assign custom_dma_burst_5_upstream_begins_xfer = ~d1_reasons_to_wait & ((fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream));
  //assign custom_dma_burst_5_upstream_readdata_from_sa = custom_dma_burst_5_upstream_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_5_upstream_readdata_from_sa = custom_dma_burst_5_upstream_readdata;

  assign fir_dma_write_master_requests_custom_dma_burst_5_upstream = (({fir_dma_write_master_address_to_slave[31 : 25] , 25'b0} == 32'h2000000) & (fir_dma_write_master_write)) & fir_dma_write_master_write;
  //assign custom_dma_burst_5_upstream_waitrequest_from_sa = custom_dma_burst_5_upstream_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_5_upstream_waitrequest_from_sa = custom_dma_burst_5_upstream_waitrequest;

  //custom_dma_burst_5_upstream_arb_share_counter set values, which is an e_mux
  assign custom_dma_burst_5_upstream_arb_share_set_values = (fir_dma_write_master_granted_custom_dma_burst_5_upstream)? fir_dma_write_master_burstcount :
    1;

  //custom_dma_burst_5_upstream_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_burst_5_upstream_non_bursting_master_requests = 0;

  //custom_dma_burst_5_upstream_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_burst_5_upstream_any_bursting_master_saved_grant = fir_dma_write_master_saved_grant_custom_dma_burst_5_upstream;

  //custom_dma_burst_5_upstream_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_burst_5_upstream_arb_share_counter_next_value = custom_dma_burst_5_upstream_firsttransfer ? (custom_dma_burst_5_upstream_arb_share_set_values - 1) : |custom_dma_burst_5_upstream_arb_share_counter ? (custom_dma_burst_5_upstream_arb_share_counter - 1) : 0;

  //custom_dma_burst_5_upstream_allgrants all slave grants, which is an e_mux
  assign custom_dma_burst_5_upstream_allgrants = |custom_dma_burst_5_upstream_grant_vector;

  //custom_dma_burst_5_upstream_end_xfer assignment, which is an e_assign
  assign custom_dma_burst_5_upstream_end_xfer = ~(custom_dma_burst_5_upstream_waits_for_read | custom_dma_burst_5_upstream_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream = custom_dma_burst_5_upstream_end_xfer & (~custom_dma_burst_5_upstream_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_burst_5_upstream_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_burst_5_upstream_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream & custom_dma_burst_5_upstream_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream & ~custom_dma_burst_5_upstream_non_bursting_master_requests);

  //custom_dma_burst_5_upstream_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_upstream_arb_share_counter <= 0;
      else if (custom_dma_burst_5_upstream_arb_counter_enable)
          custom_dma_burst_5_upstream_arb_share_counter <= custom_dma_burst_5_upstream_arb_share_counter_next_value;
    end


  //custom_dma_burst_5_upstream_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_upstream_slavearbiterlockenable <= 0;
      else if ((|custom_dma_burst_5_upstream_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream) | (end_xfer_arb_share_counter_term_custom_dma_burst_5_upstream & ~custom_dma_burst_5_upstream_non_bursting_master_requests))
          custom_dma_burst_5_upstream_slavearbiterlockenable <= |custom_dma_burst_5_upstream_arb_share_counter_next_value;
    end


  //fir_dma/write_master custom_dma_burst_5/upstream arbiterlock, which is an e_assign
  assign fir_dma_write_master_arbiterlock = custom_dma_burst_5_upstream_slavearbiterlockenable & fir_dma_write_master_continuerequest;

  //custom_dma_burst_5_upstream_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_burst_5_upstream_slavearbiterlockenable2 = |custom_dma_burst_5_upstream_arb_share_counter_next_value;

  //fir_dma/write_master custom_dma_burst_5/upstream arbiterlock2, which is an e_assign
  assign fir_dma_write_master_arbiterlock2 = custom_dma_burst_5_upstream_slavearbiterlockenable2 & fir_dma_write_master_continuerequest;

  //custom_dma_burst_5_upstream_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_burst_5_upstream_any_continuerequest = 1;

  //fir_dma_write_master_continuerequest continued request, which is an e_assign
  assign fir_dma_write_master_continuerequest = 1;

  assign fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream = fir_dma_write_master_requests_custom_dma_burst_5_upstream;
  //custom_dma_burst_5_upstream_writedata mux, which is an e_mux
  assign custom_dma_burst_5_upstream_writedata = fir_dma_write_master_writedata;

  //byteaddress mux for custom_dma_burst_5/upstream, which is an e_mux
  assign custom_dma_burst_5_upstream_byteaddress = fir_dma_write_master_address_to_slave;

  //master is always granted when requested
  assign fir_dma_write_master_granted_custom_dma_burst_5_upstream = fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream;

  //fir_dma/write_master saved-grant custom_dma_burst_5/upstream, which is an e_assign
  assign fir_dma_write_master_saved_grant_custom_dma_burst_5_upstream = fir_dma_write_master_requests_custom_dma_burst_5_upstream;

  //allow new arb cycle for custom_dma_burst_5/upstream, which is an e_assign
  assign custom_dma_burst_5_upstream_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_burst_5_upstream_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_burst_5_upstream_master_qreq_vector = 1;

  //custom_dma_burst_5_upstream_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_5_upstream_firsttransfer = custom_dma_burst_5_upstream_begins_xfer ? custom_dma_burst_5_upstream_unreg_firsttransfer : custom_dma_burst_5_upstream_reg_firsttransfer;

  //custom_dma_burst_5_upstream_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_burst_5_upstream_unreg_firsttransfer = ~(custom_dma_burst_5_upstream_slavearbiterlockenable & custom_dma_burst_5_upstream_any_continuerequest);

  //custom_dma_burst_5_upstream_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_upstream_reg_firsttransfer <= 1'b1;
      else if (custom_dma_burst_5_upstream_begins_xfer)
          custom_dma_burst_5_upstream_reg_firsttransfer <= custom_dma_burst_5_upstream_unreg_firsttransfer;
    end


  //custom_dma_burst_5_upstream_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign custom_dma_burst_5_upstream_next_bbt_burstcount = ((((custom_dma_burst_5_upstream_write) && (custom_dma_burst_5_upstream_bbt_burstcounter == 0))))? (custom_dma_burst_5_upstream_burstcount - 1) :
    ((((custom_dma_burst_5_upstream_read) && (custom_dma_burst_5_upstream_bbt_burstcounter == 0))))? 0 :
    (custom_dma_burst_5_upstream_bbt_burstcounter - 1);

  //custom_dma_burst_5_upstream_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_upstream_bbt_burstcounter <= 0;
      else if (custom_dma_burst_5_upstream_begins_xfer)
          custom_dma_burst_5_upstream_bbt_burstcounter <= custom_dma_burst_5_upstream_next_bbt_burstcount;
    end


  //custom_dma_burst_5_upstream_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_burst_5_upstream_beginbursttransfer_internal = custom_dma_burst_5_upstream_begins_xfer & (custom_dma_burst_5_upstream_bbt_burstcounter == 0);

  //custom_dma_burst_5_upstream_read assignment, which is an e_mux
  assign custom_dma_burst_5_upstream_read = 0;

  //custom_dma_burst_5_upstream_write assignment, which is an e_mux
  assign custom_dma_burst_5_upstream_write = fir_dma_write_master_granted_custom_dma_burst_5_upstream & fir_dma_write_master_write;

  //custom_dma_burst_5_upstream_address mux, which is an e_mux
  assign custom_dma_burst_5_upstream_address = fir_dma_write_master_address_to_slave;

  //d1_custom_dma_burst_5_upstream_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_burst_5_upstream_end_xfer <= 1;
      else 
        d1_custom_dma_burst_5_upstream_end_xfer <= custom_dma_burst_5_upstream_end_xfer;
    end


  //custom_dma_burst_5_upstream_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_burst_5_upstream_waits_for_read = custom_dma_burst_5_upstream_in_a_read_cycle & custom_dma_burst_5_upstream_waitrequest_from_sa;

  //custom_dma_burst_5_upstream_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_burst_5_upstream_in_a_read_cycle = 0;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_burst_5_upstream_in_a_read_cycle;

  //custom_dma_burst_5_upstream_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_burst_5_upstream_waits_for_write = custom_dma_burst_5_upstream_in_a_write_cycle & custom_dma_burst_5_upstream_waitrequest_from_sa;

  //assign custom_dma_burst_5_upstream_readdatavalid_from_sa = custom_dma_burst_5_upstream_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_burst_5_upstream_readdatavalid_from_sa = custom_dma_burst_5_upstream_readdatavalid;

  //custom_dma_burst_5_upstream_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_burst_5_upstream_in_a_write_cycle = fir_dma_write_master_granted_custom_dma_burst_5_upstream & fir_dma_write_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_burst_5_upstream_in_a_write_cycle;

  assign wait_for_custom_dma_burst_5_upstream_counter = 0;
  //custom_dma_burst_5_upstream_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_burst_5_upstream_byteenable = (fir_dma_write_master_granted_custom_dma_burst_5_upstream)? fir_dma_write_master_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign custom_dma_burst_5_upstream_burstcount = (fir_dma_write_master_granted_custom_dma_burst_5_upstream)? fir_dma_write_master_burstcount :
    1;

  //debugaccess mux, which is an e_mux
  assign custom_dma_burst_5_upstream_debugaccess = 0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_5/upstream enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //fir_dma/write_master non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (fir_dma_write_master_requests_custom_dma_burst_5_upstream && (fir_dma_write_master_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: fir_dma/write_master drove 0 on its 'burstcount' port while accessing slave custom_dma_burst_5/upstream", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_burst_5_downstream_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   custom_dma_burst_5_downstream_address,
                                                   custom_dma_burst_5_downstream_burstcount,
                                                   custom_dma_burst_5_downstream_byteenable,
                                                   custom_dma_burst_5_downstream_granted_ddr_sdram_s1,
                                                   custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1,
                                                   custom_dma_burst_5_downstream_read,
                                                   custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1,
                                                   custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                                   custom_dma_burst_5_downstream_requests_ddr_sdram_s1,
                                                   custom_dma_burst_5_downstream_write,
                                                   custom_dma_burst_5_downstream_writedata,
                                                   d1_ddr_sdram_s1_end_xfer,
                                                   ddr_sdram_s1_readdata_from_sa,
                                                   ddr_sdram_s1_waitrequest_n_from_sa,
                                                   reset_n,

                                                  // outputs:
                                                   custom_dma_burst_5_downstream_address_to_slave,
                                                   custom_dma_burst_5_downstream_latency_counter,
                                                   custom_dma_burst_5_downstream_readdata,
                                                   custom_dma_burst_5_downstream_readdatavalid,
                                                   custom_dma_burst_5_downstream_reset_n,
                                                   custom_dma_burst_5_downstream_waitrequest
                                                )
;

  output  [ 24: 0] custom_dma_burst_5_downstream_address_to_slave;
  output           custom_dma_burst_5_downstream_latency_counter;
  output  [ 31: 0] custom_dma_burst_5_downstream_readdata;
  output           custom_dma_burst_5_downstream_readdatavalid;
  output           custom_dma_burst_5_downstream_reset_n;
  output           custom_dma_burst_5_downstream_waitrequest;
  input            clk;
  input   [ 24: 0] custom_dma_burst_5_downstream_address;
  input   [  2: 0] custom_dma_burst_5_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_5_downstream_byteenable;
  input            custom_dma_burst_5_downstream_granted_ddr_sdram_s1;
  input            custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1;
  input            custom_dma_burst_5_downstream_read;
  input            custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1;
  input            custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  input            custom_dma_burst_5_downstream_requests_ddr_sdram_s1;
  input            custom_dma_burst_5_downstream_write;
  input   [ 31: 0] custom_dma_burst_5_downstream_writedata;
  input            d1_ddr_sdram_s1_end_xfer;
  input   [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  input            ddr_sdram_s1_waitrequest_n_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] custom_dma_burst_5_downstream_address_last_time;
  wire    [ 24: 0] custom_dma_burst_5_downstream_address_to_slave;
  reg     [  2: 0] custom_dma_burst_5_downstream_burstcount_last_time;
  reg     [  3: 0] custom_dma_burst_5_downstream_byteenable_last_time;
  wire             custom_dma_burst_5_downstream_is_granted_some_slave;
  reg              custom_dma_burst_5_downstream_latency_counter;
  reg              custom_dma_burst_5_downstream_read_but_no_slave_selected;
  reg              custom_dma_burst_5_downstream_read_last_time;
  wire    [ 31: 0] custom_dma_burst_5_downstream_readdata;
  wire             custom_dma_burst_5_downstream_readdatavalid;
  wire             custom_dma_burst_5_downstream_reset_n;
  wire             custom_dma_burst_5_downstream_run;
  wire             custom_dma_burst_5_downstream_waitrequest;
  reg              custom_dma_burst_5_downstream_write_last_time;
  reg     [ 31: 0] custom_dma_burst_5_downstream_writedata_last_time;
  wire             latency_load_value;
  wire             p1_custom_dma_burst_5_downstream_latency_counter;
  wire             pre_flush_custom_dma_burst_5_downstream_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1 | ~custom_dma_burst_5_downstream_requests_ddr_sdram_s1) & (custom_dma_burst_5_downstream_granted_ddr_sdram_s1 | ~custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1) & ((~custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write)))) & ((~custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1 | ~(custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write) | (1 & ddr_sdram_s1_waitrequest_n_from_sa & (custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write))));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_burst_5_downstream_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_burst_5_downstream_address_to_slave = custom_dma_burst_5_downstream_address;

  //custom_dma_burst_5_downstream_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_read_but_no_slave_selected <= 0;
      else 
        custom_dma_burst_5_downstream_read_but_no_slave_selected <= custom_dma_burst_5_downstream_read & custom_dma_burst_5_downstream_run & ~custom_dma_burst_5_downstream_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign custom_dma_burst_5_downstream_is_granted_some_slave = custom_dma_burst_5_downstream_granted_ddr_sdram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_custom_dma_burst_5_downstream_readdatavalid = custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign custom_dma_burst_5_downstream_readdatavalid = custom_dma_burst_5_downstream_read_but_no_slave_selected |
    pre_flush_custom_dma_burst_5_downstream_readdatavalid;

  //custom_dma_burst_5/downstream readdata mux, which is an e_mux
  assign custom_dma_burst_5_downstream_readdata = ddr_sdram_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_burst_5_downstream_waitrequest = ~custom_dma_burst_5_downstream_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_latency_counter <= 0;
      else 
        custom_dma_burst_5_downstream_latency_counter <= p1_custom_dma_burst_5_downstream_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_custom_dma_burst_5_downstream_latency_counter = ((custom_dma_burst_5_downstream_run & custom_dma_burst_5_downstream_read))? latency_load_value :
    (custom_dma_burst_5_downstream_latency_counter)? custom_dma_burst_5_downstream_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = 0;

  //custom_dma_burst_5_downstream_reset_n assignment, which is an e_assign
  assign custom_dma_burst_5_downstream_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_burst_5_downstream_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_address_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_address_last_time <= custom_dma_burst_5_downstream_address;
    end


  //custom_dma_burst_5/downstream waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_burst_5_downstream_waitrequest & (custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write);
    end


  //custom_dma_burst_5_downstream_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_address != custom_dma_burst_5_downstream_address_last_time))
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_5_downstream_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_burstcount_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_burstcount_last_time <= custom_dma_burst_5_downstream_burstcount;
    end


  //custom_dma_burst_5_downstream_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_burstcount != custom_dma_burst_5_downstream_burstcount_last_time))
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_5_downstream_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_byteenable_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_byteenable_last_time <= custom_dma_burst_5_downstream_byteenable;
    end


  //custom_dma_burst_5_downstream_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_byteenable != custom_dma_burst_5_downstream_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_5_downstream_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_read_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_read_last_time <= custom_dma_burst_5_downstream_read;
    end


  //custom_dma_burst_5_downstream_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_read != custom_dma_burst_5_downstream_read_last_time))
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_5_downstream_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_write_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_write_last_time <= custom_dma_burst_5_downstream_write;
    end


  //custom_dma_burst_5_downstream_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_write != custom_dma_burst_5_downstream_write_last_time))
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_burst_5_downstream_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_5_downstream_writedata_last_time <= 0;
      else 
        custom_dma_burst_5_downstream_writedata_last_time <= custom_dma_burst_5_downstream_writedata;
    end


  //custom_dma_burst_5_downstream_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_burst_5_downstream_writedata != custom_dma_burst_5_downstream_writedata_last_time) & custom_dma_burst_5_downstream_write)
        begin
          $write("%0d ns: custom_dma_burst_5_downstream_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_in_arbitrator (
                                          // inputs:
                                           clk,
                                           custom_dma_clock_0_in_endofpacket,
                                           custom_dma_clock_0_in_readdata,
                                           custom_dma_clock_0_in_waitrequest,
                                           pipeline_bridge_m1_address_to_slave,
                                           pipeline_bridge_m1_burstcount,
                                           pipeline_bridge_m1_byteenable,
                                           pipeline_bridge_m1_chipselect,
                                           pipeline_bridge_m1_latency_counter,
                                           pipeline_bridge_m1_read,
                                           pipeline_bridge_m1_write,
                                           pipeline_bridge_m1_writedata,
                                           reset_n,

                                          // outputs:
                                           custom_dma_clock_0_in_address,
                                           custom_dma_clock_0_in_byteenable,
                                           custom_dma_clock_0_in_endofpacket_from_sa,
                                           custom_dma_clock_0_in_nativeaddress,
                                           custom_dma_clock_0_in_read,
                                           custom_dma_clock_0_in_readdata_from_sa,
                                           custom_dma_clock_0_in_reset_n,
                                           custom_dma_clock_0_in_waitrequest_from_sa,
                                           custom_dma_clock_0_in_write,
                                           custom_dma_clock_0_in_writedata,
                                           d1_custom_dma_clock_0_in_end_xfer,
                                           pipeline_bridge_m1_granted_custom_dma_clock_0_in,
                                           pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in,
                                           pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in,
                                           pipeline_bridge_m1_requests_custom_dma_clock_0_in
                                        )
;

  output  [  3: 0] custom_dma_clock_0_in_address;
  output  [  1: 0] custom_dma_clock_0_in_byteenable;
  output           custom_dma_clock_0_in_endofpacket_from_sa;
  output  [  2: 0] custom_dma_clock_0_in_nativeaddress;
  output           custom_dma_clock_0_in_read;
  output  [ 15: 0] custom_dma_clock_0_in_readdata_from_sa;
  output           custom_dma_clock_0_in_reset_n;
  output           custom_dma_clock_0_in_waitrequest_from_sa;
  output           custom_dma_clock_0_in_write;
  output  [ 15: 0] custom_dma_clock_0_in_writedata;
  output           d1_custom_dma_clock_0_in_end_xfer;
  output           pipeline_bridge_m1_granted_custom_dma_clock_0_in;
  output           pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in;
  output           pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in;
  output           pipeline_bridge_m1_requests_custom_dma_clock_0_in;
  input            clk;
  input            custom_dma_clock_0_in_endofpacket;
  input   [ 15: 0] custom_dma_clock_0_in_readdata;
  input            custom_dma_clock_0_in_waitrequest;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  wire    [  3: 0] custom_dma_clock_0_in_address;
  wire             custom_dma_clock_0_in_allgrants;
  wire             custom_dma_clock_0_in_allow_new_arb_cycle;
  wire             custom_dma_clock_0_in_any_bursting_master_saved_grant;
  wire             custom_dma_clock_0_in_any_continuerequest;
  wire             custom_dma_clock_0_in_arb_counter_enable;
  reg              custom_dma_clock_0_in_arb_share_counter;
  wire             custom_dma_clock_0_in_arb_share_counter_next_value;
  wire             custom_dma_clock_0_in_arb_share_set_values;
  wire             custom_dma_clock_0_in_beginbursttransfer_internal;
  wire             custom_dma_clock_0_in_begins_xfer;
  wire    [  1: 0] custom_dma_clock_0_in_byteenable;
  wire             custom_dma_clock_0_in_end_xfer;
  wire             custom_dma_clock_0_in_endofpacket_from_sa;
  wire             custom_dma_clock_0_in_firsttransfer;
  wire             custom_dma_clock_0_in_grant_vector;
  wire             custom_dma_clock_0_in_in_a_read_cycle;
  wire             custom_dma_clock_0_in_in_a_write_cycle;
  wire             custom_dma_clock_0_in_master_qreq_vector;
  wire    [  2: 0] custom_dma_clock_0_in_nativeaddress;
  wire             custom_dma_clock_0_in_non_bursting_master_requests;
  wire             custom_dma_clock_0_in_read;
  wire    [ 15: 0] custom_dma_clock_0_in_readdata_from_sa;
  reg              custom_dma_clock_0_in_reg_firsttransfer;
  wire             custom_dma_clock_0_in_reset_n;
  reg              custom_dma_clock_0_in_slavearbiterlockenable;
  wire             custom_dma_clock_0_in_slavearbiterlockenable2;
  wire             custom_dma_clock_0_in_unreg_firsttransfer;
  wire             custom_dma_clock_0_in_waitrequest_from_sa;
  wire             custom_dma_clock_0_in_waits_for_read;
  wire             custom_dma_clock_0_in_waits_for_write;
  wire             custom_dma_clock_0_in_write;
  wire    [ 15: 0] custom_dma_clock_0_in_writedata;
  reg              d1_custom_dma_clock_0_in_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_custom_dma_clock_0_in;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_requests_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_saved_grant_custom_dma_clock_0_in;
  wire    [ 11: 0] shifted_address_to_custom_dma_clock_0_in_from_pipeline_bridge_m1;
  wire             wait_for_custom_dma_clock_0_in_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~custom_dma_clock_0_in_end_xfer;
    end


  assign custom_dma_clock_0_in_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in));
  //assign custom_dma_clock_0_in_readdata_from_sa = custom_dma_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_clock_0_in_readdata_from_sa = custom_dma_clock_0_in_readdata;

  assign pipeline_bridge_m1_requests_custom_dma_clock_0_in = ({pipeline_bridge_m1_address_to_slave[11 : 5] , 5'b0} == 12'h820) & pipeline_bridge_m1_chipselect;
  //assign custom_dma_clock_0_in_waitrequest_from_sa = custom_dma_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_clock_0_in_waitrequest_from_sa = custom_dma_clock_0_in_waitrequest;

  //custom_dma_clock_0_in_arb_share_counter set values, which is an e_mux
  assign custom_dma_clock_0_in_arb_share_set_values = 1;

  //custom_dma_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  assign custom_dma_clock_0_in_non_bursting_master_requests = pipeline_bridge_m1_requests_custom_dma_clock_0_in;

  //custom_dma_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  assign custom_dma_clock_0_in_any_bursting_master_saved_grant = 0;

  //custom_dma_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  assign custom_dma_clock_0_in_arb_share_counter_next_value = custom_dma_clock_0_in_firsttransfer ? (custom_dma_clock_0_in_arb_share_set_values - 1) : |custom_dma_clock_0_in_arb_share_counter ? (custom_dma_clock_0_in_arb_share_counter - 1) : 0;

  //custom_dma_clock_0_in_allgrants all slave grants, which is an e_mux
  assign custom_dma_clock_0_in_allgrants = |custom_dma_clock_0_in_grant_vector;

  //custom_dma_clock_0_in_end_xfer assignment, which is an e_assign
  assign custom_dma_clock_0_in_end_xfer = ~(custom_dma_clock_0_in_waits_for_read | custom_dma_clock_0_in_waits_for_write);

  //end_xfer_arb_share_counter_term_custom_dma_clock_0_in arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_custom_dma_clock_0_in = custom_dma_clock_0_in_end_xfer & (~custom_dma_clock_0_in_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //custom_dma_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  assign custom_dma_clock_0_in_arb_counter_enable = (end_xfer_arb_share_counter_term_custom_dma_clock_0_in & custom_dma_clock_0_in_allgrants) | (end_xfer_arb_share_counter_term_custom_dma_clock_0_in & ~custom_dma_clock_0_in_non_bursting_master_requests);

  //custom_dma_clock_0_in_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_in_arb_share_counter <= 0;
      else if (custom_dma_clock_0_in_arb_counter_enable)
          custom_dma_clock_0_in_arb_share_counter <= custom_dma_clock_0_in_arb_share_counter_next_value;
    end


  //custom_dma_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_in_slavearbiterlockenable <= 0;
      else if ((|custom_dma_clock_0_in_master_qreq_vector & end_xfer_arb_share_counter_term_custom_dma_clock_0_in) | (end_xfer_arb_share_counter_term_custom_dma_clock_0_in & ~custom_dma_clock_0_in_non_bursting_master_requests))
          custom_dma_clock_0_in_slavearbiterlockenable <= |custom_dma_clock_0_in_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 custom_dma_clock_0/in arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = custom_dma_clock_0_in_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //custom_dma_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign custom_dma_clock_0_in_slavearbiterlockenable2 = |custom_dma_clock_0_in_arb_share_counter_next_value;

  //pipeline_bridge/m1 custom_dma_clock_0/in arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = custom_dma_clock_0_in_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //custom_dma_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  assign custom_dma_clock_0_in_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in = pipeline_bridge_m1_requests_custom_dma_clock_0_in & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in = pipeline_bridge_m1_granted_custom_dma_clock_0_in & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~custom_dma_clock_0_in_waits_for_read;

  //custom_dma_clock_0_in_writedata mux, which is an e_mux
  assign custom_dma_clock_0_in_writedata = pipeline_bridge_m1_writedata;

  //assign custom_dma_clock_0_in_endofpacket_from_sa = custom_dma_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign custom_dma_clock_0_in_endofpacket_from_sa = custom_dma_clock_0_in_endofpacket;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_custom_dma_clock_0_in = pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in;

  //pipeline_bridge/m1 saved-grant custom_dma_clock_0/in, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_custom_dma_clock_0_in = pipeline_bridge_m1_requests_custom_dma_clock_0_in;

  //allow new arb cycle for custom_dma_clock_0/in, which is an e_assign
  assign custom_dma_clock_0_in_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign custom_dma_clock_0_in_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign custom_dma_clock_0_in_master_qreq_vector = 1;

  //custom_dma_clock_0_in_reset_n assignment, which is an e_assign
  assign custom_dma_clock_0_in_reset_n = reset_n;

  //custom_dma_clock_0_in_firsttransfer first transaction, which is an e_assign
  assign custom_dma_clock_0_in_firsttransfer = custom_dma_clock_0_in_begins_xfer ? custom_dma_clock_0_in_unreg_firsttransfer : custom_dma_clock_0_in_reg_firsttransfer;

  //custom_dma_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  assign custom_dma_clock_0_in_unreg_firsttransfer = ~(custom_dma_clock_0_in_slavearbiterlockenable & custom_dma_clock_0_in_any_continuerequest);

  //custom_dma_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_in_reg_firsttransfer <= 1'b1;
      else if (custom_dma_clock_0_in_begins_xfer)
          custom_dma_clock_0_in_reg_firsttransfer <= custom_dma_clock_0_in_unreg_firsttransfer;
    end


  //custom_dma_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign custom_dma_clock_0_in_beginbursttransfer_internal = custom_dma_clock_0_in_begins_xfer;

  //custom_dma_clock_0_in_read assignment, which is an e_mux
  assign custom_dma_clock_0_in_read = pipeline_bridge_m1_granted_custom_dma_clock_0_in & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //custom_dma_clock_0_in_write assignment, which is an e_mux
  assign custom_dma_clock_0_in_write = pipeline_bridge_m1_granted_custom_dma_clock_0_in & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_custom_dma_clock_0_in_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //custom_dma_clock_0_in_address mux, which is an e_mux
  assign custom_dma_clock_0_in_address = shifted_address_to_custom_dma_clock_0_in_from_pipeline_bridge_m1 >> 2;

  //slaveid custom_dma_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  assign custom_dma_clock_0_in_nativeaddress = pipeline_bridge_m1_address_to_slave >> 2;

  //d1_custom_dma_clock_0_in_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_custom_dma_clock_0_in_end_xfer <= 1;
      else 
        d1_custom_dma_clock_0_in_end_xfer <= custom_dma_clock_0_in_end_xfer;
    end


  //custom_dma_clock_0_in_waits_for_read in a cycle, which is an e_mux
  assign custom_dma_clock_0_in_waits_for_read = custom_dma_clock_0_in_in_a_read_cycle & custom_dma_clock_0_in_waitrequest_from_sa;

  //custom_dma_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  assign custom_dma_clock_0_in_in_a_read_cycle = pipeline_bridge_m1_granted_custom_dma_clock_0_in & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = custom_dma_clock_0_in_in_a_read_cycle;

  //custom_dma_clock_0_in_waits_for_write in a cycle, which is an e_mux
  assign custom_dma_clock_0_in_waits_for_write = custom_dma_clock_0_in_in_a_write_cycle & custom_dma_clock_0_in_waitrequest_from_sa;

  //custom_dma_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  assign custom_dma_clock_0_in_in_a_write_cycle = pipeline_bridge_m1_granted_custom_dma_clock_0_in & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = custom_dma_clock_0_in_in_a_write_cycle;

  assign wait_for_custom_dma_clock_0_in_counter = 0;
  //custom_dma_clock_0_in_byteenable byte enable port mux, which is an e_mux
  assign custom_dma_clock_0_in_byteenable = (pipeline_bridge_m1_granted_custom_dma_clock_0_in)? pipeline_bridge_m1_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_clock_0/in enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_custom_dma_clock_0_in && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave custom_dma_clock_0/in", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_out_arbitrator (
                                           // inputs:
                                            clk,
                                            custom_dma_clock_0_out_address,
                                            custom_dma_clock_0_out_byteenable,
                                            custom_dma_clock_0_out_granted_pll_s1,
                                            custom_dma_clock_0_out_qualified_request_pll_s1,
                                            custom_dma_clock_0_out_read,
                                            custom_dma_clock_0_out_read_data_valid_pll_s1,
                                            custom_dma_clock_0_out_requests_pll_s1,
                                            custom_dma_clock_0_out_write,
                                            custom_dma_clock_0_out_writedata,
                                            d1_pll_s1_end_xfer,
                                            pll_s1_readdata_from_sa,
                                            reset_n,

                                           // outputs:
                                            custom_dma_clock_0_out_address_to_slave,
                                            custom_dma_clock_0_out_readdata,
                                            custom_dma_clock_0_out_reset_n,
                                            custom_dma_clock_0_out_waitrequest
                                         )
;

  output  [  3: 0] custom_dma_clock_0_out_address_to_slave;
  output  [ 15: 0] custom_dma_clock_0_out_readdata;
  output           custom_dma_clock_0_out_reset_n;
  output           custom_dma_clock_0_out_waitrequest;
  input            clk;
  input   [  3: 0] custom_dma_clock_0_out_address;
  input   [  1: 0] custom_dma_clock_0_out_byteenable;
  input            custom_dma_clock_0_out_granted_pll_s1;
  input            custom_dma_clock_0_out_qualified_request_pll_s1;
  input            custom_dma_clock_0_out_read;
  input            custom_dma_clock_0_out_read_data_valid_pll_s1;
  input            custom_dma_clock_0_out_requests_pll_s1;
  input            custom_dma_clock_0_out_write;
  input   [ 15: 0] custom_dma_clock_0_out_writedata;
  input            d1_pll_s1_end_xfer;
  input   [ 15: 0] pll_s1_readdata_from_sa;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [  3: 0] custom_dma_clock_0_out_address_last_time;
  wire    [  3: 0] custom_dma_clock_0_out_address_to_slave;
  reg     [  1: 0] custom_dma_clock_0_out_byteenable_last_time;
  reg              custom_dma_clock_0_out_read_last_time;
  wire    [ 15: 0] custom_dma_clock_0_out_readdata;
  wire             custom_dma_clock_0_out_reset_n;
  wire             custom_dma_clock_0_out_run;
  wire             custom_dma_clock_0_out_waitrequest;
  reg              custom_dma_clock_0_out_write_last_time;
  reg     [ 15: 0] custom_dma_clock_0_out_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & ((~custom_dma_clock_0_out_qualified_request_pll_s1 | ~custom_dma_clock_0_out_read | (1 & ~d1_pll_s1_end_xfer & custom_dma_clock_0_out_read))) & ((~custom_dma_clock_0_out_qualified_request_pll_s1 | ~custom_dma_clock_0_out_write | (1 & custom_dma_clock_0_out_write)));

  //cascaded wait assignment, which is an e_assign
  assign custom_dma_clock_0_out_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign custom_dma_clock_0_out_address_to_slave = custom_dma_clock_0_out_address;

  //custom_dma_clock_0/out readdata mux, which is an e_mux
  assign custom_dma_clock_0_out_readdata = pll_s1_readdata_from_sa;

  //actual waitrequest port, which is an e_assign
  assign custom_dma_clock_0_out_waitrequest = ~custom_dma_clock_0_out_run;

  //custom_dma_clock_0_out_reset_n assignment, which is an e_assign
  assign custom_dma_clock_0_out_reset_n = reset_n;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //custom_dma_clock_0_out_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_out_address_last_time <= 0;
      else 
        custom_dma_clock_0_out_address_last_time <= custom_dma_clock_0_out_address;
    end


  //custom_dma_clock_0/out waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= custom_dma_clock_0_out_waitrequest & (custom_dma_clock_0_out_read | custom_dma_clock_0_out_write);
    end


  //custom_dma_clock_0_out_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_clock_0_out_address != custom_dma_clock_0_out_address_last_time))
        begin
          $write("%0d ns: custom_dma_clock_0_out_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_clock_0_out_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_out_byteenable_last_time <= 0;
      else 
        custom_dma_clock_0_out_byteenable_last_time <= custom_dma_clock_0_out_byteenable;
    end


  //custom_dma_clock_0_out_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_clock_0_out_byteenable != custom_dma_clock_0_out_byteenable_last_time))
        begin
          $write("%0d ns: custom_dma_clock_0_out_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_clock_0_out_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_out_read_last_time <= 0;
      else 
        custom_dma_clock_0_out_read_last_time <= custom_dma_clock_0_out_read;
    end


  //custom_dma_clock_0_out_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_clock_0_out_read != custom_dma_clock_0_out_read_last_time))
        begin
          $write("%0d ns: custom_dma_clock_0_out_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_clock_0_out_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_out_write_last_time <= 0;
      else 
        custom_dma_clock_0_out_write_last_time <= custom_dma_clock_0_out_write;
    end


  //custom_dma_clock_0_out_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_clock_0_out_write != custom_dma_clock_0_out_write_last_time))
        begin
          $write("%0d ns: custom_dma_clock_0_out_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //custom_dma_clock_0_out_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_clock_0_out_writedata_last_time <= 0;
      else 
        custom_dma_clock_0_out_writedata_last_time <= custom_dma_clock_0_out_writedata;
    end


  //custom_dma_clock_0_out_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (custom_dma_clock_0_out_writedata != custom_dma_clock_0_out_writedata_last_time) & custom_dma_clock_0_out_write)
        begin
          $write("%0d ns: custom_dma_clock_0_out_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module burstcount_fifo_for_ddr_sdram_s1_module (
                                                 // inputs:
                                                  clear_fifo,
                                                  clk,
                                                  data_in,
                                                  read,
                                                  reset_n,
                                                  sync_reset,
                                                  write,

                                                 // outputs:
                                                  data_out,
                                                  empty,
                                                  fifo_contains_ones_n,
                                                  full
                                               )
;

  output  [  2: 0] data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input   [  2: 0] data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire    [  2: 0] data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  wire             full_16;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire    [  2: 0] p0_stage_0;
  wire             p10_full_10;
  wire    [  2: 0] p10_stage_10;
  wire             p11_full_11;
  wire    [  2: 0] p11_stage_11;
  wire             p12_full_12;
  wire    [  2: 0] p12_stage_12;
  wire             p13_full_13;
  wire    [  2: 0] p13_stage_13;
  wire             p14_full_14;
  wire    [  2: 0] p14_stage_14;
  wire             p15_full_15;
  wire    [  2: 0] p15_stage_15;
  wire             p1_full_1;
  wire    [  2: 0] p1_stage_1;
  wire             p2_full_2;
  wire    [  2: 0] p2_stage_2;
  wire             p3_full_3;
  wire    [  2: 0] p3_stage_3;
  wire             p4_full_4;
  wire    [  2: 0] p4_stage_4;
  wire             p5_full_5;
  wire    [  2: 0] p5_stage_5;
  wire             p6_full_6;
  wire    [  2: 0] p6_stage_6;
  wire             p7_full_7;
  wire    [  2: 0] p7_stage_7;
  wire             p8_full_8;
  wire    [  2: 0] p8_stage_8;
  wire             p9_full_9;
  wire    [  2: 0] p9_stage_9;
  reg     [  2: 0] stage_0;
  reg     [  2: 0] stage_1;
  reg     [  2: 0] stage_10;
  reg     [  2: 0] stage_11;
  reg     [  2: 0] stage_12;
  reg     [  2: 0] stage_13;
  reg     [  2: 0] stage_14;
  reg     [  2: 0] stage_15;
  reg     [  2: 0] stage_2;
  reg     [  2: 0] stage_3;
  reg     [  2: 0] stage_4;
  reg     [  2: 0] stage_5;
  reg     [  2: 0] stage_6;
  reg     [  2: 0] stage_7;
  reg     [  2: 0] stage_8;
  reg     [  2: 0] stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_15;
  assign empty = !full_0;
  assign full_16 = 0;
  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    0;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_custom_dma_burst_3_downstream_to_ddr_sdram_s1_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  wire             full_16;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_15;
  assign empty = !full_0;
  assign full_16 = 0;
  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    0;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_custom_dma_burst_4_downstream_to_ddr_sdram_s1_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  wire             full_16;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_15;
  assign empty = !full_0;
  assign full_16 = 0;
  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    0;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_custom_dma_burst_5_downstream_to_ddr_sdram_s1_module (
                                                                           // inputs:
                                                                            clear_fifo,
                                                                            clk,
                                                                            data_in,
                                                                            read,
                                                                            reset_n,
                                                                            sync_reset,
                                                                            write,

                                                                           // outputs:
                                                                            data_out,
                                                                            empty,
                                                                            fifo_contains_ones_n,
                                                                            full
                                                                         )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_10;
  reg              full_11;
  reg              full_12;
  reg              full_13;
  reg              full_14;
  reg              full_15;
  wire             full_16;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  reg              full_7;
  reg              full_8;
  reg              full_9;
  reg     [  5: 0] how_many_ones;
  wire    [  5: 0] one_count_minus_one;
  wire    [  5: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p10_full_10;
  wire             p10_stage_10;
  wire             p11_full_11;
  wire             p11_stage_11;
  wire             p12_full_12;
  wire             p12_stage_12;
  wire             p13_full_13;
  wire             p13_stage_13;
  wire             p14_full_14;
  wire             p14_stage_14;
  wire             p15_full_15;
  wire             p15_stage_15;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  wire             p7_full_7;
  wire             p7_stage_7;
  wire             p8_full_8;
  wire             p8_stage_8;
  wire             p9_full_9;
  wire             p9_stage_9;
  reg              stage_0;
  reg              stage_1;
  reg              stage_10;
  reg              stage_11;
  reg              stage_12;
  reg              stage_13;
  reg              stage_14;
  reg              stage_15;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  reg              stage_7;
  reg              stage_8;
  reg              stage_9;
  wire    [  5: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_15;
  assign empty = !full_0;
  assign full_16 = 0;
  //data_15, which is an e_mux
  assign p15_stage_15 = ((full_16 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_15 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_15))
          if (sync_reset & full_15 & !((full_16 == 0) & read & write))
              stage_15 <= 0;
          else 
            stage_15 <= p15_stage_15;
    end


  //control_15, which is an e_mux
  assign p15_full_15 = ((read & !write) == 0)? full_14 :
    0;

  //control_reg_15, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_15 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_15 <= 0;
          else 
            full_15 <= p15_full_15;
    end


  //data_14, which is an e_mux
  assign p14_stage_14 = ((full_15 & ~clear_fifo) == 0)? data_in :
    stage_15;

  //data_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_14 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_14))
          if (sync_reset & full_14 & !((full_15 == 0) & read & write))
              stage_14 <= 0;
          else 
            stage_14 <= p14_stage_14;
    end


  //control_14, which is an e_mux
  assign p14_full_14 = ((read & !write) == 0)? full_13 :
    full_15;

  //control_reg_14, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_14 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_14 <= 0;
          else 
            full_14 <= p14_full_14;
    end


  //data_13, which is an e_mux
  assign p13_stage_13 = ((full_14 & ~clear_fifo) == 0)? data_in :
    stage_14;

  //data_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_13 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_13))
          if (sync_reset & full_13 & !((full_14 == 0) & read & write))
              stage_13 <= 0;
          else 
            stage_13 <= p13_stage_13;
    end


  //control_13, which is an e_mux
  assign p13_full_13 = ((read & !write) == 0)? full_12 :
    full_14;

  //control_reg_13, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_13 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_13 <= 0;
          else 
            full_13 <= p13_full_13;
    end


  //data_12, which is an e_mux
  assign p12_stage_12 = ((full_13 & ~clear_fifo) == 0)? data_in :
    stage_13;

  //data_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_12 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_12))
          if (sync_reset & full_12 & !((full_13 == 0) & read & write))
              stage_12 <= 0;
          else 
            stage_12 <= p12_stage_12;
    end


  //control_12, which is an e_mux
  assign p12_full_12 = ((read & !write) == 0)? full_11 :
    full_13;

  //control_reg_12, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_12 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_12 <= 0;
          else 
            full_12 <= p12_full_12;
    end


  //data_11, which is an e_mux
  assign p11_stage_11 = ((full_12 & ~clear_fifo) == 0)? data_in :
    stage_12;

  //data_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_11 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_11))
          if (sync_reset & full_11 & !((full_12 == 0) & read & write))
              stage_11 <= 0;
          else 
            stage_11 <= p11_stage_11;
    end


  //control_11, which is an e_mux
  assign p11_full_11 = ((read & !write) == 0)? full_10 :
    full_12;

  //control_reg_11, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_11 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_11 <= 0;
          else 
            full_11 <= p11_full_11;
    end


  //data_10, which is an e_mux
  assign p10_stage_10 = ((full_11 & ~clear_fifo) == 0)? data_in :
    stage_11;

  //data_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_10 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_10))
          if (sync_reset & full_10 & !((full_11 == 0) & read & write))
              stage_10 <= 0;
          else 
            stage_10 <= p10_stage_10;
    end


  //control_10, which is an e_mux
  assign p10_full_10 = ((read & !write) == 0)? full_9 :
    full_11;

  //control_reg_10, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_10 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_10 <= 0;
          else 
            full_10 <= p10_full_10;
    end


  //data_9, which is an e_mux
  assign p9_stage_9 = ((full_10 & ~clear_fifo) == 0)? data_in :
    stage_10;

  //data_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_9 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_9))
          if (sync_reset & full_9 & !((full_10 == 0) & read & write))
              stage_9 <= 0;
          else 
            stage_9 <= p9_stage_9;
    end


  //control_9, which is an e_mux
  assign p9_full_9 = ((read & !write) == 0)? full_8 :
    full_10;

  //control_reg_9, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_9 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_9 <= 0;
          else 
            full_9 <= p9_full_9;
    end


  //data_8, which is an e_mux
  assign p8_stage_8 = ((full_9 & ~clear_fifo) == 0)? data_in :
    stage_9;

  //data_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_8 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_8))
          if (sync_reset & full_8 & !((full_9 == 0) & read & write))
              stage_8 <= 0;
          else 
            stage_8 <= p8_stage_8;
    end


  //control_8, which is an e_mux
  assign p8_full_8 = ((read & !write) == 0)? full_7 :
    full_9;

  //control_reg_8, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_8 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_8 <= 0;
          else 
            full_8 <= p8_full_8;
    end


  //data_7, which is an e_mux
  assign p7_stage_7 = ((full_8 & ~clear_fifo) == 0)? data_in :
    stage_8;

  //data_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_7 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_7))
          if (sync_reset & full_7 & !((full_8 == 0) & read & write))
              stage_7 <= 0;
          else 
            stage_7 <= p7_stage_7;
    end


  //control_7, which is an e_mux
  assign p7_full_7 = ((read & !write) == 0)? full_6 :
    full_8;

  //control_reg_7, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_7 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_7 <= 0;
          else 
            full_7 <= p7_full_7;
    end


  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    stage_7;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    full_7;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_s1_arbitrator (
                                 // inputs:
                                  clk,
                                  custom_dma_burst_3_downstream_address_to_slave,
                                  custom_dma_burst_3_downstream_arbitrationshare,
                                  custom_dma_burst_3_downstream_burstcount,
                                  custom_dma_burst_3_downstream_byteenable,
                                  custom_dma_burst_3_downstream_latency_counter,
                                  custom_dma_burst_3_downstream_read,
                                  custom_dma_burst_3_downstream_write,
                                  custom_dma_burst_3_downstream_writedata,
                                  custom_dma_burst_4_downstream_address_to_slave,
                                  custom_dma_burst_4_downstream_arbitrationshare,
                                  custom_dma_burst_4_downstream_burstcount,
                                  custom_dma_burst_4_downstream_byteenable,
                                  custom_dma_burst_4_downstream_latency_counter,
                                  custom_dma_burst_4_downstream_read,
                                  custom_dma_burst_4_downstream_write,
                                  custom_dma_burst_4_downstream_writedata,
                                  custom_dma_burst_5_downstream_address_to_slave,
                                  custom_dma_burst_5_downstream_arbitrationshare,
                                  custom_dma_burst_5_downstream_burstcount,
                                  custom_dma_burst_5_downstream_byteenable,
                                  custom_dma_burst_5_downstream_latency_counter,
                                  custom_dma_burst_5_downstream_read,
                                  custom_dma_burst_5_downstream_write,
                                  custom_dma_burst_5_downstream_writedata,
                                  ddr_sdram_s1_readdata,
                                  ddr_sdram_s1_readdatavalid,
                                  ddr_sdram_s1_waitrequest_n,
                                  reset_n,

                                 // outputs:
                                  custom_dma_burst_3_downstream_granted_ddr_sdram_s1,
                                  custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1,
                                  custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1,
                                  custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                  custom_dma_burst_3_downstream_requests_ddr_sdram_s1,
                                  custom_dma_burst_4_downstream_granted_ddr_sdram_s1,
                                  custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1,
                                  custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1,
                                  custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                  custom_dma_burst_4_downstream_requests_ddr_sdram_s1,
                                  custom_dma_burst_5_downstream_granted_ddr_sdram_s1,
                                  custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1,
                                  custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1,
                                  custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register,
                                  custom_dma_burst_5_downstream_requests_ddr_sdram_s1,
                                  d1_ddr_sdram_s1_end_xfer,
                                  ddr_sdram_s1_address,
                                  ddr_sdram_s1_beginbursttransfer,
                                  ddr_sdram_s1_burstcount,
                                  ddr_sdram_s1_byteenable,
                                  ddr_sdram_s1_read,
                                  ddr_sdram_s1_readdata_from_sa,
                                  ddr_sdram_s1_reset_n,
                                  ddr_sdram_s1_waitrequest_n_from_sa,
                                  ddr_sdram_s1_write,
                                  ddr_sdram_s1_writedata
                               )
;

  output           custom_dma_burst_3_downstream_granted_ddr_sdram_s1;
  output           custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1;
  output           custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1;
  output           custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  output           custom_dma_burst_3_downstream_requests_ddr_sdram_s1;
  output           custom_dma_burst_4_downstream_granted_ddr_sdram_s1;
  output           custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1;
  output           custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1;
  output           custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  output           custom_dma_burst_4_downstream_requests_ddr_sdram_s1;
  output           custom_dma_burst_5_downstream_granted_ddr_sdram_s1;
  output           custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1;
  output           custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1;
  output           custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  output           custom_dma_burst_5_downstream_requests_ddr_sdram_s1;
  output           d1_ddr_sdram_s1_end_xfer;
  output  [ 22: 0] ddr_sdram_s1_address;
  output           ddr_sdram_s1_beginbursttransfer;
  output  [  2: 0] ddr_sdram_s1_burstcount;
  output  [  3: 0] ddr_sdram_s1_byteenable;
  output           ddr_sdram_s1_read;
  output  [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  output           ddr_sdram_s1_reset_n;
  output           ddr_sdram_s1_waitrequest_n_from_sa;
  output           ddr_sdram_s1_write;
  output  [ 31: 0] ddr_sdram_s1_writedata;
  input            clk;
  input   [ 24: 0] custom_dma_burst_3_downstream_address_to_slave;
  input   [  3: 0] custom_dma_burst_3_downstream_arbitrationshare;
  input   [  2: 0] custom_dma_burst_3_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_3_downstream_byteenable;
  input            custom_dma_burst_3_downstream_latency_counter;
  input            custom_dma_burst_3_downstream_read;
  input            custom_dma_burst_3_downstream_write;
  input   [ 31: 0] custom_dma_burst_3_downstream_writedata;
  input   [ 24: 0] custom_dma_burst_4_downstream_address_to_slave;
  input   [  3: 0] custom_dma_burst_4_downstream_arbitrationshare;
  input   [  2: 0] custom_dma_burst_4_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_4_downstream_byteenable;
  input            custom_dma_burst_4_downstream_latency_counter;
  input            custom_dma_burst_4_downstream_read;
  input            custom_dma_burst_4_downstream_write;
  input   [ 31: 0] custom_dma_burst_4_downstream_writedata;
  input   [ 24: 0] custom_dma_burst_5_downstream_address_to_slave;
  input   [  2: 0] custom_dma_burst_5_downstream_arbitrationshare;
  input   [  2: 0] custom_dma_burst_5_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_5_downstream_byteenable;
  input            custom_dma_burst_5_downstream_latency_counter;
  input            custom_dma_burst_5_downstream_read;
  input            custom_dma_burst_5_downstream_write;
  input   [ 31: 0] custom_dma_burst_5_downstream_writedata;
  input   [ 31: 0] ddr_sdram_s1_readdata;
  input            ddr_sdram_s1_readdatavalid;
  input            ddr_sdram_s1_waitrequest_n;
  input            reset_n;

  wire             custom_dma_burst_3_downstream_arbiterlock;
  wire             custom_dma_burst_3_downstream_arbiterlock2;
  wire             custom_dma_burst_3_downstream_continuerequest;
  wire             custom_dma_burst_3_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_rdv_fifo_empty_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_rdv_fifo_output_from_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire             custom_dma_burst_3_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_arbiterlock;
  wire             custom_dma_burst_4_downstream_arbiterlock2;
  wire             custom_dma_burst_4_downstream_continuerequest;
  wire             custom_dma_burst_4_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_rdv_fifo_empty_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_rdv_fifo_output_from_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire             custom_dma_burst_4_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_arbiterlock;
  wire             custom_dma_burst_5_downstream_arbiterlock2;
  wire             custom_dma_burst_5_downstream_continuerequest;
  wire             custom_dma_burst_5_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_rdv_fifo_empty_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_rdv_fifo_output_from_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire             custom_dma_burst_5_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1;
  reg              d1_ddr_sdram_s1_end_xfer;
  reg              d1_reasons_to_wait;
  wire    [ 22: 0] ddr_sdram_s1_address;
  wire             ddr_sdram_s1_allgrants;
  wire             ddr_sdram_s1_allow_new_arb_cycle;
  wire             ddr_sdram_s1_any_bursting_master_saved_grant;
  wire             ddr_sdram_s1_any_continuerequest;
  reg     [  2: 0] ddr_sdram_s1_arb_addend;
  wire             ddr_sdram_s1_arb_counter_enable;
  reg     [  3: 0] ddr_sdram_s1_arb_share_counter;
  wire    [  3: 0] ddr_sdram_s1_arb_share_counter_next_value;
  wire    [  3: 0] ddr_sdram_s1_arb_share_set_values;
  wire    [  2: 0] ddr_sdram_s1_arb_winner;
  wire             ddr_sdram_s1_arbitration_holdoff_internal;
  reg     [  1: 0] ddr_sdram_s1_bbt_burstcounter;
  wire             ddr_sdram_s1_beginbursttransfer;
  wire             ddr_sdram_s1_beginbursttransfer_internal;
  wire             ddr_sdram_s1_begins_xfer;
  wire    [  2: 0] ddr_sdram_s1_burstcount;
  wire             ddr_sdram_s1_burstcount_fifo_empty;
  wire    [  3: 0] ddr_sdram_s1_byteenable;
  wire    [  5: 0] ddr_sdram_s1_chosen_master_double_vector;
  wire    [  2: 0] ddr_sdram_s1_chosen_master_rot_left;
  reg     [  2: 0] ddr_sdram_s1_current_burst;
  wire    [  2: 0] ddr_sdram_s1_current_burst_minus_one;
  wire             ddr_sdram_s1_end_xfer;
  wire             ddr_sdram_s1_firsttransfer;
  wire    [  2: 0] ddr_sdram_s1_grant_vector;
  wire             ddr_sdram_s1_in_a_read_cycle;
  wire             ddr_sdram_s1_in_a_write_cycle;
  reg              ddr_sdram_s1_load_fifo;
  wire    [  2: 0] ddr_sdram_s1_master_qreq_vector;
  wire             ddr_sdram_s1_move_on_to_next_transaction;
  wire    [  1: 0] ddr_sdram_s1_next_bbt_burstcount;
  wire    [  2: 0] ddr_sdram_s1_next_burst_count;
  wire             ddr_sdram_s1_non_bursting_master_requests;
  wire             ddr_sdram_s1_read;
  wire    [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  wire             ddr_sdram_s1_readdatavalid_from_sa;
  reg              ddr_sdram_s1_reg_firsttransfer;
  wire             ddr_sdram_s1_reset_n;
  reg     [  2: 0] ddr_sdram_s1_saved_chosen_master_vector;
  wire    [  2: 0] ddr_sdram_s1_selected_burstcount;
  reg              ddr_sdram_s1_slavearbiterlockenable;
  wire             ddr_sdram_s1_slavearbiterlockenable2;
  wire             ddr_sdram_s1_this_cycle_is_the_last_burst;
  wire    [  2: 0] ddr_sdram_s1_transaction_burst_count;
  wire             ddr_sdram_s1_unreg_firsttransfer;
  wire             ddr_sdram_s1_waitrequest_n_from_sa;
  wire             ddr_sdram_s1_waits_for_read;
  wire             ddr_sdram_s1_waits_for_write;
  wire             ddr_sdram_s1_write;
  wire    [ 31: 0] ddr_sdram_s1_writedata;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ddr_sdram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1;
  reg              last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1;
  reg              last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1;
  wire             p0_ddr_sdram_s1_load_fifo;
  wire    [ 24: 0] shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_3_downstream;
  wire    [ 24: 0] shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_4_downstream;
  wire    [ 24: 0] shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_5_downstream;
  wire             wait_for_ddr_sdram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ddr_sdram_s1_end_xfer;
    end


  assign ddr_sdram_s1_begins_xfer = ~d1_reasons_to_wait & ((custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1 | custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1 | custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1));
  //assign ddr_sdram_s1_readdata_from_sa = ddr_sdram_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_s1_readdata_from_sa = ddr_sdram_s1_readdata;

  assign custom_dma_burst_3_downstream_requests_ddr_sdram_s1 = (1) & (custom_dma_burst_3_downstream_read | custom_dma_burst_3_downstream_write);
  //assign ddr_sdram_s1_waitrequest_n_from_sa = ddr_sdram_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_s1_waitrequest_n_from_sa = ddr_sdram_s1_waitrequest_n;

  //assign ddr_sdram_s1_readdatavalid_from_sa = ddr_sdram_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign ddr_sdram_s1_readdatavalid_from_sa = ddr_sdram_s1_readdatavalid;

  //ddr_sdram_s1_arb_share_counter set values, which is an e_mux
  assign ddr_sdram_s1_arb_share_set_values = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_arbitrationshare :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_arbitrationshare :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_arbitrationshare :
    (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_arbitrationshare :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_arbitrationshare :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_arbitrationshare :
    (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_arbitrationshare :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_arbitrationshare :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_arbitrationshare :
    1;

  //ddr_sdram_s1_non_bursting_master_requests mux, which is an e_mux
  assign ddr_sdram_s1_non_bursting_master_requests = 0;

  //ddr_sdram_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign ddr_sdram_s1_any_bursting_master_saved_grant = custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 |
    custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1;

  //ddr_sdram_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign ddr_sdram_s1_arb_share_counter_next_value = ddr_sdram_s1_firsttransfer ? (ddr_sdram_s1_arb_share_set_values - 1) : |ddr_sdram_s1_arb_share_counter ? (ddr_sdram_s1_arb_share_counter - 1) : 0;

  //ddr_sdram_s1_allgrants all slave grants, which is an e_mux
  assign ddr_sdram_s1_allgrants = (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector) |
    (|ddr_sdram_s1_grant_vector);

  //ddr_sdram_s1_end_xfer assignment, which is an e_assign
  assign ddr_sdram_s1_end_xfer = ~(ddr_sdram_s1_waits_for_read | ddr_sdram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ddr_sdram_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ddr_sdram_s1 = ddr_sdram_s1_end_xfer & (~ddr_sdram_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ddr_sdram_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign ddr_sdram_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_ddr_sdram_s1 & ddr_sdram_s1_allgrants) | (end_xfer_arb_share_counter_term_ddr_sdram_s1 & ~ddr_sdram_s1_non_bursting_master_requests);

  //ddr_sdram_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_arb_share_counter <= 0;
      else if (ddr_sdram_s1_arb_counter_enable)
          ddr_sdram_s1_arb_share_counter <= ddr_sdram_s1_arb_share_counter_next_value;
    end


  //ddr_sdram_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_slavearbiterlockenable <= 0;
      else if ((|ddr_sdram_s1_master_qreq_vector & end_xfer_arb_share_counter_term_ddr_sdram_s1) | (end_xfer_arb_share_counter_term_ddr_sdram_s1 & ~ddr_sdram_s1_non_bursting_master_requests))
          ddr_sdram_s1_slavearbiterlockenable <= |ddr_sdram_s1_arb_share_counter_next_value;
    end


  //custom_dma_burst_3/downstream ddr_sdram/s1 arbiterlock, which is an e_assign
  assign custom_dma_burst_3_downstream_arbiterlock = ddr_sdram_s1_slavearbiterlockenable & custom_dma_burst_3_downstream_continuerequest;

  //ddr_sdram_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ddr_sdram_s1_slavearbiterlockenable2 = |ddr_sdram_s1_arb_share_counter_next_value;

  //custom_dma_burst_3/downstream ddr_sdram/s1 arbiterlock2, which is an e_assign
  assign custom_dma_burst_3_downstream_arbiterlock2 = ddr_sdram_s1_slavearbiterlockenable2 & custom_dma_burst_3_downstream_continuerequest;

  //custom_dma_burst_4/downstream ddr_sdram/s1 arbiterlock, which is an e_assign
  assign custom_dma_burst_4_downstream_arbiterlock = ddr_sdram_s1_slavearbiterlockenable & custom_dma_burst_4_downstream_continuerequest;

  //custom_dma_burst_4/downstream ddr_sdram/s1 arbiterlock2, which is an e_assign
  assign custom_dma_burst_4_downstream_arbiterlock2 = ddr_sdram_s1_slavearbiterlockenable2 & custom_dma_burst_4_downstream_continuerequest;

  //custom_dma_burst_4/downstream granted ddr_sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1 <= custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 ? 1 : (ddr_sdram_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1;
    end


  //custom_dma_burst_4_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_4_downstream_continuerequest = (last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1 & 1) |
    (last_cycle_custom_dma_burst_4_downstream_granted_slave_ddr_sdram_s1 & 1);

  //ddr_sdram_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ddr_sdram_s1_any_continuerequest = custom_dma_burst_4_downstream_continuerequest |
    custom_dma_burst_5_downstream_continuerequest |
    custom_dma_burst_3_downstream_continuerequest |
    custom_dma_burst_5_downstream_continuerequest |
    custom_dma_burst_3_downstream_continuerequest |
    custom_dma_burst_4_downstream_continuerequest;

  //custom_dma_burst_5/downstream ddr_sdram/s1 arbiterlock, which is an e_assign
  assign custom_dma_burst_5_downstream_arbiterlock = ddr_sdram_s1_slavearbiterlockenable & custom_dma_burst_5_downstream_continuerequest;

  //custom_dma_burst_5/downstream ddr_sdram/s1 arbiterlock2, which is an e_assign
  assign custom_dma_burst_5_downstream_arbiterlock2 = ddr_sdram_s1_slavearbiterlockenable2 & custom_dma_burst_5_downstream_continuerequest;

  //custom_dma_burst_5/downstream granted ddr_sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1 <= custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1 ? 1 : (ddr_sdram_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1;
    end


  //custom_dma_burst_5_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_5_downstream_continuerequest = (last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1 & 1) |
    (last_cycle_custom_dma_burst_5_downstream_granted_slave_ddr_sdram_s1 & 1);

  assign custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1 = custom_dma_burst_3_downstream_requests_ddr_sdram_s1 & ~((custom_dma_burst_3_downstream_read & ((custom_dma_burst_3_downstream_latency_counter != 0) | (1 < custom_dma_burst_3_downstream_latency_counter))) | custom_dma_burst_4_downstream_arbiterlock | custom_dma_burst_5_downstream_arbiterlock);
  //unique name for ddr_sdram_s1_move_on_to_next_transaction, which is an e_assign
  assign ddr_sdram_s1_move_on_to_next_transaction = ddr_sdram_s1_this_cycle_is_the_last_burst & ddr_sdram_s1_load_fifo;

  //the currently selected burstcount for ddr_sdram_s1, which is an e_mux
  assign ddr_sdram_s1_selected_burstcount = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_burstcount :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_burstcount :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_burstcount :
    1;

  //burstcount_fifo_for_ddr_sdram_s1, which is an e_fifo_with_registered_outputs
  burstcount_fifo_for_ddr_sdram_s1_module burstcount_fifo_for_ddr_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (ddr_sdram_s1_selected_burstcount),
      .data_out             (ddr_sdram_s1_transaction_burst_count),
      .empty                (ddr_sdram_s1_burstcount_fifo_empty),
      .fifo_contains_ones_n (),
      .full                 (),
      .read                 (ddr_sdram_s1_this_cycle_is_the_last_burst),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr_sdram_s1_waits_for_read & ddr_sdram_s1_load_fifo & ~(ddr_sdram_s1_this_cycle_is_the_last_burst & ddr_sdram_s1_burstcount_fifo_empty))
    );

  //ddr_sdram_s1 current burst minus one, which is an e_assign
  assign ddr_sdram_s1_current_burst_minus_one = ddr_sdram_s1_current_burst - 1;

  //what to load in current_burst, for ddr_sdram_s1, which is an e_mux
  assign ddr_sdram_s1_next_burst_count = (((in_a_read_cycle & ~ddr_sdram_s1_waits_for_read) & ~ddr_sdram_s1_load_fifo))? ddr_sdram_s1_selected_burstcount :
    ((in_a_read_cycle & ~ddr_sdram_s1_waits_for_read & ddr_sdram_s1_this_cycle_is_the_last_burst & ddr_sdram_s1_burstcount_fifo_empty))? ddr_sdram_s1_selected_burstcount :
    (ddr_sdram_s1_this_cycle_is_the_last_burst)? ddr_sdram_s1_transaction_burst_count :
    ddr_sdram_s1_current_burst_minus_one;

  //the current burst count for ddr_sdram_s1, to be decremented, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_current_burst <= 0;
      else if (ddr_sdram_s1_readdatavalid_from_sa | (~ddr_sdram_s1_load_fifo & (in_a_read_cycle & ~ddr_sdram_s1_waits_for_read)))
          ddr_sdram_s1_current_burst <= ddr_sdram_s1_next_burst_count;
    end


  //a 1 or burstcount fifo empty, to initialize the counter, which is an e_mux
  assign p0_ddr_sdram_s1_load_fifo = (~ddr_sdram_s1_load_fifo)? 1 :
    (((in_a_read_cycle & ~ddr_sdram_s1_waits_for_read) & ddr_sdram_s1_load_fifo))? 1 :
    ~ddr_sdram_s1_burstcount_fifo_empty;

  //whether to load directly to the counter or to the fifo, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_load_fifo <= 0;
      else if ((in_a_read_cycle & ~ddr_sdram_s1_waits_for_read) & ~ddr_sdram_s1_load_fifo | ddr_sdram_s1_this_cycle_is_the_last_burst)
          ddr_sdram_s1_load_fifo <= p0_ddr_sdram_s1_load_fifo;
    end


  //the last cycle in the burst for ddr_sdram_s1, which is an e_assign
  assign ddr_sdram_s1_this_cycle_is_the_last_burst = ~(|ddr_sdram_s1_current_burst_minus_one) & ddr_sdram_s1_readdatavalid_from_sa;

  //rdv_fifo_for_custom_dma_burst_3_downstream_to_ddr_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_custom_dma_burst_3_downstream_to_ddr_sdram_s1_module rdv_fifo_for_custom_dma_burst_3_downstream_to_ddr_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_3_downstream_granted_ddr_sdram_s1),
      .data_out             (custom_dma_burst_3_downstream_rdv_fifo_output_from_ddr_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (custom_dma_burst_3_downstream_rdv_fifo_empty_ddr_sdram_s1),
      .full                 (),
      .read                 (ddr_sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr_sdram_s1_waits_for_read)
    );

  assign custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register = ~custom_dma_burst_3_downstream_rdv_fifo_empty_ddr_sdram_s1;
  //local readdatavalid custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1, which is an e_mux
  assign custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1 = (ddr_sdram_s1_readdatavalid_from_sa & custom_dma_burst_3_downstream_rdv_fifo_output_from_ddr_sdram_s1) & ~ custom_dma_burst_3_downstream_rdv_fifo_empty_ddr_sdram_s1;

  //ddr_sdram_s1_writedata mux, which is an e_mux
  assign ddr_sdram_s1_writedata = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_writedata :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_writedata :
    custom_dma_burst_5_downstream_writedata;

  assign custom_dma_burst_4_downstream_requests_ddr_sdram_s1 = (1) & (custom_dma_burst_4_downstream_read | custom_dma_burst_4_downstream_write);
  //custom_dma_burst_3/downstream granted ddr_sdram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1 <= custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 ? 1 : (ddr_sdram_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1;
    end


  //custom_dma_burst_3_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_3_downstream_continuerequest = (last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1 & 1) |
    (last_cycle_custom_dma_burst_3_downstream_granted_slave_ddr_sdram_s1 & 1);

  assign custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1 = custom_dma_burst_4_downstream_requests_ddr_sdram_s1 & ~((custom_dma_burst_4_downstream_read & ((custom_dma_burst_4_downstream_latency_counter != 0) | (1 < custom_dma_burst_4_downstream_latency_counter))) | custom_dma_burst_3_downstream_arbiterlock | custom_dma_burst_5_downstream_arbiterlock);
  //rdv_fifo_for_custom_dma_burst_4_downstream_to_ddr_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_custom_dma_burst_4_downstream_to_ddr_sdram_s1_module rdv_fifo_for_custom_dma_burst_4_downstream_to_ddr_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_4_downstream_granted_ddr_sdram_s1),
      .data_out             (custom_dma_burst_4_downstream_rdv_fifo_output_from_ddr_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (custom_dma_burst_4_downstream_rdv_fifo_empty_ddr_sdram_s1),
      .full                 (),
      .read                 (ddr_sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr_sdram_s1_waits_for_read)
    );

  assign custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register = ~custom_dma_burst_4_downstream_rdv_fifo_empty_ddr_sdram_s1;
  //local readdatavalid custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1, which is an e_mux
  assign custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1 = (ddr_sdram_s1_readdatavalid_from_sa & custom_dma_burst_4_downstream_rdv_fifo_output_from_ddr_sdram_s1) & ~ custom_dma_burst_4_downstream_rdv_fifo_empty_ddr_sdram_s1;

  assign custom_dma_burst_5_downstream_requests_ddr_sdram_s1 = (1) & (custom_dma_burst_5_downstream_read | custom_dma_burst_5_downstream_write);
  assign custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1 = custom_dma_burst_5_downstream_requests_ddr_sdram_s1 & ~((custom_dma_burst_5_downstream_read & ((custom_dma_burst_5_downstream_latency_counter != 0) | (1 < custom_dma_burst_5_downstream_latency_counter))) | custom_dma_burst_3_downstream_arbiterlock | custom_dma_burst_4_downstream_arbiterlock);
  //rdv_fifo_for_custom_dma_burst_5_downstream_to_ddr_sdram_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_custom_dma_burst_5_downstream_to_ddr_sdram_s1_module rdv_fifo_for_custom_dma_burst_5_downstream_to_ddr_sdram_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_5_downstream_granted_ddr_sdram_s1),
      .data_out             (custom_dma_burst_5_downstream_rdv_fifo_output_from_ddr_sdram_s1),
      .empty                (),
      .fifo_contains_ones_n (custom_dma_burst_5_downstream_rdv_fifo_empty_ddr_sdram_s1),
      .full                 (),
      .read                 (ddr_sdram_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~ddr_sdram_s1_waits_for_read)
    );

  assign custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register = ~custom_dma_burst_5_downstream_rdv_fifo_empty_ddr_sdram_s1;
  //local readdatavalid custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1, which is an e_mux
  assign custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1 = (ddr_sdram_s1_readdatavalid_from_sa & custom_dma_burst_5_downstream_rdv_fifo_output_from_ddr_sdram_s1) & ~ custom_dma_burst_5_downstream_rdv_fifo_empty_ddr_sdram_s1;

  //allow new arb cycle for ddr_sdram/s1, which is an e_assign
  assign ddr_sdram_s1_allow_new_arb_cycle = ~custom_dma_burst_3_downstream_arbiterlock & ~custom_dma_burst_4_downstream_arbiterlock & ~custom_dma_burst_5_downstream_arbiterlock;

  //custom_dma_burst_5/downstream assignment into master qualified-requests vector for ddr_sdram/s1, which is an e_assign
  assign ddr_sdram_s1_master_qreq_vector[0] = custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1;

  //custom_dma_burst_5/downstream grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_5_downstream_granted_ddr_sdram_s1 = ddr_sdram_s1_grant_vector[0];

  //custom_dma_burst_5/downstream saved-grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1 = ddr_sdram_s1_arb_winner[0];

  //custom_dma_burst_4/downstream assignment into master qualified-requests vector for ddr_sdram/s1, which is an e_assign
  assign ddr_sdram_s1_master_qreq_vector[1] = custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1;

  //custom_dma_burst_4/downstream grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_4_downstream_granted_ddr_sdram_s1 = ddr_sdram_s1_grant_vector[1];

  //custom_dma_burst_4/downstream saved-grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 = ddr_sdram_s1_arb_winner[1];

  //custom_dma_burst_3/downstream assignment into master qualified-requests vector for ddr_sdram/s1, which is an e_assign
  assign ddr_sdram_s1_master_qreq_vector[2] = custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1;

  //custom_dma_burst_3/downstream grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_3_downstream_granted_ddr_sdram_s1 = ddr_sdram_s1_grant_vector[2];

  //custom_dma_burst_3/downstream saved-grant ddr_sdram/s1, which is an e_assign
  assign custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 = ddr_sdram_s1_arb_winner[2];

  //ddr_sdram/s1 chosen-master double-vector, which is an e_assign
  assign ddr_sdram_s1_chosen_master_double_vector = {ddr_sdram_s1_master_qreq_vector, ddr_sdram_s1_master_qreq_vector} & ({~ddr_sdram_s1_master_qreq_vector, ~ddr_sdram_s1_master_qreq_vector} + ddr_sdram_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign ddr_sdram_s1_arb_winner = (ddr_sdram_s1_allow_new_arb_cycle & | ddr_sdram_s1_grant_vector) ? ddr_sdram_s1_grant_vector : ddr_sdram_s1_saved_chosen_master_vector;

  //saved ddr_sdram_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_saved_chosen_master_vector <= 0;
      else if (ddr_sdram_s1_allow_new_arb_cycle)
          ddr_sdram_s1_saved_chosen_master_vector <= |ddr_sdram_s1_grant_vector ? ddr_sdram_s1_grant_vector : ddr_sdram_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ddr_sdram_s1_grant_vector = {(ddr_sdram_s1_chosen_master_double_vector[2] | ddr_sdram_s1_chosen_master_double_vector[5]),
    (ddr_sdram_s1_chosen_master_double_vector[1] | ddr_sdram_s1_chosen_master_double_vector[4]),
    (ddr_sdram_s1_chosen_master_double_vector[0] | ddr_sdram_s1_chosen_master_double_vector[3])};

  //ddr_sdram/s1 chosen master rotated left, which is an e_assign
  assign ddr_sdram_s1_chosen_master_rot_left = (ddr_sdram_s1_arb_winner << 1) ? (ddr_sdram_s1_arb_winner << 1) : 1;

  //ddr_sdram/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_arb_addend <= 1;
      else if (|ddr_sdram_s1_grant_vector)
          ddr_sdram_s1_arb_addend <= ddr_sdram_s1_end_xfer? ddr_sdram_s1_chosen_master_rot_left : ddr_sdram_s1_grant_vector;
    end


  //ddr_sdram_s1_reset_n assignment, which is an e_assign
  assign ddr_sdram_s1_reset_n = reset_n;

  //ddr_sdram_s1_firsttransfer first transaction, which is an e_assign
  assign ddr_sdram_s1_firsttransfer = ddr_sdram_s1_begins_xfer ? ddr_sdram_s1_unreg_firsttransfer : ddr_sdram_s1_reg_firsttransfer;

  //ddr_sdram_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign ddr_sdram_s1_unreg_firsttransfer = ~(ddr_sdram_s1_slavearbiterlockenable & ddr_sdram_s1_any_continuerequest);

  //ddr_sdram_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_reg_firsttransfer <= 1'b1;
      else if (ddr_sdram_s1_begins_xfer)
          ddr_sdram_s1_reg_firsttransfer <= ddr_sdram_s1_unreg_firsttransfer;
    end


  //ddr_sdram_s1_next_bbt_burstcount next_bbt_burstcount, which is an e_mux
  assign ddr_sdram_s1_next_bbt_burstcount = ((((ddr_sdram_s1_write) && (ddr_sdram_s1_bbt_burstcounter == 0))))? (ddr_sdram_s1_burstcount - 1) :
    ((((ddr_sdram_s1_read) && (ddr_sdram_s1_bbt_burstcounter == 0))))? 0 :
    (ddr_sdram_s1_bbt_burstcounter - 1);

  //ddr_sdram_s1_bbt_burstcounter bbt_burstcounter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ddr_sdram_s1_bbt_burstcounter <= 0;
      else if (ddr_sdram_s1_begins_xfer)
          ddr_sdram_s1_bbt_burstcounter <= ddr_sdram_s1_next_bbt_burstcount;
    end


  //ddr_sdram_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ddr_sdram_s1_beginbursttransfer_internal = ddr_sdram_s1_begins_xfer & (ddr_sdram_s1_bbt_burstcounter == 0);

  //ddr_sdram/s1 begin burst transfer to slave, which is an e_assign
  assign ddr_sdram_s1_beginbursttransfer = ddr_sdram_s1_beginbursttransfer_internal;

  //ddr_sdram_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ddr_sdram_s1_arbitration_holdoff_internal = ddr_sdram_s1_begins_xfer & ddr_sdram_s1_firsttransfer;

  //ddr_sdram_s1_read assignment, which is an e_mux
  assign ddr_sdram_s1_read = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 & custom_dma_burst_3_downstream_read) | (custom_dma_burst_4_downstream_granted_ddr_sdram_s1 & custom_dma_burst_4_downstream_read) | (custom_dma_burst_5_downstream_granted_ddr_sdram_s1 & custom_dma_burst_5_downstream_read);

  //ddr_sdram_s1_write assignment, which is an e_mux
  assign ddr_sdram_s1_write = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 & custom_dma_burst_3_downstream_write) | (custom_dma_burst_4_downstream_granted_ddr_sdram_s1 & custom_dma_burst_4_downstream_write) | (custom_dma_burst_5_downstream_granted_ddr_sdram_s1 & custom_dma_burst_5_downstream_write);

  assign shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_3_downstream = custom_dma_burst_3_downstream_address_to_slave;
  //ddr_sdram_s1_address mux, which is an e_mux
  assign ddr_sdram_s1_address = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? (shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_3_downstream >> 2) :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? (shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_4_downstream >> 2) :
    (shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_5_downstream >> 2);

  assign shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_4_downstream = custom_dma_burst_4_downstream_address_to_slave;
  assign shifted_address_to_ddr_sdram_s1_from_custom_dma_burst_5_downstream = custom_dma_burst_5_downstream_address_to_slave;
  //d1_ddr_sdram_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ddr_sdram_s1_end_xfer <= 1;
      else 
        d1_ddr_sdram_s1_end_xfer <= ddr_sdram_s1_end_xfer;
    end


  //ddr_sdram_s1_waits_for_read in a cycle, which is an e_mux
  assign ddr_sdram_s1_waits_for_read = ddr_sdram_s1_in_a_read_cycle & ~ddr_sdram_s1_waitrequest_n_from_sa;

  //ddr_sdram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ddr_sdram_s1_in_a_read_cycle = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 & custom_dma_burst_3_downstream_read) | (custom_dma_burst_4_downstream_granted_ddr_sdram_s1 & custom_dma_burst_4_downstream_read) | (custom_dma_burst_5_downstream_granted_ddr_sdram_s1 & custom_dma_burst_5_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ddr_sdram_s1_in_a_read_cycle;

  //ddr_sdram_s1_waits_for_write in a cycle, which is an e_mux
  assign ddr_sdram_s1_waits_for_write = ddr_sdram_s1_in_a_write_cycle & ~ddr_sdram_s1_waitrequest_n_from_sa;

  //ddr_sdram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ddr_sdram_s1_in_a_write_cycle = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 & custom_dma_burst_3_downstream_write) | (custom_dma_burst_4_downstream_granted_ddr_sdram_s1 & custom_dma_burst_4_downstream_write) | (custom_dma_burst_5_downstream_granted_ddr_sdram_s1 & custom_dma_burst_5_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ddr_sdram_s1_in_a_write_cycle;

  assign wait_for_ddr_sdram_s1_counter = 0;
  //ddr_sdram_s1_byteenable byte enable port mux, which is an e_mux
  assign ddr_sdram_s1_byteenable = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_byteenable :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_byteenable :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign ddr_sdram_s1_burstcount = (custom_dma_burst_3_downstream_granted_ddr_sdram_s1)? custom_dma_burst_3_downstream_burstcount :
    (custom_dma_burst_4_downstream_granted_ddr_sdram_s1)? custom_dma_burst_4_downstream_burstcount :
    (custom_dma_burst_5_downstream_granted_ddr_sdram_s1)? custom_dma_burst_5_downstream_burstcount :
    1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ddr_sdram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //custom_dma_burst_3/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_3_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_3_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_3/downstream drove 0 on its 'arbitrationshare' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_3/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_3_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_3_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_3/downstream drove 0 on its 'burstcount' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_4/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_4_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_4_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_4/downstream drove 0 on its 'arbitrationshare' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_4/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_4_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_4_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_4/downstream drove 0 on its 'burstcount' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_5/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_5_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_5_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_5/downstream drove 0 on its 'arbitrationshare' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_5/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_5_downstream_requests_ddr_sdram_s1 && (custom_dma_burst_5_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_5/downstream drove 0 on its 'burstcount' port while accessing slave ddr_sdram/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_3_downstream_granted_ddr_sdram_s1 + custom_dma_burst_4_downstream_granted_ddr_sdram_s1 + custom_dma_burst_5_downstream_granted_ddr_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_3_downstream_saved_grant_ddr_sdram_s1 + custom_dma_burst_4_downstream_saved_grant_ddr_sdram_s1 + custom_dma_burst_5_downstream_saved_grant_ddr_sdram_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_bus_avalon_slave_arbitrator (
                                               // inputs:
                                                clk,
                                                custom_dma_burst_0_downstream_address_to_slave,
                                                custom_dma_burst_0_downstream_arbitrationshare,
                                                custom_dma_burst_0_downstream_burstcount,
                                                custom_dma_burst_0_downstream_byteenable,
                                                custom_dma_burst_0_downstream_latency_counter,
                                                custom_dma_burst_0_downstream_read,
                                                custom_dma_burst_0_downstream_write,
                                                custom_dma_burst_0_downstream_writedata,
                                                fir_dma_read_master_address_to_slave,
                                                fir_dma_read_master_latency_counter,
                                                fir_dma_read_master_read,
                                                reset_n,

                                               // outputs:
                                                adsc_n_to_the_ext_ssram,
                                                bw_n_to_the_ext_ssram,
                                                bwe_n_to_the_ext_ssram,
                                                chipenable1_n_to_the_ext_ssram,
                                                custom_dma_burst_0_downstream_granted_ext_ssram_s1,
                                                custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1,
                                                custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1,
                                                custom_dma_burst_0_downstream_requests_ext_ssram_s1,
                                                d1_ext_ssram_bus_avalon_slave_end_xfer,
                                                ext_ssram_bus_address,
                                                ext_ssram_bus_data,
                                                fir_dma_read_master_granted_ext_ssram_s1,
                                                fir_dma_read_master_qualified_request_ext_ssram_s1,
                                                fir_dma_read_master_read_data_valid_ext_ssram_s1,
                                                fir_dma_read_master_requests_ext_ssram_s1,
                                                incoming_ext_ssram_bus_data,
                                                outputenable_n_to_the_ext_ssram
                                             )
;

  output           adsc_n_to_the_ext_ssram;
  output  [  3: 0] bw_n_to_the_ext_ssram;
  output           bwe_n_to_the_ext_ssram;
  output           chipenable1_n_to_the_ext_ssram;
  output           custom_dma_burst_0_downstream_granted_ext_ssram_s1;
  output           custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1;
  output           custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1;
  output           custom_dma_burst_0_downstream_requests_ext_ssram_s1;
  output           d1_ext_ssram_bus_avalon_slave_end_xfer;
  output  [ 20: 0] ext_ssram_bus_address;
  inout   [ 31: 0] ext_ssram_bus_data;
  output           fir_dma_read_master_granted_ext_ssram_s1;
  output           fir_dma_read_master_qualified_request_ext_ssram_s1;
  output           fir_dma_read_master_read_data_valid_ext_ssram_s1;
  output           fir_dma_read_master_requests_ext_ssram_s1;
  output  [ 31: 0] incoming_ext_ssram_bus_data;
  output           outputenable_n_to_the_ext_ssram;
  input            clk;
  input   [ 20: 0] custom_dma_burst_0_downstream_address_to_slave;
  input   [  3: 0] custom_dma_burst_0_downstream_arbitrationshare;
  input            custom_dma_burst_0_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_0_downstream_byteenable;
  input   [  2: 0] custom_dma_burst_0_downstream_latency_counter;
  input            custom_dma_burst_0_downstream_read;
  input            custom_dma_burst_0_downstream_write;
  input   [ 31: 0] custom_dma_burst_0_downstream_writedata;
  input   [ 31: 0] fir_dma_read_master_address_to_slave;
  input   [  2: 0] fir_dma_read_master_latency_counter;
  input            fir_dma_read_master_read;
  input            reset_n;

  reg              adsc_n_to_the_ext_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg     [  3: 0] bw_n_to_the_ext_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              bwe_n_to_the_ext_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              chipenable1_n_to_the_ext_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             custom_dma_burst_0_downstream_arbiterlock;
  wire             custom_dma_burst_0_downstream_arbiterlock2;
  wire             custom_dma_burst_0_downstream_continuerequest;
  wire             custom_dma_burst_0_downstream_granted_ext_ssram_s1;
  wire             custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1;
  wire             custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1;
  reg     [  3: 0] custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register;
  wire             custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register_in;
  wire             custom_dma_burst_0_downstream_requests_ext_ssram_s1;
  wire             custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1;
  reg              d1_ext_ssram_bus_avalon_slave_end_xfer;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 31: 0] d1_outgoing_ext_ssram_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave;
  reg     [ 20: 0] ext_ssram_bus_address /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             ext_ssram_bus_avalon_slave_allgrants;
  wire             ext_ssram_bus_avalon_slave_allow_new_arb_cycle;
  wire             ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant;
  wire             ext_ssram_bus_avalon_slave_any_continuerequest;
  reg     [  1: 0] ext_ssram_bus_avalon_slave_arb_addend;
  wire             ext_ssram_bus_avalon_slave_arb_counter_enable;
  reg     [  3: 0] ext_ssram_bus_avalon_slave_arb_share_counter;
  wire    [  3: 0] ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
  wire    [  3: 0] ext_ssram_bus_avalon_slave_arb_share_set_values;
  wire    [  1: 0] ext_ssram_bus_avalon_slave_arb_winner;
  wire             ext_ssram_bus_avalon_slave_arbitration_holdoff_internal;
  wire             ext_ssram_bus_avalon_slave_beginbursttransfer_internal;
  wire             ext_ssram_bus_avalon_slave_begins_xfer;
  wire    [  3: 0] ext_ssram_bus_avalon_slave_chosen_master_double_vector;
  wire    [  1: 0] ext_ssram_bus_avalon_slave_chosen_master_rot_left;
  wire             ext_ssram_bus_avalon_slave_end_xfer;
  wire             ext_ssram_bus_avalon_slave_firsttransfer;
  wire    [  1: 0] ext_ssram_bus_avalon_slave_grant_vector;
  wire    [  1: 0] ext_ssram_bus_avalon_slave_master_qreq_vector;
  wire             ext_ssram_bus_avalon_slave_non_bursting_master_requests;
  wire             ext_ssram_bus_avalon_slave_read_pending;
  reg              ext_ssram_bus_avalon_slave_reg_firsttransfer;
  reg     [  1: 0] ext_ssram_bus_avalon_slave_saved_chosen_master_vector;
  reg              ext_ssram_bus_avalon_slave_slavearbiterlockenable;
  wire             ext_ssram_bus_avalon_slave_slavearbiterlockenable2;
  wire             ext_ssram_bus_avalon_slave_unreg_firsttransfer;
  wire             ext_ssram_bus_avalon_slave_write_pending;
  wire    [ 31: 0] ext_ssram_bus_data;
  wire             ext_ssram_s1_in_a_read_cycle;
  wire             ext_ssram_s1_in_a_write_cycle;
  wire             ext_ssram_s1_waits_for_read;
  wire             ext_ssram_s1_waits_for_write;
  wire             ext_ssram_s1_with_write_latency;
  wire             fir_dma_read_master_arbiterlock;
  wire             fir_dma_read_master_arbiterlock2;
  wire             fir_dma_read_master_continuerequest;
  wire             fir_dma_read_master_granted_ext_ssram_s1;
  wire             fir_dma_read_master_qualified_request_ext_ssram_s1;
  wire             fir_dma_read_master_read_data_valid_ext_ssram_s1;
  reg     [  3: 0] fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register;
  wire             fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register_in;
  wire             fir_dma_read_master_requests_ext_ssram_s1;
  wire             fir_dma_read_master_saved_grant_ext_ssram_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 31: 0] incoming_ext_ssram_bus_data /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  reg              last_cycle_custom_dma_burst_0_downstream_granted_slave_ext_ssram_s1;
  reg              last_cycle_fir_dma_read_master_granted_slave_ext_ssram_s1;
  wire    [ 31: 0] outgoing_ext_ssram_bus_data;
  reg              outputenable_n_to_the_ext_ssram /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             p1_adsc_n_to_the_ext_ssram;
  wire    [  3: 0] p1_bw_n_to_the_ext_ssram;
  wire             p1_bwe_n_to_the_ext_ssram;
  wire             p1_chipenable1_n_to_the_ext_ssram;
  wire    [  3: 0] p1_custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register;
  wire    [ 20: 0] p1_ext_ssram_bus_address;
  wire    [  3: 0] p1_fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register;
  wire             p1_outputenable_n_to_the_ext_ssram;
  wire             time_to_write;
  wire             wait_for_ext_ssram_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~ext_ssram_bus_avalon_slave_end_xfer;
    end


  assign ext_ssram_bus_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 | fir_dma_read_master_qualified_request_ext_ssram_s1));
  assign custom_dma_burst_0_downstream_requests_ext_ssram_s1 = (1) & (custom_dma_burst_0_downstream_read | custom_dma_burst_0_downstream_write);
  //~chipenable1_n_to_the_ext_ssram of type chipselect to ~p1_chipenable1_n_to_the_ext_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          chipenable1_n_to_the_ext_ssram <= ~0;
      else 
        chipenable1_n_to_the_ext_ssram <= p1_chipenable1_n_to_the_ext_ssram;
    end


  assign ext_ssram_bus_avalon_slave_write_pending = 0;
  //ext_ssram_bus/avalon_slave read pending calc, which is an e_assign
  assign ext_ssram_bus_avalon_slave_read_pending = (|custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | (|fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[1 : 0]);

  //ext_ssram_bus_avalon_slave_arb_share_counter set values, which is an e_mux
  assign ext_ssram_bus_avalon_slave_arb_share_set_values = (custom_dma_burst_0_downstream_granted_ext_ssram_s1)? custom_dma_burst_0_downstream_arbitrationshare :
    (custom_dma_burst_0_downstream_granted_ext_ssram_s1)? custom_dma_burst_0_downstream_arbitrationshare :
    1;

  //ext_ssram_bus_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign ext_ssram_bus_avalon_slave_non_bursting_master_requests = 0 |
    fir_dma_read_master_requests_ext_ssram_s1 |
    fir_dma_read_master_requests_ext_ssram_s1;

  //ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant = custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1 |
    custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1;

  //ext_ssram_bus_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign ext_ssram_bus_avalon_slave_arb_share_counter_next_value = ext_ssram_bus_avalon_slave_firsttransfer ? (ext_ssram_bus_avalon_slave_arb_share_set_values - 1) : |ext_ssram_bus_avalon_slave_arb_share_counter ? (ext_ssram_bus_avalon_slave_arb_share_counter - 1) : 0;

  //ext_ssram_bus_avalon_slave_allgrants all slave grants, which is an e_mux
  assign ext_ssram_bus_avalon_slave_allgrants = (|ext_ssram_bus_avalon_slave_grant_vector) |
    (|ext_ssram_bus_avalon_slave_grant_vector) |
    (|ext_ssram_bus_avalon_slave_grant_vector) |
    (|ext_ssram_bus_avalon_slave_grant_vector);

  //ext_ssram_bus_avalon_slave_end_xfer assignment, which is an e_assign
  assign ext_ssram_bus_avalon_slave_end_xfer = ~(ext_ssram_s1_waits_for_read | ext_ssram_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave = ext_ssram_bus_avalon_slave_end_xfer & (~ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //ext_ssram_bus_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign ext_ssram_bus_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave & ext_ssram_bus_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave & ~ext_ssram_bus_avalon_slave_non_bursting_master_requests);

  //ext_ssram_bus_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_avalon_slave_arb_share_counter <= 0;
      else if (ext_ssram_bus_avalon_slave_arb_counter_enable)
          ext_ssram_bus_avalon_slave_arb_share_counter <= ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
    end


  //ext_ssram_bus_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|ext_ssram_bus_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave) | (end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave & ~ext_ssram_bus_avalon_slave_non_bursting_master_requests))
          ext_ssram_bus_avalon_slave_slavearbiterlockenable <= |ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
    end


  //custom_dma_burst_0/downstream ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  assign custom_dma_burst_0_downstream_arbiterlock = ext_ssram_bus_avalon_slave_slavearbiterlockenable & custom_dma_burst_0_downstream_continuerequest;

  //ext_ssram_bus_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign ext_ssram_bus_avalon_slave_slavearbiterlockenable2 = |ext_ssram_bus_avalon_slave_arb_share_counter_next_value;

  //custom_dma_burst_0/downstream ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign custom_dma_burst_0_downstream_arbiterlock2 = ext_ssram_bus_avalon_slave_slavearbiterlockenable2 & custom_dma_burst_0_downstream_continuerequest;

  //fir_dma/read_master ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  assign fir_dma_read_master_arbiterlock = ext_ssram_bus_avalon_slave_slavearbiterlockenable & fir_dma_read_master_continuerequest;

  //fir_dma/read_master ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  assign fir_dma_read_master_arbiterlock2 = ext_ssram_bus_avalon_slave_slavearbiterlockenable2 & fir_dma_read_master_continuerequest;

  //fir_dma/read_master granted ext_ssram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_fir_dma_read_master_granted_slave_ext_ssram_s1 <= 0;
      else 
        last_cycle_fir_dma_read_master_granted_slave_ext_ssram_s1 <= fir_dma_read_master_saved_grant_ext_ssram_s1 ? 1 : (ext_ssram_bus_avalon_slave_arbitration_holdoff_internal | 0) ? 0 : last_cycle_fir_dma_read_master_granted_slave_ext_ssram_s1;
    end


  //fir_dma_read_master_continuerequest continued request, which is an e_mux
  assign fir_dma_read_master_continuerequest = last_cycle_fir_dma_read_master_granted_slave_ext_ssram_s1 & fir_dma_read_master_requests_ext_ssram_s1;

  //ext_ssram_bus_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign ext_ssram_bus_avalon_slave_any_continuerequest = fir_dma_read_master_continuerequest |
    custom_dma_burst_0_downstream_continuerequest;

  assign custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 = custom_dma_burst_0_downstream_requests_ext_ssram_s1 & ~((custom_dma_burst_0_downstream_read & (ext_ssram_bus_avalon_slave_write_pending | (ext_ssram_bus_avalon_slave_read_pending & !((((|custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | (|fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[1 : 0]))))))) | ((ext_ssram_bus_avalon_slave_read_pending) & custom_dma_burst_0_downstream_write) | fir_dma_read_master_arbiterlock);
  //custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register_in = custom_dma_burst_0_downstream_granted_ext_ssram_s1 & custom_dma_burst_0_downstream_read & ~ext_ssram_s1_waits_for_read;

  //shift register p1 custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register = {custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register, custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register_in};

  //custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register <= 0;
      else 
        custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register <= p1_custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register;
    end


  //local readdatavalid custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1, which is an e_mux
  assign custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1 = custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[3];

  //ext_ssram_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_ext_ssram_bus_data <= 0;
      else 
        incoming_ext_ssram_bus_data <= ext_ssram_bus_data;
    end


  //ext_ssram_s1_with_write_latency assignment, which is an e_assign
  assign ext_ssram_s1_with_write_latency = in_a_write_cycle & (custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 | fir_dma_read_master_qualified_request_ext_ssram_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (ext_ssram_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_ext_ssram_bus_data register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_ext_ssram_bus_data <= 0;
      else 
        d1_outgoing_ext_ssram_bus_data <= outgoing_ext_ssram_bus_data;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_ext_ssram_bus_data tristate driver, which is an e_assign
  assign ext_ssram_bus_data = (d1_in_a_write_cycle)? d1_outgoing_ext_ssram_bus_data:{32{1'bz}};

  //outgoing_ext_ssram_bus_data mux, which is an e_mux
  assign outgoing_ext_ssram_bus_data = custom_dma_burst_0_downstream_writedata;

  assign fir_dma_read_master_requests_ext_ssram_s1 = (({fir_dma_read_master_address_to_slave[31 : 21] , 21'b0} == 32'h6000000) & (fir_dma_read_master_read)) & fir_dma_read_master_read;
  //custom_dma_burst_0/downstream granted ext_ssram/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_0_downstream_granted_slave_ext_ssram_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_0_downstream_granted_slave_ext_ssram_s1 <= custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1 ? 1 : (ext_ssram_bus_avalon_slave_arbitration_holdoff_internal | ~custom_dma_burst_0_downstream_requests_ext_ssram_s1) ? 0 : last_cycle_custom_dma_burst_0_downstream_granted_slave_ext_ssram_s1;
    end


  //custom_dma_burst_0_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_0_downstream_continuerequest = last_cycle_custom_dma_burst_0_downstream_granted_slave_ext_ssram_s1 & 1;

  assign fir_dma_read_master_qualified_request_ext_ssram_s1 = fir_dma_read_master_requests_ext_ssram_s1 & ~((fir_dma_read_master_read & (ext_ssram_bus_avalon_slave_write_pending | (ext_ssram_bus_avalon_slave_read_pending & !((((|custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | (|fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[1 : 0]))))))) | custom_dma_burst_0_downstream_arbiterlock);
  //fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register_in = fir_dma_read_master_granted_ext_ssram_s1 & fir_dma_read_master_read & ~ext_ssram_s1_waits_for_read;

  //shift register p1 fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register = {fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register, fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register_in};

  //fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register <= 0;
      else 
        fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register <= p1_fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register;
    end


  //local readdatavalid fir_dma_read_master_read_data_valid_ext_ssram_s1, which is an e_mux
  assign fir_dma_read_master_read_data_valid_ext_ssram_s1 = fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[3];

  //allow new arb cycle for ext_ssram_bus/avalon_slave, which is an e_assign
  assign ext_ssram_bus_avalon_slave_allow_new_arb_cycle = ~custom_dma_burst_0_downstream_arbiterlock & ~fir_dma_read_master_arbiterlock;

  //fir_dma/read_master assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  assign ext_ssram_bus_avalon_slave_master_qreq_vector[0] = fir_dma_read_master_qualified_request_ext_ssram_s1;

  //fir_dma/read_master grant ext_ssram/s1, which is an e_assign
  assign fir_dma_read_master_granted_ext_ssram_s1 = ext_ssram_bus_avalon_slave_grant_vector[0];

  //fir_dma/read_master saved-grant ext_ssram/s1, which is an e_assign
  assign fir_dma_read_master_saved_grant_ext_ssram_s1 = ext_ssram_bus_avalon_slave_arb_winner[0] && fir_dma_read_master_requests_ext_ssram_s1;

  //custom_dma_burst_0/downstream assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  assign ext_ssram_bus_avalon_slave_master_qreq_vector[1] = custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1;

  //custom_dma_burst_0/downstream grant ext_ssram/s1, which is an e_assign
  assign custom_dma_burst_0_downstream_granted_ext_ssram_s1 = ext_ssram_bus_avalon_slave_grant_vector[1];

  //custom_dma_burst_0/downstream saved-grant ext_ssram/s1, which is an e_assign
  assign custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1 = ext_ssram_bus_avalon_slave_arb_winner[1];

  //ext_ssram_bus/avalon_slave chosen-master double-vector, which is an e_assign
  assign ext_ssram_bus_avalon_slave_chosen_master_double_vector = {ext_ssram_bus_avalon_slave_master_qreq_vector, ext_ssram_bus_avalon_slave_master_qreq_vector} & ({~ext_ssram_bus_avalon_slave_master_qreq_vector, ~ext_ssram_bus_avalon_slave_master_qreq_vector} + ext_ssram_bus_avalon_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign ext_ssram_bus_avalon_slave_arb_winner = (ext_ssram_bus_avalon_slave_allow_new_arb_cycle & | ext_ssram_bus_avalon_slave_grant_vector) ? ext_ssram_bus_avalon_slave_grant_vector : ext_ssram_bus_avalon_slave_saved_chosen_master_vector;

  //saved ext_ssram_bus_avalon_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_avalon_slave_saved_chosen_master_vector <= 0;
      else if (ext_ssram_bus_avalon_slave_allow_new_arb_cycle)
          ext_ssram_bus_avalon_slave_saved_chosen_master_vector <= |ext_ssram_bus_avalon_slave_grant_vector ? ext_ssram_bus_avalon_slave_grant_vector : ext_ssram_bus_avalon_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign ext_ssram_bus_avalon_slave_grant_vector = {(ext_ssram_bus_avalon_slave_chosen_master_double_vector[1] | ext_ssram_bus_avalon_slave_chosen_master_double_vector[3]),
    (ext_ssram_bus_avalon_slave_chosen_master_double_vector[0] | ext_ssram_bus_avalon_slave_chosen_master_double_vector[2])};

  //ext_ssram_bus/avalon_slave chosen master rotated left, which is an e_assign
  assign ext_ssram_bus_avalon_slave_chosen_master_rot_left = (ext_ssram_bus_avalon_slave_arb_winner << 1) ? (ext_ssram_bus_avalon_slave_arb_winner << 1) : 1;

  //ext_ssram_bus/avalon_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_avalon_slave_arb_addend <= 1;
      else if (|ext_ssram_bus_avalon_slave_grant_vector)
          ext_ssram_bus_avalon_slave_arb_addend <= ext_ssram_bus_avalon_slave_end_xfer? ext_ssram_bus_avalon_slave_chosen_master_rot_left : ext_ssram_bus_avalon_slave_grant_vector;
    end


  //~adsc_n_to_the_ext_ssram of type begintransfer to ~p1_adsc_n_to_the_ext_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          adsc_n_to_the_ext_ssram <= ~0;
      else 
        adsc_n_to_the_ext_ssram <= p1_adsc_n_to_the_ext_ssram;
    end


  assign p1_adsc_n_to_the_ext_ssram = ~ext_ssram_bus_avalon_slave_begins_xfer;
  //~outputenable_n_to_the_ext_ssram of type outputenable to ~p1_outputenable_n_to_the_ext_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          outputenable_n_to_the_ext_ssram <= ~0;
      else 
        outputenable_n_to_the_ext_ssram <= p1_outputenable_n_to_the_ext_ssram;
    end


  //~p1_outputenable_n_to_the_ext_ssram assignment, which is an e_mux
  assign p1_outputenable_n_to_the_ext_ssram = ~((|custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | (|fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | ext_ssram_s1_in_a_read_cycle);

  assign p1_chipenable1_n_to_the_ext_ssram = ~(custom_dma_burst_0_downstream_granted_ext_ssram_s1 | fir_dma_read_master_granted_ext_ssram_s1 | (|custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1_shift_register[1 : 0]) | (|fir_dma_read_master_read_data_valid_ext_ssram_s1_shift_register[1 : 0]));
  //ext_ssram_bus_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign ext_ssram_bus_avalon_slave_firsttransfer = ext_ssram_bus_avalon_slave_begins_xfer ? ext_ssram_bus_avalon_slave_unreg_firsttransfer : ext_ssram_bus_avalon_slave_reg_firsttransfer;

  //ext_ssram_bus_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign ext_ssram_bus_avalon_slave_unreg_firsttransfer = ~(ext_ssram_bus_avalon_slave_slavearbiterlockenable & ext_ssram_bus_avalon_slave_any_continuerequest);

  //ext_ssram_bus_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (ext_ssram_bus_avalon_slave_begins_xfer)
          ext_ssram_bus_avalon_slave_reg_firsttransfer <= ext_ssram_bus_avalon_slave_unreg_firsttransfer;
    end


  //ext_ssram_bus_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign ext_ssram_bus_avalon_slave_beginbursttransfer_internal = ext_ssram_bus_avalon_slave_begins_xfer;

  //ext_ssram_bus_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign ext_ssram_bus_avalon_slave_arbitration_holdoff_internal = ext_ssram_bus_avalon_slave_begins_xfer & ext_ssram_bus_avalon_slave_firsttransfer;

  //~bwe_n_to_the_ext_ssram of type write to ~p1_bwe_n_to_the_ext_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          bwe_n_to_the_ext_ssram <= ~0;
      else 
        bwe_n_to_the_ext_ssram <= p1_bwe_n_to_the_ext_ssram;
    end


  //~bw_n_to_the_ext_ssram of type byteenable to ~p1_bw_n_to_the_ext_ssram, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          bw_n_to_the_ext_ssram <= ~0;
      else 
        bw_n_to_the_ext_ssram <= p1_bw_n_to_the_ext_ssram;
    end


  //~p1_bwe_n_to_the_ext_ssram assignment, which is an e_mux
  assign p1_bwe_n_to_the_ext_ssram = ~(custom_dma_burst_0_downstream_granted_ext_ssram_s1 & custom_dma_burst_0_downstream_write);

  //ext_ssram_bus_address of type address to p1_ext_ssram_bus_address, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          ext_ssram_bus_address <= 0;
      else 
        ext_ssram_bus_address <= p1_ext_ssram_bus_address;
    end


  //p1_ext_ssram_bus_address mux, which is an e_mux
  assign p1_ext_ssram_bus_address = (custom_dma_burst_0_downstream_granted_ext_ssram_s1)? custom_dma_burst_0_downstream_address_to_slave :
    fir_dma_read_master_address_to_slave;

  //d1_ext_ssram_bus_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_ext_ssram_bus_avalon_slave_end_xfer <= 1;
      else 
        d1_ext_ssram_bus_avalon_slave_end_xfer <= ext_ssram_bus_avalon_slave_end_xfer;
    end


  //ext_ssram_s1_waits_for_read in a cycle, which is an e_mux
  assign ext_ssram_s1_waits_for_read = ext_ssram_s1_in_a_read_cycle & 0;

  //ext_ssram_s1_in_a_read_cycle assignment, which is an e_assign
  assign ext_ssram_s1_in_a_read_cycle = (custom_dma_burst_0_downstream_granted_ext_ssram_s1 & custom_dma_burst_0_downstream_read) | (fir_dma_read_master_granted_ext_ssram_s1 & fir_dma_read_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = ext_ssram_s1_in_a_read_cycle;

  //ext_ssram_s1_waits_for_write in a cycle, which is an e_mux
  assign ext_ssram_s1_waits_for_write = ext_ssram_s1_in_a_write_cycle & 0;

  //ext_ssram_s1_in_a_write_cycle assignment, which is an e_assign
  assign ext_ssram_s1_in_a_write_cycle = custom_dma_burst_0_downstream_granted_ext_ssram_s1 & custom_dma_burst_0_downstream_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = ext_ssram_s1_in_a_write_cycle;

  assign wait_for_ext_ssram_s1_counter = 0;
  //~p1_bw_n_to_the_ext_ssram byte enable port mux, which is an e_mux
  assign p1_bw_n_to_the_ext_ssram = ~((custom_dma_burst_0_downstream_granted_ext_ssram_s1)? custom_dma_burst_0_downstream_byteenable :
    -1);


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //ext_ssram/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //custom_dma_burst_0/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_0_downstream_requests_ext_ssram_s1 && (custom_dma_burst_0_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_0/downstream drove 0 on its 'arbitrationshare' port while accessing slave ext_ssram/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_0/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_0_downstream_requests_ext_ssram_s1 && (custom_dma_burst_0_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_0/downstream drove 0 on its 'burstcount' port while accessing slave ext_ssram/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_0_downstream_granted_ext_ssram_s1 + fir_dma_read_master_granted_ext_ssram_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_0_downstream_saved_grant_ext_ssram_s1 + fir_dma_read_master_saved_grant_ext_ssram_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_bus_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module fir_dma_control_arbitrator (
                                    // inputs:
                                     clk,
                                     fir_dma_control_irq,
                                     fir_dma_control_readdata,
                                     pipeline_bridge_m1_address_to_slave,
                                     pipeline_bridge_m1_burstcount,
                                     pipeline_bridge_m1_byteenable,
                                     pipeline_bridge_m1_chipselect,
                                     pipeline_bridge_m1_latency_counter,
                                     pipeline_bridge_m1_read,
                                     pipeline_bridge_m1_write,
                                     pipeline_bridge_m1_writedata,
                                     reset_n,

                                    // outputs:
                                     d1_fir_dma_control_end_xfer,
                                     fir_dma_control_address,
                                     fir_dma_control_byteenable,
                                     fir_dma_control_irq_from_sa,
                                     fir_dma_control_read,
                                     fir_dma_control_readdata_from_sa,
                                     fir_dma_control_reset,
                                     fir_dma_control_write,
                                     fir_dma_control_writedata,
                                     pipeline_bridge_m1_granted_fir_dma_control,
                                     pipeline_bridge_m1_qualified_request_fir_dma_control,
                                     pipeline_bridge_m1_read_data_valid_fir_dma_control,
                                     pipeline_bridge_m1_requests_fir_dma_control
                                  )
;

  output           d1_fir_dma_control_end_xfer;
  output  [  2: 0] fir_dma_control_address;
  output  [  3: 0] fir_dma_control_byteenable;
  output           fir_dma_control_irq_from_sa;
  output           fir_dma_control_read;
  output  [ 31: 0] fir_dma_control_readdata_from_sa;
  output           fir_dma_control_reset;
  output           fir_dma_control_write;
  output  [ 31: 0] fir_dma_control_writedata;
  output           pipeline_bridge_m1_granted_fir_dma_control;
  output           pipeline_bridge_m1_qualified_request_fir_dma_control;
  output           pipeline_bridge_m1_read_data_valid_fir_dma_control;
  output           pipeline_bridge_m1_requests_fir_dma_control;
  input            clk;
  input            fir_dma_control_irq;
  input   [ 31: 0] fir_dma_control_readdata;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_fir_dma_control_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_fir_dma_control;
  wire    [  2: 0] fir_dma_control_address;
  wire             fir_dma_control_allgrants;
  wire             fir_dma_control_allow_new_arb_cycle;
  wire             fir_dma_control_any_bursting_master_saved_grant;
  wire             fir_dma_control_any_continuerequest;
  wire             fir_dma_control_arb_counter_enable;
  reg              fir_dma_control_arb_share_counter;
  wire             fir_dma_control_arb_share_counter_next_value;
  wire             fir_dma_control_arb_share_set_values;
  wire             fir_dma_control_beginbursttransfer_internal;
  wire             fir_dma_control_begins_xfer;
  wire    [  3: 0] fir_dma_control_byteenable;
  wire             fir_dma_control_end_xfer;
  wire             fir_dma_control_firsttransfer;
  wire             fir_dma_control_grant_vector;
  wire             fir_dma_control_in_a_read_cycle;
  wire             fir_dma_control_in_a_write_cycle;
  wire             fir_dma_control_irq_from_sa;
  wire             fir_dma_control_master_qreq_vector;
  wire             fir_dma_control_non_bursting_master_requests;
  wire             fir_dma_control_read;
  wire    [ 31: 0] fir_dma_control_readdata_from_sa;
  reg              fir_dma_control_reg_firsttransfer;
  wire             fir_dma_control_reset;
  reg              fir_dma_control_slavearbiterlockenable;
  wire             fir_dma_control_slavearbiterlockenable2;
  wire             fir_dma_control_unreg_firsttransfer;
  wire             fir_dma_control_waits_for_read;
  wire             fir_dma_control_waits_for_write;
  wire             fir_dma_control_write;
  wire    [ 31: 0] fir_dma_control_writedata;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             p1_pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_fir_dma_control;
  wire             pipeline_bridge_m1_qualified_request_fir_dma_control;
  wire             pipeline_bridge_m1_read_data_valid_fir_dma_control;
  reg              pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register;
  wire             pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register_in;
  wire             pipeline_bridge_m1_requests_fir_dma_control;
  wire             pipeline_bridge_m1_saved_grant_fir_dma_control;
  wire    [ 11: 0] shifted_address_to_fir_dma_control_from_pipeline_bridge_m1;
  wire             wait_for_fir_dma_control_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~fir_dma_control_end_xfer;
    end


  assign fir_dma_control_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_fir_dma_control));
  //assign fir_dma_control_readdata_from_sa = fir_dma_control_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign fir_dma_control_readdata_from_sa = fir_dma_control_readdata;

  assign pipeline_bridge_m1_requests_fir_dma_control = ({pipeline_bridge_m1_address_to_slave[11 : 5] , 5'b0} == 12'h840) & pipeline_bridge_m1_chipselect;
  //fir_dma_control_arb_share_counter set values, which is an e_mux
  assign fir_dma_control_arb_share_set_values = 1;

  //fir_dma_control_non_bursting_master_requests mux, which is an e_mux
  assign fir_dma_control_non_bursting_master_requests = pipeline_bridge_m1_requests_fir_dma_control;

  //fir_dma_control_any_bursting_master_saved_grant mux, which is an e_mux
  assign fir_dma_control_any_bursting_master_saved_grant = 0;

  //fir_dma_control_arb_share_counter_next_value assignment, which is an e_assign
  assign fir_dma_control_arb_share_counter_next_value = fir_dma_control_firsttransfer ? (fir_dma_control_arb_share_set_values - 1) : |fir_dma_control_arb_share_counter ? (fir_dma_control_arb_share_counter - 1) : 0;

  //fir_dma_control_allgrants all slave grants, which is an e_mux
  assign fir_dma_control_allgrants = |fir_dma_control_grant_vector;

  //fir_dma_control_end_xfer assignment, which is an e_assign
  assign fir_dma_control_end_xfer = ~(fir_dma_control_waits_for_read | fir_dma_control_waits_for_write);

  //end_xfer_arb_share_counter_term_fir_dma_control arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_fir_dma_control = fir_dma_control_end_xfer & (~fir_dma_control_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //fir_dma_control_arb_share_counter arbitration counter enable, which is an e_assign
  assign fir_dma_control_arb_counter_enable = (end_xfer_arb_share_counter_term_fir_dma_control & fir_dma_control_allgrants) | (end_xfer_arb_share_counter_term_fir_dma_control & ~fir_dma_control_non_bursting_master_requests);

  //fir_dma_control_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_control_arb_share_counter <= 0;
      else if (fir_dma_control_arb_counter_enable)
          fir_dma_control_arb_share_counter <= fir_dma_control_arb_share_counter_next_value;
    end


  //fir_dma_control_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_control_slavearbiterlockenable <= 0;
      else if ((|fir_dma_control_master_qreq_vector & end_xfer_arb_share_counter_term_fir_dma_control) | (end_xfer_arb_share_counter_term_fir_dma_control & ~fir_dma_control_non_bursting_master_requests))
          fir_dma_control_slavearbiterlockenable <= |fir_dma_control_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 fir_dma/control arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = fir_dma_control_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //fir_dma_control_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign fir_dma_control_slavearbiterlockenable2 = |fir_dma_control_arb_share_counter_next_value;

  //pipeline_bridge/m1 fir_dma/control arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = fir_dma_control_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //fir_dma_control_any_continuerequest at least one master continues requesting, which is an e_assign
  assign fir_dma_control_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_fir_dma_control = pipeline_bridge_m1_requests_fir_dma_control & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((1 < pipeline_bridge_m1_latency_counter))));
  //pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register_in mux for readlatency shift register, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register_in = pipeline_bridge_m1_granted_fir_dma_control & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~fir_dma_control_waits_for_read;

  //shift register p1 pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register = {pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register, pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register_in};

  //pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register <= 0;
      else 
        pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register <= p1_pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register;
    end


  //local readdatavalid pipeline_bridge_m1_read_data_valid_fir_dma_control, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_fir_dma_control = pipeline_bridge_m1_read_data_valid_fir_dma_control_shift_register;

  //fir_dma_control_writedata mux, which is an e_mux
  assign fir_dma_control_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_fir_dma_control = pipeline_bridge_m1_qualified_request_fir_dma_control;

  //pipeline_bridge/m1 saved-grant fir_dma/control, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_fir_dma_control = pipeline_bridge_m1_requests_fir_dma_control;

  //allow new arb cycle for fir_dma/control, which is an e_assign
  assign fir_dma_control_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign fir_dma_control_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign fir_dma_control_master_qreq_vector = 1;

  //~fir_dma_control_reset assignment, which is an e_assign
  assign fir_dma_control_reset = ~reset_n;

  //fir_dma_control_firsttransfer first transaction, which is an e_assign
  assign fir_dma_control_firsttransfer = fir_dma_control_begins_xfer ? fir_dma_control_unreg_firsttransfer : fir_dma_control_reg_firsttransfer;

  //fir_dma_control_unreg_firsttransfer first transaction, which is an e_assign
  assign fir_dma_control_unreg_firsttransfer = ~(fir_dma_control_slavearbiterlockenable & fir_dma_control_any_continuerequest);

  //fir_dma_control_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_control_reg_firsttransfer <= 1'b1;
      else if (fir_dma_control_begins_xfer)
          fir_dma_control_reg_firsttransfer <= fir_dma_control_unreg_firsttransfer;
    end


  //fir_dma_control_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign fir_dma_control_beginbursttransfer_internal = fir_dma_control_begins_xfer;

  //fir_dma_control_read assignment, which is an e_mux
  assign fir_dma_control_read = pipeline_bridge_m1_granted_fir_dma_control & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //fir_dma_control_write assignment, which is an e_mux
  assign fir_dma_control_write = pipeline_bridge_m1_granted_fir_dma_control & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  assign shifted_address_to_fir_dma_control_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //fir_dma_control_address mux, which is an e_mux
  assign fir_dma_control_address = shifted_address_to_fir_dma_control_from_pipeline_bridge_m1 >> 2;

  //d1_fir_dma_control_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_fir_dma_control_end_xfer <= 1;
      else 
        d1_fir_dma_control_end_xfer <= fir_dma_control_end_xfer;
    end


  //fir_dma_control_waits_for_read in a cycle, which is an e_mux
  assign fir_dma_control_waits_for_read = fir_dma_control_in_a_read_cycle & 0;

  //fir_dma_control_in_a_read_cycle assignment, which is an e_assign
  assign fir_dma_control_in_a_read_cycle = pipeline_bridge_m1_granted_fir_dma_control & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = fir_dma_control_in_a_read_cycle;

  //fir_dma_control_waits_for_write in a cycle, which is an e_mux
  assign fir_dma_control_waits_for_write = fir_dma_control_in_a_write_cycle & 0;

  //fir_dma_control_in_a_write_cycle assignment, which is an e_assign
  assign fir_dma_control_in_a_write_cycle = pipeline_bridge_m1_granted_fir_dma_control & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = fir_dma_control_in_a_write_cycle;

  assign wait_for_fir_dma_control_counter = 0;
  //fir_dma_control_byteenable byte enable port mux, which is an e_mux
  assign fir_dma_control_byteenable = (pipeline_bridge_m1_granted_fir_dma_control)? pipeline_bridge_m1_byteenable :
    -1;

  //assign fir_dma_control_irq_from_sa = fir_dma_control_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign fir_dma_control_irq_from_sa = fir_dma_control_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //fir_dma/control enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_fir_dma_control && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave fir_dma/control", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module fir_dma_read_master_arbitrator (
                                        // inputs:
                                         clk,
                                         d1_ext_ssram_bus_avalon_slave_end_xfer,
                                         fir_dma_read_master_address,
                                         fir_dma_read_master_byteenable,
                                         fir_dma_read_master_granted_ext_ssram_s1,
                                         fir_dma_read_master_qualified_request_ext_ssram_s1,
                                         fir_dma_read_master_read,
                                         fir_dma_read_master_read_data_valid_ext_ssram_s1,
                                         fir_dma_read_master_requests_ext_ssram_s1,
                                         incoming_ext_ssram_bus_data,
                                         reset_n,

                                        // outputs:
                                         fir_dma_read_master_address_to_slave,
                                         fir_dma_read_master_latency_counter,
                                         fir_dma_read_master_readdata,
                                         fir_dma_read_master_readdatavalid,
                                         fir_dma_read_master_waitrequest
                                      )
;

  output  [ 31: 0] fir_dma_read_master_address_to_slave;
  output  [  2: 0] fir_dma_read_master_latency_counter;
  output  [ 31: 0] fir_dma_read_master_readdata;
  output           fir_dma_read_master_readdatavalid;
  output           fir_dma_read_master_waitrequest;
  input            clk;
  input            d1_ext_ssram_bus_avalon_slave_end_xfer;
  input   [ 31: 0] fir_dma_read_master_address;
  input   [  3: 0] fir_dma_read_master_byteenable;
  input            fir_dma_read_master_granted_ext_ssram_s1;
  input            fir_dma_read_master_qualified_request_ext_ssram_s1;
  input            fir_dma_read_master_read;
  input            fir_dma_read_master_read_data_valid_ext_ssram_s1;
  input            fir_dma_read_master_requests_ext_ssram_s1;
  input   [ 31: 0] incoming_ext_ssram_bus_data;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] fir_dma_read_master_address_last_time;
  wire    [ 31: 0] fir_dma_read_master_address_to_slave;
  reg     [  3: 0] fir_dma_read_master_byteenable_last_time;
  wire             fir_dma_read_master_is_granted_some_slave;
  reg     [  2: 0] fir_dma_read_master_latency_counter;
  reg              fir_dma_read_master_read_but_no_slave_selected;
  reg              fir_dma_read_master_read_last_time;
  wire    [ 31: 0] fir_dma_read_master_readdata;
  wire             fir_dma_read_master_readdatavalid;
  wire             fir_dma_read_master_run;
  wire             fir_dma_read_master_waitrequest;
  wire    [  2: 0] latency_load_value;
  wire    [  2: 0] p1_fir_dma_read_master_latency_counter;
  wire             pre_flush_fir_dma_read_master_readdatavalid;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (fir_dma_read_master_qualified_request_ext_ssram_s1 | ~fir_dma_read_master_requests_ext_ssram_s1) & (fir_dma_read_master_granted_ext_ssram_s1 | ~fir_dma_read_master_qualified_request_ext_ssram_s1) & ((~fir_dma_read_master_qualified_request_ext_ssram_s1 | ~(fir_dma_read_master_read) | (1 & (fir_dma_read_master_read))));

  //cascaded wait assignment, which is an e_assign
  assign fir_dma_read_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign fir_dma_read_master_address_to_slave = {11'b110000,
    fir_dma_read_master_address[20 : 0]};

  //fir_dma_read_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_read_but_no_slave_selected <= 0;
      else 
        fir_dma_read_master_read_but_no_slave_selected <= fir_dma_read_master_read & fir_dma_read_master_run & ~fir_dma_read_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign fir_dma_read_master_is_granted_some_slave = fir_dma_read_master_granted_ext_ssram_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_fir_dma_read_master_readdatavalid = fir_dma_read_master_read_data_valid_ext_ssram_s1;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign fir_dma_read_master_readdatavalid = fir_dma_read_master_read_but_no_slave_selected |
    pre_flush_fir_dma_read_master_readdatavalid;

  //fir_dma/read_master readdata mux, which is an e_mux
  assign fir_dma_read_master_readdata = incoming_ext_ssram_bus_data;

  //actual waitrequest port, which is an e_assign
  assign fir_dma_read_master_waitrequest = ~fir_dma_read_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_latency_counter <= 0;
      else 
        fir_dma_read_master_latency_counter <= p1_fir_dma_read_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_fir_dma_read_master_latency_counter = ((fir_dma_read_master_run & fir_dma_read_master_read))? latency_load_value :
    (fir_dma_read_master_latency_counter)? fir_dma_read_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {3 {fir_dma_read_master_requests_ext_ssram_s1}} & 4;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //fir_dma_read_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_address_last_time <= 0;
      else 
        fir_dma_read_master_address_last_time <= fir_dma_read_master_address;
    end


  //fir_dma/read_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= fir_dma_read_master_waitrequest & (fir_dma_read_master_read);
    end


  //fir_dma_read_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_read_master_address != fir_dma_read_master_address_last_time))
        begin
          $write("%0d ns: fir_dma_read_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_read_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_byteenable_last_time <= 0;
      else 
        fir_dma_read_master_byteenable_last_time <= fir_dma_read_master_byteenable;
    end


  //fir_dma_read_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_read_master_byteenable != fir_dma_read_master_byteenable_last_time))
        begin
          $write("%0d ns: fir_dma_read_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_read_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_read_master_read_last_time <= 0;
      else 
        fir_dma_read_master_read_last_time <= fir_dma_read_master_read;
    end


  //fir_dma_read_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_read_master_read != fir_dma_read_master_read_last_time))
        begin
          $write("%0d ns: fir_dma_read_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module fir_dma_write_master_arbitrator (
                                         // inputs:
                                          clk,
                                          custom_dma_burst_5_upstream_waitrequest_from_sa,
                                          d1_custom_dma_burst_5_upstream_end_xfer,
                                          fir_dma_write_master_address,
                                          fir_dma_write_master_burstcount,
                                          fir_dma_write_master_byteenable,
                                          fir_dma_write_master_granted_custom_dma_burst_5_upstream,
                                          fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream,
                                          fir_dma_write_master_requests_custom_dma_burst_5_upstream,
                                          fir_dma_write_master_write,
                                          fir_dma_write_master_writedata,
                                          reset_n,

                                         // outputs:
                                          fir_dma_write_master_address_to_slave,
                                          fir_dma_write_master_waitrequest
                                       )
;

  output  [ 31: 0] fir_dma_write_master_address_to_slave;
  output           fir_dma_write_master_waitrequest;
  input            clk;
  input            custom_dma_burst_5_upstream_waitrequest_from_sa;
  input            d1_custom_dma_burst_5_upstream_end_xfer;
  input   [ 31: 0] fir_dma_write_master_address;
  input   [  2: 0] fir_dma_write_master_burstcount;
  input   [  3: 0] fir_dma_write_master_byteenable;
  input            fir_dma_write_master_granted_custom_dma_burst_5_upstream;
  input            fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream;
  input            fir_dma_write_master_requests_custom_dma_burst_5_upstream;
  input            fir_dma_write_master_write;
  input   [ 31: 0] fir_dma_write_master_writedata;
  input            reset_n;

  reg              active_and_waiting_last_time;
  reg     [ 31: 0] fir_dma_write_master_address_last_time;
  wire    [ 31: 0] fir_dma_write_master_address_to_slave;
  reg     [  2: 0] fir_dma_write_master_burstcount_last_time;
  reg     [  3: 0] fir_dma_write_master_byteenable_last_time;
  wire             fir_dma_write_master_run;
  wire             fir_dma_write_master_waitrequest;
  reg              fir_dma_write_master_write_last_time;
  reg     [ 31: 0] fir_dma_write_master_writedata_last_time;
  wire             r_0;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & ((~fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream | ~(fir_dma_write_master_write) | (1 & ~custom_dma_burst_5_upstream_waitrequest_from_sa & (fir_dma_write_master_write))));

  //cascaded wait assignment, which is an e_assign
  assign fir_dma_write_master_run = r_0;

  //optimize select-logic by passing only those address bits which matter.
  assign fir_dma_write_master_address_to_slave = {7'b1,
    fir_dma_write_master_address[24 : 0]};

  //actual waitrequest port, which is an e_assign
  assign fir_dma_write_master_waitrequest = ~fir_dma_write_master_run;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //fir_dma_write_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_write_master_address_last_time <= 0;
      else 
        fir_dma_write_master_address_last_time <= fir_dma_write_master_address;
    end


  //fir_dma/write_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= fir_dma_write_master_waitrequest & (fir_dma_write_master_write);
    end


  //fir_dma_write_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_write_master_address != fir_dma_write_master_address_last_time))
        begin
          $write("%0d ns: fir_dma_write_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_write_master_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_write_master_burstcount_last_time <= 0;
      else 
        fir_dma_write_master_burstcount_last_time <= fir_dma_write_master_burstcount;
    end


  //fir_dma_write_master_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_write_master_burstcount != fir_dma_write_master_burstcount_last_time))
        begin
          $write("%0d ns: fir_dma_write_master_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_write_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_write_master_byteenable_last_time <= 0;
      else 
        fir_dma_write_master_byteenable_last_time <= fir_dma_write_master_byteenable;
    end


  //fir_dma_write_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_write_master_byteenable != fir_dma_write_master_byteenable_last_time))
        begin
          $write("%0d ns: fir_dma_write_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_write_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_write_master_write_last_time <= 0;
      else 
        fir_dma_write_master_write_last_time <= fir_dma_write_master_write;
    end


  //fir_dma_write_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_write_master_write != fir_dma_write_master_write_last_time))
        begin
          $write("%0d ns: fir_dma_write_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //fir_dma_write_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fir_dma_write_master_writedata_last_time <= 0;
      else 
        fir_dma_write_master_writedata_last_time <= fir_dma_write_master_writedata;
    end


  //fir_dma_write_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (fir_dma_write_master_writedata != fir_dma_write_master_writedata_last_time) & fir_dma_write_master_write)
        begin
          $write("%0d ns: fir_dma_write_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_avalon_jtag_slave_arbitrator (
                                                // inputs:
                                                 clk,
                                                 jtag_uart_avalon_jtag_slave_dataavailable,
                                                 jtag_uart_avalon_jtag_slave_irq,
                                                 jtag_uart_avalon_jtag_slave_readdata,
                                                 jtag_uart_avalon_jtag_slave_readyfordata,
                                                 jtag_uart_avalon_jtag_slave_waitrequest,
                                                 pipeline_bridge_m1_address_to_slave,
                                                 pipeline_bridge_m1_burstcount,
                                                 pipeline_bridge_m1_chipselect,
                                                 pipeline_bridge_m1_latency_counter,
                                                 pipeline_bridge_m1_read,
                                                 pipeline_bridge_m1_write,
                                                 pipeline_bridge_m1_writedata,
                                                 reset_n,

                                                // outputs:
                                                 d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                                 jtag_uart_avalon_jtag_slave_address,
                                                 jtag_uart_avalon_jtag_slave_chipselect,
                                                 jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
                                                 jtag_uart_avalon_jtag_slave_irq_from_sa,
                                                 jtag_uart_avalon_jtag_slave_read_n,
                                                 jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
                                                 jtag_uart_avalon_jtag_slave_reset_n,
                                                 jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                                 jtag_uart_avalon_jtag_slave_write_n,
                                                 jtag_uart_avalon_jtag_slave_writedata,
                                                 pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                                 pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                                 pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                                 pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave
                                              )
;

  output           d1_jtag_uart_avalon_jtag_slave_end_xfer;
  output           jtag_uart_avalon_jtag_slave_address;
  output           jtag_uart_avalon_jtag_slave_chipselect;
  output           jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_avalon_jtag_slave_reset_n;
  output           jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  output           pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  output           pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  output           pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  output           pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  input            clk;
  input            jtag_uart_avalon_jtag_slave_dataavailable;
  input            jtag_uart_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  input            jtag_uart_avalon_jtag_slave_readyfordata;
  input            jtag_uart_avalon_jtag_slave_waitrequest;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;

  reg              d1_jtag_uart_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_allgrants;
  wire             jtag_uart_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_avalon_jtag_slave_arb_counter_enable;
  reg              jtag_uart_avalon_jtag_slave_arb_share_counter;
  wire             jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
  wire             jtag_uart_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  reg              jtag_uart_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave;
  wire    [ 11: 0] shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1;
  wire             wait_for_jtag_uart_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave));
  //assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata;

  assign pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave = ({pipeline_bridge_m1_address_to_slave[11 : 3] , 3'b0} == 12'h868) & pipeline_bridge_m1_chipselect;
  //assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest;

  //jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_non_bursting_master_requests = pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_avalon_jtag_slave_firsttransfer ? (jtag_uart_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_avalon_jtag_slave_arb_share_counter ? (jtag_uart_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_allgrants = |jtag_uart_avalon_jtag_slave_grant_vector;

  //jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_end_xfer = ~(jtag_uart_avalon_jtag_slave_waits_for_read | jtag_uart_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave = jtag_uart_avalon_jtag_slave_end_xfer & (~jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & jtag_uart_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave & ~jtag_uart_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = jtag_uart_avalon_jtag_slave_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;

  //pipeline_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave = pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave = pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~jtag_uart_avalon_jtag_slave_waits_for_read;

  //jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave = pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;

  //pipeline_bridge/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave = pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_avalon_jtag_slave_chipselect = pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  //jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_firsttransfer = jtag_uart_avalon_jtag_slave_begins_xfer ? jtag_uart_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_avalon_jtag_slave_begins_xfer)
          jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_read_n = ~(pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect));

  //~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_write_n = ~(pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect));

  assign shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_address = shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1 >> 2;

  //d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_read = jtag_uart_avalon_jtag_slave_in_a_read_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_read_cycle = pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_avalon_jtag_slave_waits_for_write = jtag_uart_avalon_jtag_slave_in_a_write_cycle & jtag_uart_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_in_a_write_cycle = pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_custom_dma_burst_1_downstream_to_pipeline_bridge_s1_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_custom_dma_burst_2_downstream_to_pipeline_bridge_s1_module (
                                                                                 // inputs:
                                                                                  clear_fifo,
                                                                                  clk,
                                                                                  data_in,
                                                                                  read,
                                                                                  reset_n,
                                                                                  sync_reset,
                                                                                  write,

                                                                                 // outputs:
                                                                                  data_out,
                                                                                  empty,
                                                                                  fifo_contains_ones_n,
                                                                                  full
                                                                               )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  wire             full_4;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_3;
  assign empty = !full_0;
  assign full_4 = 0;
  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    0;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_s1_arbitrator (
                                       // inputs:
                                        clk,
                                        custom_dma_burst_1_downstream_address_to_slave,
                                        custom_dma_burst_1_downstream_arbitrationshare,
                                        custom_dma_burst_1_downstream_burstcount,
                                        custom_dma_burst_1_downstream_byteenable,
                                        custom_dma_burst_1_downstream_debugaccess,
                                        custom_dma_burst_1_downstream_latency_counter,
                                        custom_dma_burst_1_downstream_nativeaddress,
                                        custom_dma_burst_1_downstream_read,
                                        custom_dma_burst_1_downstream_write,
                                        custom_dma_burst_1_downstream_writedata,
                                        custom_dma_burst_2_downstream_address_to_slave,
                                        custom_dma_burst_2_downstream_arbitrationshare,
                                        custom_dma_burst_2_downstream_burstcount,
                                        custom_dma_burst_2_downstream_byteenable,
                                        custom_dma_burst_2_downstream_debugaccess,
                                        custom_dma_burst_2_downstream_latency_counter,
                                        custom_dma_burst_2_downstream_nativeaddress,
                                        custom_dma_burst_2_downstream_read,
                                        custom_dma_burst_2_downstream_write,
                                        custom_dma_burst_2_downstream_writedata,
                                        pipeline_bridge_s1_endofpacket,
                                        pipeline_bridge_s1_readdata,
                                        pipeline_bridge_s1_readdatavalid,
                                        pipeline_bridge_s1_waitrequest,
                                        reset_n,

                                       // outputs:
                                        custom_dma_burst_1_downstream_granted_pipeline_bridge_s1,
                                        custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1,
                                        custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1,
                                        custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register,
                                        custom_dma_burst_1_downstream_requests_pipeline_bridge_s1,
                                        custom_dma_burst_2_downstream_granted_pipeline_bridge_s1,
                                        custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1,
                                        custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1,
                                        custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register,
                                        custom_dma_burst_2_downstream_requests_pipeline_bridge_s1,
                                        d1_pipeline_bridge_s1_end_xfer,
                                        pipeline_bridge_s1_address,
                                        pipeline_bridge_s1_arbiterlock,
                                        pipeline_bridge_s1_arbiterlock2,
                                        pipeline_bridge_s1_burstcount,
                                        pipeline_bridge_s1_byteenable,
                                        pipeline_bridge_s1_chipselect,
                                        pipeline_bridge_s1_debugaccess,
                                        pipeline_bridge_s1_endofpacket_from_sa,
                                        pipeline_bridge_s1_nativeaddress,
                                        pipeline_bridge_s1_read,
                                        pipeline_bridge_s1_readdata_from_sa,
                                        pipeline_bridge_s1_reset_n,
                                        pipeline_bridge_s1_waitrequest_from_sa,
                                        pipeline_bridge_s1_write,
                                        pipeline_bridge_s1_writedata
                                     )
;

  output           custom_dma_burst_1_downstream_granted_pipeline_bridge_s1;
  output           custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1;
  output           custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1;
  output           custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  output           custom_dma_burst_1_downstream_requests_pipeline_bridge_s1;
  output           custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;
  output           custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1;
  output           custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1;
  output           custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  output           custom_dma_burst_2_downstream_requests_pipeline_bridge_s1;
  output           d1_pipeline_bridge_s1_end_xfer;
  output  [  9: 0] pipeline_bridge_s1_address;
  output           pipeline_bridge_s1_arbiterlock;
  output           pipeline_bridge_s1_arbiterlock2;
  output           pipeline_bridge_s1_burstcount;
  output  [  3: 0] pipeline_bridge_s1_byteenable;
  output           pipeline_bridge_s1_chipselect;
  output           pipeline_bridge_s1_debugaccess;
  output           pipeline_bridge_s1_endofpacket_from_sa;
  output  [  9: 0] pipeline_bridge_s1_nativeaddress;
  output           pipeline_bridge_s1_read;
  output  [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  output           pipeline_bridge_s1_reset_n;
  output           pipeline_bridge_s1_waitrequest_from_sa;
  output           pipeline_bridge_s1_write;
  output  [ 31: 0] pipeline_bridge_s1_writedata;
  input            clk;
  input   [ 11: 0] custom_dma_burst_1_downstream_address_to_slave;
  input   [  3: 0] custom_dma_burst_1_downstream_arbitrationshare;
  input            custom_dma_burst_1_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_1_downstream_byteenable;
  input            custom_dma_burst_1_downstream_debugaccess;
  input            custom_dma_burst_1_downstream_latency_counter;
  input   [ 11: 0] custom_dma_burst_1_downstream_nativeaddress;
  input            custom_dma_burst_1_downstream_read;
  input            custom_dma_burst_1_downstream_write;
  input   [ 31: 0] custom_dma_burst_1_downstream_writedata;
  input   [ 11: 0] custom_dma_burst_2_downstream_address_to_slave;
  input   [  3: 0] custom_dma_burst_2_downstream_arbitrationshare;
  input            custom_dma_burst_2_downstream_burstcount;
  input   [  3: 0] custom_dma_burst_2_downstream_byteenable;
  input            custom_dma_burst_2_downstream_debugaccess;
  input            custom_dma_burst_2_downstream_latency_counter;
  input   [ 11: 0] custom_dma_burst_2_downstream_nativeaddress;
  input            custom_dma_burst_2_downstream_read;
  input            custom_dma_burst_2_downstream_write;
  input   [ 31: 0] custom_dma_burst_2_downstream_writedata;
  input            pipeline_bridge_s1_endofpacket;
  input   [ 31: 0] pipeline_bridge_s1_readdata;
  input            pipeline_bridge_s1_readdatavalid;
  input            pipeline_bridge_s1_waitrequest;
  input            reset_n;

  wire             custom_dma_burst_1_downstream_arbiterlock;
  wire             custom_dma_burst_1_downstream_arbiterlock2;
  wire             custom_dma_burst_1_downstream_continuerequest;
  wire             custom_dma_burst_1_downstream_granted_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_rdv_fifo_empty_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_rdv_fifo_output_from_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  wire             custom_dma_burst_1_downstream_requests_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_arbiterlock;
  wire             custom_dma_burst_2_downstream_arbiterlock2;
  wire             custom_dma_burst_2_downstream_continuerequest;
  wire             custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_rdv_fifo_empty_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_rdv_fifo_output_from_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  wire             custom_dma_burst_2_downstream_requests_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1;
  reg              d1_pipeline_bridge_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pipeline_bridge_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_custom_dma_burst_1_downstream_granted_slave_pipeline_bridge_s1;
  reg              last_cycle_custom_dma_burst_2_downstream_granted_slave_pipeline_bridge_s1;
  wire    [  9: 0] pipeline_bridge_s1_address;
  wire             pipeline_bridge_s1_allgrants;
  wire             pipeline_bridge_s1_allow_new_arb_cycle;
  wire             pipeline_bridge_s1_any_bursting_master_saved_grant;
  wire             pipeline_bridge_s1_any_continuerequest;
  reg     [  1: 0] pipeline_bridge_s1_arb_addend;
  wire             pipeline_bridge_s1_arb_counter_enable;
  reg     [  3: 0] pipeline_bridge_s1_arb_share_counter;
  wire    [  3: 0] pipeline_bridge_s1_arb_share_counter_next_value;
  wire    [  3: 0] pipeline_bridge_s1_arb_share_set_values;
  wire    [  1: 0] pipeline_bridge_s1_arb_winner;
  wire             pipeline_bridge_s1_arbiterlock;
  wire             pipeline_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_s1_arbitration_holdoff_internal;
  wire             pipeline_bridge_s1_beginbursttransfer_internal;
  wire             pipeline_bridge_s1_begins_xfer;
  wire             pipeline_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_s1_byteenable;
  wire             pipeline_bridge_s1_chipselect;
  wire    [  3: 0] pipeline_bridge_s1_chosen_master_double_vector;
  wire    [  1: 0] pipeline_bridge_s1_chosen_master_rot_left;
  wire             pipeline_bridge_s1_debugaccess;
  wire             pipeline_bridge_s1_end_xfer;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  wire             pipeline_bridge_s1_firsttransfer;
  wire    [  1: 0] pipeline_bridge_s1_grant_vector;
  wire             pipeline_bridge_s1_in_a_read_cycle;
  wire             pipeline_bridge_s1_in_a_write_cycle;
  wire    [  1: 0] pipeline_bridge_s1_master_qreq_vector;
  wire             pipeline_bridge_s1_move_on_to_next_transaction;
  wire    [  9: 0] pipeline_bridge_s1_nativeaddress;
  wire             pipeline_bridge_s1_non_bursting_master_requests;
  wire             pipeline_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_s1_readdatavalid_from_sa;
  reg              pipeline_bridge_s1_reg_firsttransfer;
  wire             pipeline_bridge_s1_reset_n;
  reg     [  1: 0] pipeline_bridge_s1_saved_chosen_master_vector;
  reg              pipeline_bridge_s1_slavearbiterlockenable;
  wire             pipeline_bridge_s1_slavearbiterlockenable2;
  wire             pipeline_bridge_s1_unreg_firsttransfer;
  wire             pipeline_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_s1_waits_for_read;
  wire             pipeline_bridge_s1_waits_for_write;
  wire             pipeline_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_s1_writedata;
  wire    [ 11: 0] shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_1_downstream;
  wire    [ 11: 0] shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_2_downstream;
  wire             wait_for_pipeline_bridge_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pipeline_bridge_s1_end_xfer;
    end


  assign pipeline_bridge_s1_begins_xfer = ~d1_reasons_to_wait & ((custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1 | custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1));
  //assign pipeline_bridge_s1_readdata_from_sa = pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_readdata_from_sa = pipeline_bridge_s1_readdata;

  assign custom_dma_burst_1_downstream_requests_pipeline_bridge_s1 = (1) & (custom_dma_burst_1_downstream_read | custom_dma_burst_1_downstream_write);
  //assign pipeline_bridge_s1_waitrequest_from_sa = pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_waitrequest_from_sa = pipeline_bridge_s1_waitrequest;

  //assign pipeline_bridge_s1_readdatavalid_from_sa = pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_readdatavalid_from_sa = pipeline_bridge_s1_readdatavalid;

  //pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  assign pipeline_bridge_s1_arb_share_set_values = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_arbitrationshare :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_arbitrationshare :
    (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_arbitrationshare :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_arbitrationshare :
    (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_arbitrationshare :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_arbitrationshare :
    1;

  //pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  assign pipeline_bridge_s1_non_bursting_master_requests = 0;

  //pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pipeline_bridge_s1_any_bursting_master_saved_grant = custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 |
    custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1 |
    custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 |
    custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1 |
    custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 |
    custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1;

  //pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pipeline_bridge_s1_arb_share_counter_next_value = pipeline_bridge_s1_firsttransfer ? (pipeline_bridge_s1_arb_share_set_values - 1) : |pipeline_bridge_s1_arb_share_counter ? (pipeline_bridge_s1_arb_share_counter - 1) : 0;

  //pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  assign pipeline_bridge_s1_allgrants = (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector) |
    (|pipeline_bridge_s1_grant_vector);

  //pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  assign pipeline_bridge_s1_end_xfer = ~(pipeline_bridge_s1_waits_for_read | pipeline_bridge_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pipeline_bridge_s1 = pipeline_bridge_s1_end_xfer & (~pipeline_bridge_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pipeline_bridge_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & pipeline_bridge_s1_allgrants) | (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & ~pipeline_bridge_s1_non_bursting_master_requests);

  //pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_arb_share_counter <= 0;
      else if (pipeline_bridge_s1_arb_counter_enable)
          pipeline_bridge_s1_arb_share_counter <= pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_slavearbiterlockenable <= 0;
      else if ((|pipeline_bridge_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pipeline_bridge_s1) | (end_xfer_arb_share_counter_term_pipeline_bridge_s1 & ~pipeline_bridge_s1_non_bursting_master_requests))
          pipeline_bridge_s1_slavearbiterlockenable <= |pipeline_bridge_s1_arb_share_counter_next_value;
    end


  //custom_dma_burst_1/downstream pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign custom_dma_burst_1_downstream_arbiterlock = pipeline_bridge_s1_slavearbiterlockenable & custom_dma_burst_1_downstream_continuerequest;

  //pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pipeline_bridge_s1_slavearbiterlockenable2 = |pipeline_bridge_s1_arb_share_counter_next_value;

  //custom_dma_burst_1/downstream pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign custom_dma_burst_1_downstream_arbiterlock2 = pipeline_bridge_s1_slavearbiterlockenable2 & custom_dma_burst_1_downstream_continuerequest;

  //custom_dma_burst_2/downstream pipeline_bridge/s1 arbiterlock, which is an e_assign
  assign custom_dma_burst_2_downstream_arbiterlock = pipeline_bridge_s1_slavearbiterlockenable & custom_dma_burst_2_downstream_continuerequest;

  //custom_dma_burst_2/downstream pipeline_bridge/s1 arbiterlock2, which is an e_assign
  assign custom_dma_burst_2_downstream_arbiterlock2 = pipeline_bridge_s1_slavearbiterlockenable2 & custom_dma_burst_2_downstream_continuerequest;

  //custom_dma_burst_2/downstream granted pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_2_downstream_granted_slave_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_2_downstream_granted_slave_pipeline_bridge_s1 <= custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1 ? 1 : (pipeline_bridge_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_custom_dma_burst_2_downstream_granted_slave_pipeline_bridge_s1;
    end


  //custom_dma_burst_2_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_2_downstream_continuerequest = last_cycle_custom_dma_burst_2_downstream_granted_slave_pipeline_bridge_s1 & 1;

  //pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign pipeline_bridge_s1_any_continuerequest = custom_dma_burst_2_downstream_continuerequest |
    custom_dma_burst_1_downstream_continuerequest;

  assign custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1 = custom_dma_burst_1_downstream_requests_pipeline_bridge_s1 & ~((custom_dma_burst_1_downstream_read & ((custom_dma_burst_1_downstream_latency_counter != 0) | (1 < custom_dma_burst_1_downstream_latency_counter))) | custom_dma_burst_2_downstream_arbiterlock);
  //unique name for pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  assign pipeline_bridge_s1_move_on_to_next_transaction = pipeline_bridge_s1_readdatavalid_from_sa;

  //rdv_fifo_for_custom_dma_burst_1_downstream_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_custom_dma_burst_1_downstream_to_pipeline_bridge_s1_module rdv_fifo_for_custom_dma_burst_1_downstream_to_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1),
      .data_out             (custom_dma_burst_1_downstream_rdv_fifo_output_from_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (custom_dma_burst_1_downstream_rdv_fifo_empty_pipeline_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_s1_waits_for_read)
    );

  assign custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register = ~custom_dma_burst_1_downstream_rdv_fifo_empty_pipeline_bridge_s1;
  //local readdatavalid custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1, which is an e_mux
  assign custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1 = (pipeline_bridge_s1_readdatavalid_from_sa & custom_dma_burst_1_downstream_rdv_fifo_output_from_pipeline_bridge_s1) & ~ custom_dma_burst_1_downstream_rdv_fifo_empty_pipeline_bridge_s1;

  //pipeline_bridge_s1_writedata mux, which is an e_mux
  assign pipeline_bridge_s1_writedata = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_writedata :
    custom_dma_burst_2_downstream_writedata;

  //assign pipeline_bridge_s1_endofpacket_from_sa = pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pipeline_bridge_s1_endofpacket_from_sa = pipeline_bridge_s1_endofpacket;

  assign custom_dma_burst_2_downstream_requests_pipeline_bridge_s1 = (1) & (custom_dma_burst_2_downstream_read | custom_dma_burst_2_downstream_write);
  //custom_dma_burst_1/downstream granted pipeline_bridge/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_custom_dma_burst_1_downstream_granted_slave_pipeline_bridge_s1 <= 0;
      else 
        last_cycle_custom_dma_burst_1_downstream_granted_slave_pipeline_bridge_s1 <= custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 ? 1 : (pipeline_bridge_s1_arbitration_holdoff_internal | 0) ? 0 : last_cycle_custom_dma_burst_1_downstream_granted_slave_pipeline_bridge_s1;
    end


  //custom_dma_burst_1_downstream_continuerequest continued request, which is an e_mux
  assign custom_dma_burst_1_downstream_continuerequest = last_cycle_custom_dma_burst_1_downstream_granted_slave_pipeline_bridge_s1 & 1;

  assign custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1 = custom_dma_burst_2_downstream_requests_pipeline_bridge_s1 & ~((custom_dma_burst_2_downstream_read & ((custom_dma_burst_2_downstream_latency_counter != 0) | (1 < custom_dma_burst_2_downstream_latency_counter))) | custom_dma_burst_1_downstream_arbiterlock);
  //rdv_fifo_for_custom_dma_burst_2_downstream_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_custom_dma_burst_2_downstream_to_pipeline_bridge_s1_module rdv_fifo_for_custom_dma_burst_2_downstream_to_pipeline_bridge_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1),
      .data_out             (custom_dma_burst_2_downstream_rdv_fifo_output_from_pipeline_bridge_s1),
      .empty                (),
      .fifo_contains_ones_n (custom_dma_burst_2_downstream_rdv_fifo_empty_pipeline_bridge_s1),
      .full                 (),
      .read                 (pipeline_bridge_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~pipeline_bridge_s1_waits_for_read)
    );

  assign custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register = ~custom_dma_burst_2_downstream_rdv_fifo_empty_pipeline_bridge_s1;
  //local readdatavalid custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1, which is an e_mux
  assign custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1 = (pipeline_bridge_s1_readdatavalid_from_sa & custom_dma_burst_2_downstream_rdv_fifo_output_from_pipeline_bridge_s1) & ~ custom_dma_burst_2_downstream_rdv_fifo_empty_pipeline_bridge_s1;

  //allow new arb cycle for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_allow_new_arb_cycle = ~custom_dma_burst_1_downstream_arbiterlock & ~custom_dma_burst_2_downstream_arbiterlock;

  //custom_dma_burst_2/downstream assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_master_qreq_vector[0] = custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1;

  //custom_dma_burst_2/downstream grant pipeline_bridge/s1, which is an e_assign
  assign custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 = pipeline_bridge_s1_grant_vector[0];

  //custom_dma_burst_2/downstream saved-grant pipeline_bridge/s1, which is an e_assign
  assign custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1 = pipeline_bridge_s1_arb_winner[0];

  //custom_dma_burst_1/downstream assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  assign pipeline_bridge_s1_master_qreq_vector[1] = custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1;

  //custom_dma_burst_1/downstream grant pipeline_bridge/s1, which is an e_assign
  assign custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 = pipeline_bridge_s1_grant_vector[1];

  //custom_dma_burst_1/downstream saved-grant pipeline_bridge/s1, which is an e_assign
  assign custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 = pipeline_bridge_s1_arb_winner[1];

  //pipeline_bridge/s1 chosen-master double-vector, which is an e_assign
  assign pipeline_bridge_s1_chosen_master_double_vector = {pipeline_bridge_s1_master_qreq_vector, pipeline_bridge_s1_master_qreq_vector} & ({~pipeline_bridge_s1_master_qreq_vector, ~pipeline_bridge_s1_master_qreq_vector} + pipeline_bridge_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign pipeline_bridge_s1_arb_winner = (pipeline_bridge_s1_allow_new_arb_cycle & | pipeline_bridge_s1_grant_vector) ? pipeline_bridge_s1_grant_vector : pipeline_bridge_s1_saved_chosen_master_vector;

  //saved pipeline_bridge_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_saved_chosen_master_vector <= 0;
      else if (pipeline_bridge_s1_allow_new_arb_cycle)
          pipeline_bridge_s1_saved_chosen_master_vector <= |pipeline_bridge_s1_grant_vector ? pipeline_bridge_s1_grant_vector : pipeline_bridge_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign pipeline_bridge_s1_grant_vector = {(pipeline_bridge_s1_chosen_master_double_vector[1] | pipeline_bridge_s1_chosen_master_double_vector[3]),
    (pipeline_bridge_s1_chosen_master_double_vector[0] | pipeline_bridge_s1_chosen_master_double_vector[2])};

  //pipeline_bridge/s1 chosen master rotated left, which is an e_assign
  assign pipeline_bridge_s1_chosen_master_rot_left = (pipeline_bridge_s1_arb_winner << 1) ? (pipeline_bridge_s1_arb_winner << 1) : 1;

  //pipeline_bridge/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_arb_addend <= 1;
      else if (|pipeline_bridge_s1_grant_vector)
          pipeline_bridge_s1_arb_addend <= pipeline_bridge_s1_end_xfer? pipeline_bridge_s1_chosen_master_rot_left : pipeline_bridge_s1_grant_vector;
    end


  //pipeline_bridge_s1_reset_n assignment, which is an e_assign
  assign pipeline_bridge_s1_reset_n = reset_n;

  assign pipeline_bridge_s1_chipselect = custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 | custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;
  //pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_s1_firsttransfer = pipeline_bridge_s1_begins_xfer ? pipeline_bridge_s1_unreg_firsttransfer : pipeline_bridge_s1_reg_firsttransfer;

  //pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pipeline_bridge_s1_unreg_firsttransfer = ~(pipeline_bridge_s1_slavearbiterlockenable & pipeline_bridge_s1_any_continuerequest);

  //pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_s1_reg_firsttransfer <= 1'b1;
      else if (pipeline_bridge_s1_begins_xfer)
          pipeline_bridge_s1_reg_firsttransfer <= pipeline_bridge_s1_unreg_firsttransfer;
    end


  //pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pipeline_bridge_s1_beginbursttransfer_internal = pipeline_bridge_s1_begins_xfer;

  //pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign pipeline_bridge_s1_arbitration_holdoff_internal = pipeline_bridge_s1_begins_xfer & pipeline_bridge_s1_firsttransfer;

  //pipeline_bridge_s1_read assignment, which is an e_mux
  assign pipeline_bridge_s1_read = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_1_downstream_read) | (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_2_downstream_read);

  //pipeline_bridge_s1_write assignment, which is an e_mux
  assign pipeline_bridge_s1_write = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_1_downstream_write) | (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_2_downstream_write);

  assign shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_1_downstream = custom_dma_burst_1_downstream_address_to_slave;
  //pipeline_bridge_s1_address mux, which is an e_mux
  assign pipeline_bridge_s1_address = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? (shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_1_downstream >> 2) :
    (shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_2_downstream >> 2);

  assign shifted_address_to_pipeline_bridge_s1_from_custom_dma_burst_2_downstream = custom_dma_burst_2_downstream_address_to_slave;
  //slaveid pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  assign pipeline_bridge_s1_nativeaddress = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_nativeaddress :
    custom_dma_burst_2_downstream_nativeaddress;

  //d1_pipeline_bridge_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pipeline_bridge_s1_end_xfer <= 1;
      else 
        d1_pipeline_bridge_s1_end_xfer <= pipeline_bridge_s1_end_xfer;
    end


  //pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  assign pipeline_bridge_s1_waits_for_read = pipeline_bridge_s1_in_a_read_cycle & pipeline_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  assign pipeline_bridge_s1_in_a_read_cycle = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_1_downstream_read) | (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_2_downstream_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pipeline_bridge_s1_in_a_read_cycle;

  //pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  assign pipeline_bridge_s1_waits_for_write = pipeline_bridge_s1_in_a_write_cycle & pipeline_bridge_s1_waitrequest_from_sa;

  //pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  assign pipeline_bridge_s1_in_a_write_cycle = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_1_downstream_write) | (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 & custom_dma_burst_2_downstream_write);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pipeline_bridge_s1_in_a_write_cycle;

  assign wait_for_pipeline_bridge_s1_counter = 0;
  //pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  assign pipeline_bridge_s1_byteenable = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_byteenable :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_byteenable :
    -1;

  //burstcount mux, which is an e_mux
  assign pipeline_bridge_s1_burstcount = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_burstcount :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_burstcount :
    1;

  //pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  assign pipeline_bridge_s1_arbiterlock = (custom_dma_burst_1_downstream_arbiterlock)? custom_dma_burst_1_downstream_arbiterlock :
    custom_dma_burst_2_downstream_arbiterlock;

  //pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  assign pipeline_bridge_s1_arbiterlock2 = (custom_dma_burst_1_downstream_arbiterlock2)? custom_dma_burst_1_downstream_arbiterlock2 :
    custom_dma_burst_2_downstream_arbiterlock2;

  //debugaccess mux, which is an e_mux
  assign pipeline_bridge_s1_debugaccess = (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_1_downstream_debugaccess :
    (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1)? custom_dma_burst_2_downstream_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //custom_dma_burst_1/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_1_downstream_requests_pipeline_bridge_s1 && (custom_dma_burst_1_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_1/downstream drove 0 on its 'arbitrationshare' port while accessing slave pipeline_bridge/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_1/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_1_downstream_requests_pipeline_bridge_s1 && (custom_dma_burst_1_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_1/downstream drove 0 on its 'burstcount' port while accessing slave pipeline_bridge/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_2/downstream non-zero arbitrationshare assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_2_downstream_requests_pipeline_bridge_s1 && (custom_dma_burst_2_downstream_arbitrationshare == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_2/downstream drove 0 on its 'arbitrationshare' port while accessing slave pipeline_bridge/s1", $time);
          $stop;
        end
    end


  //custom_dma_burst_2/downstream non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_2_downstream_requests_pipeline_bridge_s1 && (custom_dma_burst_2_downstream_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: custom_dma_burst_2/downstream drove 0 on its 'burstcount' port while accessing slave pipeline_bridge/s1", $time);
          $stop;
        end
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1 + custom_dma_burst_2_downstream_granted_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (custom_dma_burst_1_downstream_saved_grant_pipeline_bridge_s1 + custom_dma_burst_2_downstream_saved_grant_pipeline_bridge_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_m1_arbitrator (
                                       // inputs:
                                        clk,
                                        cpu_jtag_debug_module_readdata_from_sa,
                                        custom_dma_clock_0_in_endofpacket_from_sa,
                                        custom_dma_clock_0_in_readdata_from_sa,
                                        custom_dma_clock_0_in_waitrequest_from_sa,
                                        d1_cpu_jtag_debug_module_end_xfer,
                                        d1_custom_dma_clock_0_in_end_xfer,
                                        d1_fir_dma_control_end_xfer,
                                        d1_jtag_uart_avalon_jtag_slave_end_xfer,
                                        d1_sysid_control_slave_end_xfer,
                                        d1_timestamp_timer_s1_end_xfer,
                                        fir_dma_control_readdata_from_sa,
                                        jtag_uart_avalon_jtag_slave_readdata_from_sa,
                                        jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
                                        pipeline_bridge_m1_address,
                                        pipeline_bridge_m1_burstcount,
                                        pipeline_bridge_m1_byteenable,
                                        pipeline_bridge_m1_chipselect,
                                        pipeline_bridge_m1_granted_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_granted_custom_dma_clock_0_in,
                                        pipeline_bridge_m1_granted_fir_dma_control,
                                        pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
                                        pipeline_bridge_m1_granted_sysid_control_slave,
                                        pipeline_bridge_m1_granted_timestamp_timer_s1,
                                        pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in,
                                        pipeline_bridge_m1_qualified_request_fir_dma_control,
                                        pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
                                        pipeline_bridge_m1_qualified_request_sysid_control_slave,
                                        pipeline_bridge_m1_qualified_request_timestamp_timer_s1,
                                        pipeline_bridge_m1_read,
                                        pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in,
                                        pipeline_bridge_m1_read_data_valid_fir_dma_control,
                                        pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
                                        pipeline_bridge_m1_read_data_valid_sysid_control_slave,
                                        pipeline_bridge_m1_read_data_valid_timestamp_timer_s1,
                                        pipeline_bridge_m1_requests_cpu_jtag_debug_module,
                                        pipeline_bridge_m1_requests_custom_dma_clock_0_in,
                                        pipeline_bridge_m1_requests_fir_dma_control,
                                        pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
                                        pipeline_bridge_m1_requests_sysid_control_slave,
                                        pipeline_bridge_m1_requests_timestamp_timer_s1,
                                        pipeline_bridge_m1_write,
                                        pipeline_bridge_m1_writedata,
                                        reset_n,
                                        sysid_control_slave_readdata_from_sa,
                                        timestamp_timer_s1_readdata_from_sa,

                                       // outputs:
                                        pipeline_bridge_m1_address_to_slave,
                                        pipeline_bridge_m1_endofpacket,
                                        pipeline_bridge_m1_latency_counter,
                                        pipeline_bridge_m1_readdata,
                                        pipeline_bridge_m1_readdatavalid,
                                        pipeline_bridge_m1_waitrequest
                                     )
;

  output  [ 11: 0] pipeline_bridge_m1_address_to_slave;
  output           pipeline_bridge_m1_endofpacket;
  output           pipeline_bridge_m1_latency_counter;
  output  [ 31: 0] pipeline_bridge_m1_readdata;
  output           pipeline_bridge_m1_readdatavalid;
  output           pipeline_bridge_m1_waitrequest;
  input            clk;
  input   [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  input            custom_dma_clock_0_in_endofpacket_from_sa;
  input   [ 15: 0] custom_dma_clock_0_in_readdata_from_sa;
  input            custom_dma_clock_0_in_waitrequest_from_sa;
  input            d1_cpu_jtag_debug_module_end_xfer;
  input            d1_custom_dma_clock_0_in_end_xfer;
  input            d1_fir_dma_control_end_xfer;
  input            d1_jtag_uart_avalon_jtag_slave_end_xfer;
  input            d1_sysid_control_slave_end_xfer;
  input            d1_timestamp_timer_s1_end_xfer;
  input   [ 31: 0] fir_dma_control_readdata_from_sa;
  input   [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  input   [ 11: 0] pipeline_bridge_m1_address;
  input            pipeline_bridge_m1_burstcount;
  input   [  3: 0] pipeline_bridge_m1_byteenable;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_granted_custom_dma_clock_0_in;
  input            pipeline_bridge_m1_granted_fir_dma_control;
  input            pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  input            pipeline_bridge_m1_granted_sysid_control_slave;
  input            pipeline_bridge_m1_granted_timestamp_timer_s1;
  input            pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in;
  input            pipeline_bridge_m1_qualified_request_fir_dma_control;
  input            pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  input            pipeline_bridge_m1_qualified_request_sysid_control_slave;
  input            pipeline_bridge_m1_qualified_request_timestamp_timer_s1;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in;
  input            pipeline_bridge_m1_read_data_valid_fir_dma_control;
  input            pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  input            pipeline_bridge_m1_read_data_valid_sysid_control_slave;
  input            pipeline_bridge_m1_read_data_valid_timestamp_timer_s1;
  input            pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  input            pipeline_bridge_m1_requests_custom_dma_clock_0_in;
  input            pipeline_bridge_m1_requests_fir_dma_control;
  input            pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  input            pipeline_bridge_m1_requests_sysid_control_slave;
  input            pipeline_bridge_m1_requests_timestamp_timer_s1;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata_from_sa;
  input   [ 15: 0] timestamp_timer_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  wire             latency_load_value;
  wire             p1_pipeline_bridge_m1_latency_counter;
  reg     [ 11: 0] pipeline_bridge_m1_address_last_time;
  wire    [ 11: 0] pipeline_bridge_m1_address_to_slave;
  reg              pipeline_bridge_m1_burstcount_last_time;
  reg     [  3: 0] pipeline_bridge_m1_byteenable_last_time;
  reg              pipeline_bridge_m1_chipselect_last_time;
  wire             pipeline_bridge_m1_endofpacket;
  wire             pipeline_bridge_m1_is_granted_some_slave;
  reg              pipeline_bridge_m1_latency_counter;
  reg              pipeline_bridge_m1_read_but_no_slave_selected;
  reg              pipeline_bridge_m1_read_last_time;
  wire    [ 31: 0] pipeline_bridge_m1_readdata;
  wire             pipeline_bridge_m1_readdatavalid;
  wire             pipeline_bridge_m1_run;
  wire             pipeline_bridge_m1_waitrequest;
  reg              pipeline_bridge_m1_write_last_time;
  reg     [ 31: 0] pipeline_bridge_m1_writedata_last_time;
  wire             pre_flush_pipeline_bridge_m1_readdatavalid;
  wire             r_0;
  wire             r_1;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~pipeline_bridge_m1_requests_cpu_jtag_debug_module) & ((~pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~(pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) | (1 & ~d1_cpu_jtag_debug_module_end_xfer & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))) & ((~pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module | ~(pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect) | (1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect)))) & 1 & (pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in | ~pipeline_bridge_m1_requests_custom_dma_clock_0_in) & ((~pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in | ~pipeline_bridge_m1_chipselect | (1 & ~custom_dma_clock_0_in_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in | ~pipeline_bridge_m1_chipselect | (1 & ~custom_dma_clock_0_in_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_fir_dma_control | ~pipeline_bridge_m1_requests_fir_dma_control) & ((~pipeline_bridge_m1_qualified_request_fir_dma_control | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_fir_dma_control | ~pipeline_bridge_m1_chipselect | (1 & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave) & ((~pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pipeline_bridge_m1_chipselect | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & ((~pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave | ~pipeline_bridge_m1_chipselect | (1 & ~jtag_uart_avalon_jtag_slave_waitrequest_from_sa & pipeline_bridge_m1_chipselect))) & 1 & (pipeline_bridge_m1_qualified_request_sysid_control_slave | ~pipeline_bridge_m1_requests_sysid_control_slave) & ((~pipeline_bridge_m1_qualified_request_sysid_control_slave | ~(pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) | (1 & ~d1_sysid_control_slave_end_xfer & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))) & ((~pipeline_bridge_m1_qualified_request_sysid_control_slave | ~(pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect) | (1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect))));

  //cascaded wait assignment, which is an e_assign
  assign pipeline_bridge_m1_run = r_0 & r_1;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (pipeline_bridge_m1_qualified_request_timestamp_timer_s1 | ~pipeline_bridge_m1_requests_timestamp_timer_s1) & ((~pipeline_bridge_m1_qualified_request_timestamp_timer_s1 | ~(pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) | (1 & ~d1_timestamp_timer_s1_end_xfer & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))) & ((~pipeline_bridge_m1_qualified_request_timestamp_timer_s1 | ~(pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect) | (1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect))));

  //optimize select-logic by passing only those address bits which matter.
  assign pipeline_bridge_m1_address_to_slave = pipeline_bridge_m1_address[11 : 0];

  //pipeline_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_but_no_slave_selected <= 0;
      else 
        pipeline_bridge_m1_read_but_no_slave_selected <= (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & pipeline_bridge_m1_run & ~pipeline_bridge_m1_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign pipeline_bridge_m1_is_granted_some_slave = pipeline_bridge_m1_granted_cpu_jtag_debug_module |
    pipeline_bridge_m1_granted_custom_dma_clock_0_in |
    pipeline_bridge_m1_granted_fir_dma_control |
    pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave |
    pipeline_bridge_m1_granted_sysid_control_slave |
    pipeline_bridge_m1_granted_timestamp_timer_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_pipeline_bridge_m1_readdatavalid = pipeline_bridge_m1_read_data_valid_fir_dma_control;

  //latent slave read data valid which is not flushed, which is an e_mux
  assign pipeline_bridge_m1_readdatavalid = pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_sysid_control_slave |
    pipeline_bridge_m1_read_but_no_slave_selected |
    pre_flush_pipeline_bridge_m1_readdatavalid |
    pipeline_bridge_m1_read_data_valid_timestamp_timer_s1;

  //pipeline_bridge/m1 readdata mux, which is an e_mux
  assign pipeline_bridge_m1_readdata = ({32 {~((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | cpu_jtag_debug_module_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | custom_dma_clock_0_in_readdata_from_sa) &
    ({32 {~pipeline_bridge_m1_read_data_valid_fir_dma_control}} | fir_dma_control_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | jtag_uart_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_sysid_control_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | sysid_control_slave_readdata_from_sa) &
    ({32 {~((pipeline_bridge_m1_qualified_request_timestamp_timer_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))}} | timestamp_timer_s1_readdata_from_sa);

  //actual waitrequest port, which is an e_assign
  assign pipeline_bridge_m1_waitrequest = ~pipeline_bridge_m1_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_latency_counter <= 0;
      else 
        pipeline_bridge_m1_latency_counter <= p1_pipeline_bridge_m1_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_pipeline_bridge_m1_latency_counter = ((pipeline_bridge_m1_run & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect)))? latency_load_value :
    (pipeline_bridge_m1_latency_counter)? pipeline_bridge_m1_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {1 {pipeline_bridge_m1_requests_fir_dma_control}} & 1;

  //mux pipeline_bridge_m1_endofpacket, which is an e_mux
  assign pipeline_bridge_m1_endofpacket = custom_dma_clock_0_in_endofpacket_from_sa;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pipeline_bridge_m1_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_address_last_time <= 0;
      else 
        pipeline_bridge_m1_address_last_time <= pipeline_bridge_m1_address;
    end


  //pipeline_bridge/m1 waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= pipeline_bridge_m1_waitrequest & pipeline_bridge_m1_chipselect;
    end


  //pipeline_bridge_m1_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_address != pipeline_bridge_m1_address_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_chipselect check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_chipselect_last_time <= 0;
      else 
        pipeline_bridge_m1_chipselect_last_time <= pipeline_bridge_m1_chipselect;
    end


  //pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_chipselect != pipeline_bridge_m1_chipselect_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_chipselect did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_burstcount check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_burstcount_last_time <= 0;
      else 
        pipeline_bridge_m1_burstcount_last_time <= pipeline_bridge_m1_burstcount;
    end


  //pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_burstcount != pipeline_bridge_m1_burstcount_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_burstcount did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_byteenable_last_time <= 0;
      else 
        pipeline_bridge_m1_byteenable_last_time <= pipeline_bridge_m1_byteenable;
    end


  //pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_byteenable != pipeline_bridge_m1_byteenable_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_read_last_time <= 0;
      else 
        pipeline_bridge_m1_read_last_time <= pipeline_bridge_m1_read;
    end


  //pipeline_bridge_m1_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_read != pipeline_bridge_m1_read_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_write_last_time <= 0;
      else 
        pipeline_bridge_m1_write_last_time <= pipeline_bridge_m1_write;
    end


  //pipeline_bridge_m1_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_write != pipeline_bridge_m1_write_last_time))
        begin
          $write("%0d ns: pipeline_bridge_m1_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //pipeline_bridge_m1_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pipeline_bridge_m1_writedata_last_time <= 0;
      else 
        pipeline_bridge_m1_writedata_last_time <= pipeline_bridge_m1_writedata;
    end


  //pipeline_bridge_m1_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (pipeline_bridge_m1_writedata != pipeline_bridge_m1_writedata_last_time) & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect))
        begin
          $write("%0d ns: pipeline_bridge_m1_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pll_s1_arbitrator (
                           // inputs:
                            clk,
                            custom_dma_clock_0_out_address_to_slave,
                            custom_dma_clock_0_out_nativeaddress,
                            custom_dma_clock_0_out_read,
                            custom_dma_clock_0_out_write,
                            custom_dma_clock_0_out_writedata,
                            pll_s1_readdata,
                            pll_s1_resetrequest,
                            reset_n,

                           // outputs:
                            custom_dma_clock_0_out_granted_pll_s1,
                            custom_dma_clock_0_out_qualified_request_pll_s1,
                            custom_dma_clock_0_out_read_data_valid_pll_s1,
                            custom_dma_clock_0_out_requests_pll_s1,
                            d1_pll_s1_end_xfer,
                            pll_s1_address,
                            pll_s1_chipselect,
                            pll_s1_read,
                            pll_s1_readdata_from_sa,
                            pll_s1_reset_n,
                            pll_s1_resetrequest_from_sa,
                            pll_s1_write,
                            pll_s1_writedata
                         )
;

  output           custom_dma_clock_0_out_granted_pll_s1;
  output           custom_dma_clock_0_out_qualified_request_pll_s1;
  output           custom_dma_clock_0_out_read_data_valid_pll_s1;
  output           custom_dma_clock_0_out_requests_pll_s1;
  output           d1_pll_s1_end_xfer;
  output  [  2: 0] pll_s1_address;
  output           pll_s1_chipselect;
  output           pll_s1_read;
  output  [ 15: 0] pll_s1_readdata_from_sa;
  output           pll_s1_reset_n;
  output           pll_s1_resetrequest_from_sa;
  output           pll_s1_write;
  output  [ 15: 0] pll_s1_writedata;
  input            clk;
  input   [  3: 0] custom_dma_clock_0_out_address_to_slave;
  input   [  2: 0] custom_dma_clock_0_out_nativeaddress;
  input            custom_dma_clock_0_out_read;
  input            custom_dma_clock_0_out_write;
  input   [ 15: 0] custom_dma_clock_0_out_writedata;
  input   [ 15: 0] pll_s1_readdata;
  input            pll_s1_resetrequest;
  input            reset_n;

  wire             custom_dma_clock_0_out_arbiterlock;
  wire             custom_dma_clock_0_out_arbiterlock2;
  wire             custom_dma_clock_0_out_continuerequest;
  wire             custom_dma_clock_0_out_granted_pll_s1;
  wire             custom_dma_clock_0_out_qualified_request_pll_s1;
  wire             custom_dma_clock_0_out_read_data_valid_pll_s1;
  wire             custom_dma_clock_0_out_requests_pll_s1;
  wire             custom_dma_clock_0_out_saved_grant_pll_s1;
  reg              d1_pll_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_pll_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_allgrants;
  wire             pll_s1_allow_new_arb_cycle;
  wire             pll_s1_any_bursting_master_saved_grant;
  wire             pll_s1_any_continuerequest;
  wire             pll_s1_arb_counter_enable;
  reg              pll_s1_arb_share_counter;
  wire             pll_s1_arb_share_counter_next_value;
  wire             pll_s1_arb_share_set_values;
  wire             pll_s1_beginbursttransfer_internal;
  wire             pll_s1_begins_xfer;
  wire             pll_s1_chipselect;
  wire             pll_s1_end_xfer;
  wire             pll_s1_firsttransfer;
  wire             pll_s1_grant_vector;
  wire             pll_s1_in_a_read_cycle;
  wire             pll_s1_in_a_write_cycle;
  wire             pll_s1_master_qreq_vector;
  wire             pll_s1_non_bursting_master_requests;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  reg              pll_s1_reg_firsttransfer;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest_from_sa;
  reg              pll_s1_slavearbiterlockenable;
  wire             pll_s1_slavearbiterlockenable2;
  wire             pll_s1_unreg_firsttransfer;
  wire             pll_s1_waits_for_read;
  wire             pll_s1_waits_for_write;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             wait_for_pll_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~pll_s1_end_xfer;
    end


  assign pll_s1_begins_xfer = ~d1_reasons_to_wait & ((custom_dma_clock_0_out_qualified_request_pll_s1));
  //assign pll_s1_readdata_from_sa = pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_readdata_from_sa = pll_s1_readdata;

  assign custom_dma_clock_0_out_requests_pll_s1 = (1) & (custom_dma_clock_0_out_read | custom_dma_clock_0_out_write);
  //pll_s1_arb_share_counter set values, which is an e_mux
  assign pll_s1_arb_share_set_values = 1;

  //pll_s1_non_bursting_master_requests mux, which is an e_mux
  assign pll_s1_non_bursting_master_requests = custom_dma_clock_0_out_requests_pll_s1;

  //pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign pll_s1_any_bursting_master_saved_grant = 0;

  //pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign pll_s1_arb_share_counter_next_value = pll_s1_firsttransfer ? (pll_s1_arb_share_set_values - 1) : |pll_s1_arb_share_counter ? (pll_s1_arb_share_counter - 1) : 0;

  //pll_s1_allgrants all slave grants, which is an e_mux
  assign pll_s1_allgrants = |pll_s1_grant_vector;

  //pll_s1_end_xfer assignment, which is an e_assign
  assign pll_s1_end_xfer = ~(pll_s1_waits_for_read | pll_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_pll_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_pll_s1 = pll_s1_end_xfer & (~pll_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign pll_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_pll_s1 & pll_s1_allgrants) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests);

  //pll_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_arb_share_counter <= 0;
      else if (pll_s1_arb_counter_enable)
          pll_s1_arb_share_counter <= pll_s1_arb_share_counter_next_value;
    end


  //pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_slavearbiterlockenable <= 0;
      else if ((|pll_s1_master_qreq_vector & end_xfer_arb_share_counter_term_pll_s1) | (end_xfer_arb_share_counter_term_pll_s1 & ~pll_s1_non_bursting_master_requests))
          pll_s1_slavearbiterlockenable <= |pll_s1_arb_share_counter_next_value;
    end


  //custom_dma_clock_0/out pll/s1 arbiterlock, which is an e_assign
  assign custom_dma_clock_0_out_arbiterlock = pll_s1_slavearbiterlockenable & custom_dma_clock_0_out_continuerequest;

  //pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign pll_s1_slavearbiterlockenable2 = |pll_s1_arb_share_counter_next_value;

  //custom_dma_clock_0/out pll/s1 arbiterlock2, which is an e_assign
  assign custom_dma_clock_0_out_arbiterlock2 = pll_s1_slavearbiterlockenable2 & custom_dma_clock_0_out_continuerequest;

  //pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign pll_s1_any_continuerequest = 1;

  //custom_dma_clock_0_out_continuerequest continued request, which is an e_assign
  assign custom_dma_clock_0_out_continuerequest = 1;

  assign custom_dma_clock_0_out_qualified_request_pll_s1 = custom_dma_clock_0_out_requests_pll_s1;
  //pll_s1_writedata mux, which is an e_mux
  assign pll_s1_writedata = custom_dma_clock_0_out_writedata;

  //master is always granted when requested
  assign custom_dma_clock_0_out_granted_pll_s1 = custom_dma_clock_0_out_qualified_request_pll_s1;

  //custom_dma_clock_0/out saved-grant pll/s1, which is an e_assign
  assign custom_dma_clock_0_out_saved_grant_pll_s1 = custom_dma_clock_0_out_requests_pll_s1;

  //allow new arb cycle for pll/s1, which is an e_assign
  assign pll_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign pll_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign pll_s1_master_qreq_vector = 1;

  //pll_s1_reset_n assignment, which is an e_assign
  assign pll_s1_reset_n = reset_n;

  //assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest;

  assign pll_s1_chipselect = custom_dma_clock_0_out_granted_pll_s1;
  //pll_s1_firsttransfer first transaction, which is an e_assign
  assign pll_s1_firsttransfer = pll_s1_begins_xfer ? pll_s1_unreg_firsttransfer : pll_s1_reg_firsttransfer;

  //pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign pll_s1_unreg_firsttransfer = ~(pll_s1_slavearbiterlockenable & pll_s1_any_continuerequest);

  //pll_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pll_s1_reg_firsttransfer <= 1'b1;
      else if (pll_s1_begins_xfer)
          pll_s1_reg_firsttransfer <= pll_s1_unreg_firsttransfer;
    end


  //pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign pll_s1_beginbursttransfer_internal = pll_s1_begins_xfer;

  //pll_s1_read assignment, which is an e_mux
  assign pll_s1_read = custom_dma_clock_0_out_granted_pll_s1 & custom_dma_clock_0_out_read;

  //pll_s1_write assignment, which is an e_mux
  assign pll_s1_write = custom_dma_clock_0_out_granted_pll_s1 & custom_dma_clock_0_out_write;

  //pll_s1_address mux, which is an e_mux
  assign pll_s1_address = custom_dma_clock_0_out_nativeaddress;

  //d1_pll_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_pll_s1_end_xfer <= 1;
      else 
        d1_pll_s1_end_xfer <= pll_s1_end_xfer;
    end


  //pll_s1_waits_for_read in a cycle, which is an e_mux
  assign pll_s1_waits_for_read = pll_s1_in_a_read_cycle & pll_s1_begins_xfer;

  //pll_s1_in_a_read_cycle assignment, which is an e_assign
  assign pll_s1_in_a_read_cycle = custom_dma_clock_0_out_granted_pll_s1 & custom_dma_clock_0_out_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = pll_s1_in_a_read_cycle;

  //pll_s1_waits_for_write in a cycle, which is an e_mux
  assign pll_s1_waits_for_write = pll_s1_in_a_write_cycle & 0;

  //pll_s1_in_a_write_cycle assignment, which is an e_assign
  assign pll_s1_in_a_write_cycle = custom_dma_clock_0_out_granted_pll_s1 & custom_dma_clock_0_out_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = pll_s1_in_a_write_cycle;

  assign wait_for_pll_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //pll/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid_control_slave_arbitrator (
                                        // inputs:
                                         clk,
                                         pipeline_bridge_m1_address_to_slave,
                                         pipeline_bridge_m1_burstcount,
                                         pipeline_bridge_m1_chipselect,
                                         pipeline_bridge_m1_latency_counter,
                                         pipeline_bridge_m1_read,
                                         pipeline_bridge_m1_write,
                                         reset_n,
                                         sysid_control_slave_readdata,

                                        // outputs:
                                         d1_sysid_control_slave_end_xfer,
                                         pipeline_bridge_m1_granted_sysid_control_slave,
                                         pipeline_bridge_m1_qualified_request_sysid_control_slave,
                                         pipeline_bridge_m1_read_data_valid_sysid_control_slave,
                                         pipeline_bridge_m1_requests_sysid_control_slave,
                                         sysid_control_slave_address,
                                         sysid_control_slave_readdata_from_sa
                                      )
;

  output           d1_sysid_control_slave_end_xfer;
  output           pipeline_bridge_m1_granted_sysid_control_slave;
  output           pipeline_bridge_m1_qualified_request_sysid_control_slave;
  output           pipeline_bridge_m1_read_data_valid_sysid_control_slave;
  output           pipeline_bridge_m1_requests_sysid_control_slave;
  output           sysid_control_slave_address;
  output  [ 31: 0] sysid_control_slave_readdata_from_sa;
  input            clk;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input            reset_n;
  input   [ 31: 0] sysid_control_slave_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_sysid_control_slave_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sysid_control_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_sysid_control_slave;
  wire             pipeline_bridge_m1_qualified_request_sysid_control_slave;
  wire             pipeline_bridge_m1_read_data_valid_sysid_control_slave;
  wire             pipeline_bridge_m1_requests_sysid_control_slave;
  wire             pipeline_bridge_m1_saved_grant_sysid_control_slave;
  wire    [ 11: 0] shifted_address_to_sysid_control_slave_from_pipeline_bridge_m1;
  wire             sysid_control_slave_address;
  wire             sysid_control_slave_allgrants;
  wire             sysid_control_slave_allow_new_arb_cycle;
  wire             sysid_control_slave_any_bursting_master_saved_grant;
  wire             sysid_control_slave_any_continuerequest;
  wire             sysid_control_slave_arb_counter_enable;
  reg              sysid_control_slave_arb_share_counter;
  wire             sysid_control_slave_arb_share_counter_next_value;
  wire             sysid_control_slave_arb_share_set_values;
  wire             sysid_control_slave_beginbursttransfer_internal;
  wire             sysid_control_slave_begins_xfer;
  wire             sysid_control_slave_end_xfer;
  wire             sysid_control_slave_firsttransfer;
  wire             sysid_control_slave_grant_vector;
  wire             sysid_control_slave_in_a_read_cycle;
  wire             sysid_control_slave_in_a_write_cycle;
  wire             sysid_control_slave_master_qreq_vector;
  wire             sysid_control_slave_non_bursting_master_requests;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  reg              sysid_control_slave_reg_firsttransfer;
  reg              sysid_control_slave_slavearbiterlockenable;
  wire             sysid_control_slave_slavearbiterlockenable2;
  wire             sysid_control_slave_unreg_firsttransfer;
  wire             sysid_control_slave_waits_for_read;
  wire             sysid_control_slave_waits_for_write;
  wire             wait_for_sysid_control_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sysid_control_slave_end_xfer;
    end


  assign sysid_control_slave_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_sysid_control_slave));
  //assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sysid_control_slave_readdata_from_sa = sysid_control_slave_readdata;

  assign pipeline_bridge_m1_requests_sysid_control_slave = (({pipeline_bridge_m1_address_to_slave[11 : 3] , 3'b0} == 12'h860) & pipeline_bridge_m1_chipselect) & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);
  //sysid_control_slave_arb_share_counter set values, which is an e_mux
  assign sysid_control_slave_arb_share_set_values = 1;

  //sysid_control_slave_non_bursting_master_requests mux, which is an e_mux
  assign sysid_control_slave_non_bursting_master_requests = pipeline_bridge_m1_requests_sysid_control_slave;

  //sysid_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign sysid_control_slave_any_bursting_master_saved_grant = 0;

  //sysid_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign sysid_control_slave_arb_share_counter_next_value = sysid_control_slave_firsttransfer ? (sysid_control_slave_arb_share_set_values - 1) : |sysid_control_slave_arb_share_counter ? (sysid_control_slave_arb_share_counter - 1) : 0;

  //sysid_control_slave_allgrants all slave grants, which is an e_mux
  assign sysid_control_slave_allgrants = |sysid_control_slave_grant_vector;

  //sysid_control_slave_end_xfer assignment, which is an e_assign
  assign sysid_control_slave_end_xfer = ~(sysid_control_slave_waits_for_read | sysid_control_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_sysid_control_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sysid_control_slave = sysid_control_slave_end_xfer & (~sysid_control_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sysid_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign sysid_control_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_sysid_control_slave & sysid_control_slave_allgrants) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests);

  //sysid_control_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_arb_share_counter <= 0;
      else if (sysid_control_slave_arb_counter_enable)
          sysid_control_slave_arb_share_counter <= sysid_control_slave_arb_share_counter_next_value;
    end


  //sysid_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_slavearbiterlockenable <= 0;
      else if ((|sysid_control_slave_master_qreq_vector & end_xfer_arb_share_counter_term_sysid_control_slave) | (end_xfer_arb_share_counter_term_sysid_control_slave & ~sysid_control_slave_non_bursting_master_requests))
          sysid_control_slave_slavearbiterlockenable <= |sysid_control_slave_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 sysid/control_slave arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = sysid_control_slave_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //sysid_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sysid_control_slave_slavearbiterlockenable2 = |sysid_control_slave_arb_share_counter_next_value;

  //pipeline_bridge/m1 sysid/control_slave arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = sysid_control_slave_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //sysid_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign sysid_control_slave_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_sysid_control_slave = pipeline_bridge_m1_requests_sysid_control_slave & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_sysid_control_slave, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_sysid_control_slave = pipeline_bridge_m1_granted_sysid_control_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~sysid_control_slave_waits_for_read;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_sysid_control_slave = pipeline_bridge_m1_qualified_request_sysid_control_slave;

  //pipeline_bridge/m1 saved-grant sysid/control_slave, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_sysid_control_slave = pipeline_bridge_m1_requests_sysid_control_slave;

  //allow new arb cycle for sysid/control_slave, which is an e_assign
  assign sysid_control_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign sysid_control_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign sysid_control_slave_master_qreq_vector = 1;

  //sysid_control_slave_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_firsttransfer = sysid_control_slave_begins_xfer ? sysid_control_slave_unreg_firsttransfer : sysid_control_slave_reg_firsttransfer;

  //sysid_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign sysid_control_slave_unreg_firsttransfer = ~(sysid_control_slave_slavearbiterlockenable & sysid_control_slave_any_continuerequest);

  //sysid_control_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sysid_control_slave_reg_firsttransfer <= 1'b1;
      else if (sysid_control_slave_begins_xfer)
          sysid_control_slave_reg_firsttransfer <= sysid_control_slave_unreg_firsttransfer;
    end


  //sysid_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sysid_control_slave_beginbursttransfer_internal = sysid_control_slave_begins_xfer;

  assign shifted_address_to_sysid_control_slave_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //sysid_control_slave_address mux, which is an e_mux
  assign sysid_control_slave_address = shifted_address_to_sysid_control_slave_from_pipeline_bridge_m1 >> 2;

  //d1_sysid_control_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sysid_control_slave_end_xfer <= 1;
      else 
        d1_sysid_control_slave_end_xfer <= sysid_control_slave_end_xfer;
    end


  //sysid_control_slave_waits_for_read in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_read = sysid_control_slave_in_a_read_cycle & sysid_control_slave_begins_xfer;

  //sysid_control_slave_in_a_read_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_read_cycle = pipeline_bridge_m1_granted_sysid_control_slave & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sysid_control_slave_in_a_read_cycle;

  //sysid_control_slave_waits_for_write in a cycle, which is an e_mux
  assign sysid_control_slave_waits_for_write = sysid_control_slave_in_a_write_cycle & 0;

  //sysid_control_slave_in_a_write_cycle assignment, which is an e_assign
  assign sysid_control_slave_in_a_write_cycle = pipeline_bridge_m1_granted_sysid_control_slave & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sysid_control_slave_in_a_write_cycle;

  assign wait_for_sysid_control_slave_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sysid/control_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_sysid_control_slave && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sysid/control_slave", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module timestamp_timer_s1_arbitrator (
                                       // inputs:
                                        clk,
                                        pipeline_bridge_m1_address_to_slave,
                                        pipeline_bridge_m1_burstcount,
                                        pipeline_bridge_m1_chipselect,
                                        pipeline_bridge_m1_latency_counter,
                                        pipeline_bridge_m1_read,
                                        pipeline_bridge_m1_write,
                                        pipeline_bridge_m1_writedata,
                                        reset_n,
                                        timestamp_timer_s1_irq,
                                        timestamp_timer_s1_readdata,

                                       // outputs:
                                        d1_timestamp_timer_s1_end_xfer,
                                        pipeline_bridge_m1_granted_timestamp_timer_s1,
                                        pipeline_bridge_m1_qualified_request_timestamp_timer_s1,
                                        pipeline_bridge_m1_read_data_valid_timestamp_timer_s1,
                                        pipeline_bridge_m1_requests_timestamp_timer_s1,
                                        timestamp_timer_s1_address,
                                        timestamp_timer_s1_chipselect,
                                        timestamp_timer_s1_irq_from_sa,
                                        timestamp_timer_s1_readdata_from_sa,
                                        timestamp_timer_s1_reset_n,
                                        timestamp_timer_s1_write_n,
                                        timestamp_timer_s1_writedata
                                     )
;

  output           d1_timestamp_timer_s1_end_xfer;
  output           pipeline_bridge_m1_granted_timestamp_timer_s1;
  output           pipeline_bridge_m1_qualified_request_timestamp_timer_s1;
  output           pipeline_bridge_m1_read_data_valid_timestamp_timer_s1;
  output           pipeline_bridge_m1_requests_timestamp_timer_s1;
  output  [  2: 0] timestamp_timer_s1_address;
  output           timestamp_timer_s1_chipselect;
  output           timestamp_timer_s1_irq_from_sa;
  output  [ 15: 0] timestamp_timer_s1_readdata_from_sa;
  output           timestamp_timer_s1_reset_n;
  output           timestamp_timer_s1_write_n;
  output  [ 15: 0] timestamp_timer_s1_writedata;
  input            clk;
  input   [ 11: 0] pipeline_bridge_m1_address_to_slave;
  input            pipeline_bridge_m1_burstcount;
  input            pipeline_bridge_m1_chipselect;
  input            pipeline_bridge_m1_latency_counter;
  input            pipeline_bridge_m1_read;
  input            pipeline_bridge_m1_write;
  input   [ 31: 0] pipeline_bridge_m1_writedata;
  input            reset_n;
  input            timestamp_timer_s1_irq;
  input   [ 15: 0] timestamp_timer_s1_readdata;

  reg              d1_reasons_to_wait;
  reg              d1_timestamp_timer_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_timestamp_timer_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             pipeline_bridge_m1_arbiterlock;
  wire             pipeline_bridge_m1_arbiterlock2;
  wire             pipeline_bridge_m1_continuerequest;
  wire             pipeline_bridge_m1_granted_timestamp_timer_s1;
  wire             pipeline_bridge_m1_qualified_request_timestamp_timer_s1;
  wire             pipeline_bridge_m1_read_data_valid_timestamp_timer_s1;
  wire             pipeline_bridge_m1_requests_timestamp_timer_s1;
  wire             pipeline_bridge_m1_saved_grant_timestamp_timer_s1;
  wire    [ 11: 0] shifted_address_to_timestamp_timer_s1_from_pipeline_bridge_m1;
  wire    [  2: 0] timestamp_timer_s1_address;
  wire             timestamp_timer_s1_allgrants;
  wire             timestamp_timer_s1_allow_new_arb_cycle;
  wire             timestamp_timer_s1_any_bursting_master_saved_grant;
  wire             timestamp_timer_s1_any_continuerequest;
  wire             timestamp_timer_s1_arb_counter_enable;
  reg              timestamp_timer_s1_arb_share_counter;
  wire             timestamp_timer_s1_arb_share_counter_next_value;
  wire             timestamp_timer_s1_arb_share_set_values;
  wire             timestamp_timer_s1_beginbursttransfer_internal;
  wire             timestamp_timer_s1_begins_xfer;
  wire             timestamp_timer_s1_chipselect;
  wire             timestamp_timer_s1_end_xfer;
  wire             timestamp_timer_s1_firsttransfer;
  wire             timestamp_timer_s1_grant_vector;
  wire             timestamp_timer_s1_in_a_read_cycle;
  wire             timestamp_timer_s1_in_a_write_cycle;
  wire             timestamp_timer_s1_irq_from_sa;
  wire             timestamp_timer_s1_master_qreq_vector;
  wire             timestamp_timer_s1_non_bursting_master_requests;
  wire    [ 15: 0] timestamp_timer_s1_readdata_from_sa;
  reg              timestamp_timer_s1_reg_firsttransfer;
  wire             timestamp_timer_s1_reset_n;
  reg              timestamp_timer_s1_slavearbiterlockenable;
  wire             timestamp_timer_s1_slavearbiterlockenable2;
  wire             timestamp_timer_s1_unreg_firsttransfer;
  wire             timestamp_timer_s1_waits_for_read;
  wire             timestamp_timer_s1_waits_for_write;
  wire             timestamp_timer_s1_write_n;
  wire    [ 15: 0] timestamp_timer_s1_writedata;
  wire             wait_for_timestamp_timer_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~timestamp_timer_s1_end_xfer;
    end


  assign timestamp_timer_s1_begins_xfer = ~d1_reasons_to_wait & ((pipeline_bridge_m1_qualified_request_timestamp_timer_s1));
  //assign timestamp_timer_s1_readdata_from_sa = timestamp_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign timestamp_timer_s1_readdata_from_sa = timestamp_timer_s1_readdata;

  assign pipeline_bridge_m1_requests_timestamp_timer_s1 = ({pipeline_bridge_m1_address_to_slave[11 : 5] , 5'b0} == 12'h800) & pipeline_bridge_m1_chipselect;
  //timestamp_timer_s1_arb_share_counter set values, which is an e_mux
  assign timestamp_timer_s1_arb_share_set_values = 1;

  //timestamp_timer_s1_non_bursting_master_requests mux, which is an e_mux
  assign timestamp_timer_s1_non_bursting_master_requests = pipeline_bridge_m1_requests_timestamp_timer_s1;

  //timestamp_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign timestamp_timer_s1_any_bursting_master_saved_grant = 0;

  //timestamp_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign timestamp_timer_s1_arb_share_counter_next_value = timestamp_timer_s1_firsttransfer ? (timestamp_timer_s1_arb_share_set_values - 1) : |timestamp_timer_s1_arb_share_counter ? (timestamp_timer_s1_arb_share_counter - 1) : 0;

  //timestamp_timer_s1_allgrants all slave grants, which is an e_mux
  assign timestamp_timer_s1_allgrants = |timestamp_timer_s1_grant_vector;

  //timestamp_timer_s1_end_xfer assignment, which is an e_assign
  assign timestamp_timer_s1_end_xfer = ~(timestamp_timer_s1_waits_for_read | timestamp_timer_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_timestamp_timer_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_timestamp_timer_s1 = timestamp_timer_s1_end_xfer & (~timestamp_timer_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //timestamp_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign timestamp_timer_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_timestamp_timer_s1 & timestamp_timer_s1_allgrants) | (end_xfer_arb_share_counter_term_timestamp_timer_s1 & ~timestamp_timer_s1_non_bursting_master_requests);

  //timestamp_timer_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timestamp_timer_s1_arb_share_counter <= 0;
      else if (timestamp_timer_s1_arb_counter_enable)
          timestamp_timer_s1_arb_share_counter <= timestamp_timer_s1_arb_share_counter_next_value;
    end


  //timestamp_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timestamp_timer_s1_slavearbiterlockenable <= 0;
      else if ((|timestamp_timer_s1_master_qreq_vector & end_xfer_arb_share_counter_term_timestamp_timer_s1) | (end_xfer_arb_share_counter_term_timestamp_timer_s1 & ~timestamp_timer_s1_non_bursting_master_requests))
          timestamp_timer_s1_slavearbiterlockenable <= |timestamp_timer_s1_arb_share_counter_next_value;
    end


  //pipeline_bridge/m1 timestamp_timer/s1 arbiterlock, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock = timestamp_timer_s1_slavearbiterlockenable & pipeline_bridge_m1_continuerequest;

  //timestamp_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign timestamp_timer_s1_slavearbiterlockenable2 = |timestamp_timer_s1_arb_share_counter_next_value;

  //pipeline_bridge/m1 timestamp_timer/s1 arbiterlock2, which is an e_assign
  assign pipeline_bridge_m1_arbiterlock2 = timestamp_timer_s1_slavearbiterlockenable2 & pipeline_bridge_m1_continuerequest;

  //timestamp_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign timestamp_timer_s1_any_continuerequest = 1;

  //pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  assign pipeline_bridge_m1_continuerequest = 1;

  assign pipeline_bridge_m1_qualified_request_timestamp_timer_s1 = pipeline_bridge_m1_requests_timestamp_timer_s1 & ~(((pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ((pipeline_bridge_m1_latency_counter != 0))));
  //local readdatavalid pipeline_bridge_m1_read_data_valid_timestamp_timer_s1, which is an e_mux
  assign pipeline_bridge_m1_read_data_valid_timestamp_timer_s1 = pipeline_bridge_m1_granted_timestamp_timer_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect) & ~timestamp_timer_s1_waits_for_read;

  //timestamp_timer_s1_writedata mux, which is an e_mux
  assign timestamp_timer_s1_writedata = pipeline_bridge_m1_writedata;

  //master is always granted when requested
  assign pipeline_bridge_m1_granted_timestamp_timer_s1 = pipeline_bridge_m1_qualified_request_timestamp_timer_s1;

  //pipeline_bridge/m1 saved-grant timestamp_timer/s1, which is an e_assign
  assign pipeline_bridge_m1_saved_grant_timestamp_timer_s1 = pipeline_bridge_m1_requests_timestamp_timer_s1;

  //allow new arb cycle for timestamp_timer/s1, which is an e_assign
  assign timestamp_timer_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign timestamp_timer_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign timestamp_timer_s1_master_qreq_vector = 1;

  //timestamp_timer_s1_reset_n assignment, which is an e_assign
  assign timestamp_timer_s1_reset_n = reset_n;

  assign timestamp_timer_s1_chipselect = pipeline_bridge_m1_granted_timestamp_timer_s1;
  //timestamp_timer_s1_firsttransfer first transaction, which is an e_assign
  assign timestamp_timer_s1_firsttransfer = timestamp_timer_s1_begins_xfer ? timestamp_timer_s1_unreg_firsttransfer : timestamp_timer_s1_reg_firsttransfer;

  //timestamp_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign timestamp_timer_s1_unreg_firsttransfer = ~(timestamp_timer_s1_slavearbiterlockenable & timestamp_timer_s1_any_continuerequest);

  //timestamp_timer_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timestamp_timer_s1_reg_firsttransfer <= 1'b1;
      else if (timestamp_timer_s1_begins_xfer)
          timestamp_timer_s1_reg_firsttransfer <= timestamp_timer_s1_unreg_firsttransfer;
    end


  //timestamp_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign timestamp_timer_s1_beginbursttransfer_internal = timestamp_timer_s1_begins_xfer;

  //~timestamp_timer_s1_write_n assignment, which is an e_mux
  assign timestamp_timer_s1_write_n = ~(pipeline_bridge_m1_granted_timestamp_timer_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect));

  assign shifted_address_to_timestamp_timer_s1_from_pipeline_bridge_m1 = pipeline_bridge_m1_address_to_slave;
  //timestamp_timer_s1_address mux, which is an e_mux
  assign timestamp_timer_s1_address = shifted_address_to_timestamp_timer_s1_from_pipeline_bridge_m1 >> 2;

  //d1_timestamp_timer_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_timestamp_timer_s1_end_xfer <= 1;
      else 
        d1_timestamp_timer_s1_end_xfer <= timestamp_timer_s1_end_xfer;
    end


  //timestamp_timer_s1_waits_for_read in a cycle, which is an e_mux
  assign timestamp_timer_s1_waits_for_read = timestamp_timer_s1_in_a_read_cycle & timestamp_timer_s1_begins_xfer;

  //timestamp_timer_s1_in_a_read_cycle assignment, which is an e_assign
  assign timestamp_timer_s1_in_a_read_cycle = pipeline_bridge_m1_granted_timestamp_timer_s1 & (pipeline_bridge_m1_read & pipeline_bridge_m1_chipselect);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = timestamp_timer_s1_in_a_read_cycle;

  //timestamp_timer_s1_waits_for_write in a cycle, which is an e_mux
  assign timestamp_timer_s1_waits_for_write = timestamp_timer_s1_in_a_write_cycle & 0;

  //timestamp_timer_s1_in_a_write_cycle assignment, which is an e_assign
  assign timestamp_timer_s1_in_a_write_cycle = pipeline_bridge_m1_granted_timestamp_timer_s1 & (pipeline_bridge_m1_write & pipeline_bridge_m1_chipselect);

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = timestamp_timer_s1_in_a_write_cycle;

  assign wait_for_timestamp_timer_s1_counter = 0;
  //assign timestamp_timer_s1_irq_from_sa = timestamp_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign timestamp_timer_s1_irq_from_sa = timestamp_timer_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //timestamp_timer/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
  always @(posedge clk)
    begin
      if (pipeline_bridge_m1_requests_timestamp_timer_s1 && (pipeline_bridge_m1_burstcount == 0) && enable_nonzero_assertions)
        begin
          $write("%0d ns: pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave timestamp_timer/s1", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_reset_system_clk_domain_synch_module (
                                                         // inputs:
                                                          clk,
                                                          data_in,
                                                          reset_n,

                                                         // outputs:
                                                          data_out
                                                       )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_reset_external_clk_domain_synch_module (
                                                           // inputs:
                                                            clk,
                                                            data_in,
                                                            reset_n,

                                                           // outputs:
                                                            data_out
                                                         )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma (
                    // 1) global signals:
                     external_clk,
                     reset_n,
                     sdram_write_clk,
                     ssram_clk,
                     system_clk,

                    // the_ddr_sdram
                     clk_to_sdram_from_the_ddr_sdram,
                     clk_to_sdram_n_from_the_ddr_sdram,
                     ddr_a_from_the_ddr_sdram,
                     ddr_ba_from_the_ddr_sdram,
                     ddr_cas_n_from_the_ddr_sdram,
                     ddr_cke_from_the_ddr_sdram,
                     ddr_cs_n_from_the_ddr_sdram,
                     ddr_dm_from_the_ddr_sdram,
                     ddr_dq_to_and_from_the_ddr_sdram,
                     ddr_dqs_to_and_from_the_ddr_sdram,
                     ddr_ras_n_from_the_ddr_sdram,
                     ddr_we_n_from_the_ddr_sdram,
                     dqs_delay_ctrl_to_the_ddr_sdram,
                     dqsupdate_to_the_ddr_sdram,
                     stratix_dll_control_from_the_ddr_sdram,
                     write_clk_to_the_ddr_sdram,

                    // the_ext_ssram_bus_avalon_slave
                     adsc_n_to_the_ext_ssram,
                     bw_n_to_the_ext_ssram,
                     bwe_n_to_the_ext_ssram,
                     chipenable1_n_to_the_ext_ssram,
                     ext_ssram_bus_address,
                     ext_ssram_bus_data,
                     outputenable_n_to_the_ext_ssram
                  )
;

  output           adsc_n_to_the_ext_ssram;
  output  [  3: 0] bw_n_to_the_ext_ssram;
  output           bwe_n_to_the_ext_ssram;
  output           chipenable1_n_to_the_ext_ssram;
  output           clk_to_sdram_from_the_ddr_sdram;
  output           clk_to_sdram_n_from_the_ddr_sdram;
  output  [ 12: 0] ddr_a_from_the_ddr_sdram;
  output  [  1: 0] ddr_ba_from_the_ddr_sdram;
  output           ddr_cas_n_from_the_ddr_sdram;
  output           ddr_cke_from_the_ddr_sdram;
  output           ddr_cs_n_from_the_ddr_sdram;
  output  [  1: 0] ddr_dm_from_the_ddr_sdram;
  inout   [ 15: 0] ddr_dq_to_and_from_the_ddr_sdram;
  inout   [  1: 0] ddr_dqs_to_and_from_the_ddr_sdram;
  output           ddr_ras_n_from_the_ddr_sdram;
  output           ddr_we_n_from_the_ddr_sdram;
  output  [ 20: 0] ext_ssram_bus_address;
  inout   [ 31: 0] ext_ssram_bus_data;
  output           outputenable_n_to_the_ext_ssram;
  output           sdram_write_clk;
  output           ssram_clk;
  output           stratix_dll_control_from_the_ddr_sdram;
  output           system_clk;
  input   [  5: 0] dqs_delay_ctrl_to_the_ddr_sdram;
  input            dqsupdate_to_the_ddr_sdram;
  input            external_clk;
  input            reset_n;
  input            write_clk_to_the_ddr_sdram;

  wire             adsc_n_to_the_ext_ssram;
  wire    [  3: 0] bw_n_to_the_ext_ssram;
  wire             bwe_n_to_the_ext_ssram;
  wire             chipenable1_n_to_the_ext_ssram;
  wire             clk_to_sdram_from_the_ddr_sdram;
  wire             clk_to_sdram_n_from_the_ddr_sdram;
  wire    [ 26: 0] cpu_data_master_address;
  wire    [ 26: 0] cpu_data_master_address_to_slave;
  wire    [  3: 0] cpu_data_master_burstcount;
  wire    [  3: 0] cpu_data_master_byteenable;
  wire             cpu_data_master_debugaccess;
  wire             cpu_data_master_granted_custom_dma_burst_0_upstream;
  wire             cpu_data_master_granted_custom_dma_burst_2_upstream;
  wire             cpu_data_master_granted_custom_dma_burst_4_upstream;
  wire    [ 31: 0] cpu_data_master_irq;
  wire             cpu_data_master_latency_counter;
  wire             cpu_data_master_qualified_request_custom_dma_burst_0_upstream;
  wire             cpu_data_master_qualified_request_custom_dma_burst_2_upstream;
  wire             cpu_data_master_qualified_request_custom_dma_burst_4_upstream;
  wire             cpu_data_master_read;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_0_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_2_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_4_upstream;
  wire             cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register;
  wire    [ 31: 0] cpu_data_master_readdata;
  wire             cpu_data_master_readdatavalid;
  wire             cpu_data_master_requests_custom_dma_burst_0_upstream;
  wire             cpu_data_master_requests_custom_dma_burst_2_upstream;
  wire             cpu_data_master_requests_custom_dma_burst_4_upstream;
  wire             cpu_data_master_waitrequest;
  wire             cpu_data_master_write;
  wire    [ 31: 0] cpu_data_master_writedata;
  wire    [ 26: 0] cpu_instruction_master_address;
  wire    [ 26: 0] cpu_instruction_master_address_to_slave;
  wire    [  3: 0] cpu_instruction_master_burstcount;
  wire             cpu_instruction_master_granted_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_granted_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_latency_counter;
  wire             cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_read;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register;
  wire    [ 31: 0] cpu_instruction_master_readdata;
  wire             cpu_instruction_master_readdatavalid;
  wire             cpu_instruction_master_requests_custom_dma_burst_1_upstream;
  wire             cpu_instruction_master_requests_custom_dma_burst_3_upstream;
  wire             cpu_instruction_master_waitrequest;
  wire    [  8: 0] cpu_jtag_debug_module_address;
  wire             cpu_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_jtag_debug_module_byteenable;
  wire             cpu_jtag_debug_module_chipselect;
  wire             cpu_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_jtag_debug_module_readdata_from_sa;
  wire             cpu_jtag_debug_module_reset_n;
  wire             cpu_jtag_debug_module_resetrequest;
  wire             cpu_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_jtag_debug_module_write;
  wire    [ 31: 0] cpu_jtag_debug_module_writedata;
  wire    [ 20: 0] custom_dma_burst_0_downstream_address;
  wire    [ 20: 0] custom_dma_burst_0_downstream_address_to_slave;
  wire    [  3: 0] custom_dma_burst_0_downstream_arbitrationshare;
  wire             custom_dma_burst_0_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_0_downstream_byteenable;
  wire             custom_dma_burst_0_downstream_debugaccess;
  wire             custom_dma_burst_0_downstream_granted_ext_ssram_s1;
  wire    [  2: 0] custom_dma_burst_0_downstream_latency_counter;
  wire    [ 20: 0] custom_dma_burst_0_downstream_nativeaddress;
  wire             custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1;
  wire             custom_dma_burst_0_downstream_read;
  wire             custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1;
  wire    [ 31: 0] custom_dma_burst_0_downstream_readdata;
  wire             custom_dma_burst_0_downstream_readdatavalid;
  wire             custom_dma_burst_0_downstream_requests_ext_ssram_s1;
  wire             custom_dma_burst_0_downstream_reset_n;
  wire             custom_dma_burst_0_downstream_waitrequest;
  wire             custom_dma_burst_0_downstream_write;
  wire    [ 31: 0] custom_dma_burst_0_downstream_writedata;
  wire    [ 20: 0] custom_dma_burst_0_upstream_address;
  wire    [  3: 0] custom_dma_burst_0_upstream_burstcount;
  wire    [ 22: 0] custom_dma_burst_0_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_0_upstream_byteenable;
  wire             custom_dma_burst_0_upstream_debugaccess;
  wire             custom_dma_burst_0_upstream_read;
  wire    [ 31: 0] custom_dma_burst_0_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_0_upstream_readdata_from_sa;
  wire             custom_dma_burst_0_upstream_readdatavalid;
  wire             custom_dma_burst_0_upstream_waitrequest;
  wire             custom_dma_burst_0_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_0_upstream_write;
  wire    [ 31: 0] custom_dma_burst_0_upstream_writedata;
  wire    [ 11: 0] custom_dma_burst_1_downstream_address;
  wire    [ 11: 0] custom_dma_burst_1_downstream_address_to_slave;
  wire    [  3: 0] custom_dma_burst_1_downstream_arbitrationshare;
  wire             custom_dma_burst_1_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_1_downstream_byteenable;
  wire             custom_dma_burst_1_downstream_debugaccess;
  wire             custom_dma_burst_1_downstream_granted_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_latency_counter;
  wire    [ 11: 0] custom_dma_burst_1_downstream_nativeaddress;
  wire             custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_read;
  wire             custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  wire    [ 31: 0] custom_dma_burst_1_downstream_readdata;
  wire             custom_dma_burst_1_downstream_readdatavalid;
  wire             custom_dma_burst_1_downstream_requests_pipeline_bridge_s1;
  wire             custom_dma_burst_1_downstream_reset_n;
  wire             custom_dma_burst_1_downstream_waitrequest;
  wire             custom_dma_burst_1_downstream_write;
  wire    [ 31: 0] custom_dma_burst_1_downstream_writedata;
  wire    [ 11: 0] custom_dma_burst_1_upstream_address;
  wire    [ 13: 0] custom_dma_burst_1_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_1_upstream_byteenable;
  wire             custom_dma_burst_1_upstream_debugaccess;
  wire             custom_dma_burst_1_upstream_read;
  wire    [ 31: 0] custom_dma_burst_1_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_1_upstream_readdata_from_sa;
  wire             custom_dma_burst_1_upstream_readdatavalid;
  wire             custom_dma_burst_1_upstream_waitrequest;
  wire             custom_dma_burst_1_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_1_upstream_write;
  wire    [ 31: 0] custom_dma_burst_1_upstream_writedata;
  wire    [ 11: 0] custom_dma_burst_2_downstream_address;
  wire    [ 11: 0] custom_dma_burst_2_downstream_address_to_slave;
  wire    [  3: 0] custom_dma_burst_2_downstream_arbitrationshare;
  wire             custom_dma_burst_2_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_2_downstream_byteenable;
  wire             custom_dma_burst_2_downstream_debugaccess;
  wire             custom_dma_burst_2_downstream_granted_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_latency_counter;
  wire    [ 11: 0] custom_dma_burst_2_downstream_nativeaddress;
  wire             custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_read;
  wire             custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register;
  wire    [ 31: 0] custom_dma_burst_2_downstream_readdata;
  wire             custom_dma_burst_2_downstream_readdatavalid;
  wire             custom_dma_burst_2_downstream_requests_pipeline_bridge_s1;
  wire             custom_dma_burst_2_downstream_reset_n;
  wire             custom_dma_burst_2_downstream_waitrequest;
  wire             custom_dma_burst_2_downstream_write;
  wire    [ 31: 0] custom_dma_burst_2_downstream_writedata;
  wire    [ 11: 0] custom_dma_burst_2_upstream_address;
  wire    [  3: 0] custom_dma_burst_2_upstream_burstcount;
  wire    [ 13: 0] custom_dma_burst_2_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_2_upstream_byteenable;
  wire             custom_dma_burst_2_upstream_debugaccess;
  wire             custom_dma_burst_2_upstream_read;
  wire    [ 31: 0] custom_dma_burst_2_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_2_upstream_readdata_from_sa;
  wire             custom_dma_burst_2_upstream_readdatavalid;
  wire             custom_dma_burst_2_upstream_waitrequest;
  wire             custom_dma_burst_2_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_2_upstream_write;
  wire    [ 31: 0] custom_dma_burst_2_upstream_writedata;
  wire    [ 24: 0] custom_dma_burst_3_downstream_address;
  wire    [ 24: 0] custom_dma_burst_3_downstream_address_to_slave;
  wire    [  3: 0] custom_dma_burst_3_downstream_arbitrationshare;
  wire    [  2: 0] custom_dma_burst_3_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_3_downstream_byteenable;
  wire             custom_dma_burst_3_downstream_debugaccess;
  wire             custom_dma_burst_3_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_latency_counter;
  wire    [ 24: 0] custom_dma_burst_3_downstream_nativeaddress;
  wire             custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_read;
  wire             custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire    [ 31: 0] custom_dma_burst_3_downstream_readdata;
  wire             custom_dma_burst_3_downstream_readdatavalid;
  wire             custom_dma_burst_3_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_3_downstream_reset_n;
  wire             custom_dma_burst_3_downstream_waitrequest;
  wire             custom_dma_burst_3_downstream_write;
  wire    [ 31: 0] custom_dma_burst_3_downstream_writedata;
  wire    [ 24: 0] custom_dma_burst_3_upstream_address;
  wire    [ 26: 0] custom_dma_burst_3_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_3_upstream_byteenable;
  wire             custom_dma_burst_3_upstream_debugaccess;
  wire             custom_dma_burst_3_upstream_read;
  wire    [ 31: 0] custom_dma_burst_3_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_3_upstream_readdata_from_sa;
  wire             custom_dma_burst_3_upstream_readdatavalid;
  wire             custom_dma_burst_3_upstream_waitrequest;
  wire             custom_dma_burst_3_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_3_upstream_write;
  wire    [ 31: 0] custom_dma_burst_3_upstream_writedata;
  wire    [ 24: 0] custom_dma_burst_4_downstream_address;
  wire    [ 24: 0] custom_dma_burst_4_downstream_address_to_slave;
  wire    [  3: 0] custom_dma_burst_4_downstream_arbitrationshare;
  wire    [  2: 0] custom_dma_burst_4_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_4_downstream_byteenable;
  wire             custom_dma_burst_4_downstream_debugaccess;
  wire             custom_dma_burst_4_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_latency_counter;
  wire    [ 24: 0] custom_dma_burst_4_downstream_nativeaddress;
  wire             custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_read;
  wire             custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire    [ 31: 0] custom_dma_burst_4_downstream_readdata;
  wire             custom_dma_burst_4_downstream_readdatavalid;
  wire             custom_dma_burst_4_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_4_downstream_reset_n;
  wire             custom_dma_burst_4_downstream_waitrequest;
  wire             custom_dma_burst_4_downstream_write;
  wire    [ 31: 0] custom_dma_burst_4_downstream_writedata;
  wire    [ 24: 0] custom_dma_burst_4_upstream_address;
  wire    [  3: 0] custom_dma_burst_4_upstream_burstcount;
  wire    [ 26: 0] custom_dma_burst_4_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_4_upstream_byteenable;
  wire             custom_dma_burst_4_upstream_debugaccess;
  wire             custom_dma_burst_4_upstream_read;
  wire    [ 31: 0] custom_dma_burst_4_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_4_upstream_readdata_from_sa;
  wire             custom_dma_burst_4_upstream_readdatavalid;
  wire             custom_dma_burst_4_upstream_waitrequest;
  wire             custom_dma_burst_4_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_4_upstream_write;
  wire    [ 31: 0] custom_dma_burst_4_upstream_writedata;
  wire    [ 24: 0] custom_dma_burst_5_downstream_address;
  wire    [ 24: 0] custom_dma_burst_5_downstream_address_to_slave;
  wire    [  2: 0] custom_dma_burst_5_downstream_arbitrationshare;
  wire    [  2: 0] custom_dma_burst_5_downstream_burstcount;
  wire    [  3: 0] custom_dma_burst_5_downstream_byteenable;
  wire             custom_dma_burst_5_downstream_debugaccess;
  wire             custom_dma_burst_5_downstream_granted_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_latency_counter;
  wire    [ 24: 0] custom_dma_burst_5_downstream_nativeaddress;
  wire             custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_read;
  wire             custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register;
  wire    [ 31: 0] custom_dma_burst_5_downstream_readdata;
  wire             custom_dma_burst_5_downstream_readdatavalid;
  wire             custom_dma_burst_5_downstream_requests_ddr_sdram_s1;
  wire             custom_dma_burst_5_downstream_reset_n;
  wire             custom_dma_burst_5_downstream_waitrequest;
  wire             custom_dma_burst_5_downstream_write;
  wire    [ 31: 0] custom_dma_burst_5_downstream_writedata;
  wire    [ 24: 0] custom_dma_burst_5_upstream_address;
  wire    [  2: 0] custom_dma_burst_5_upstream_burstcount;
  wire    [ 26: 0] custom_dma_burst_5_upstream_byteaddress;
  wire    [  3: 0] custom_dma_burst_5_upstream_byteenable;
  wire             custom_dma_burst_5_upstream_debugaccess;
  wire             custom_dma_burst_5_upstream_read;
  wire    [ 31: 0] custom_dma_burst_5_upstream_readdata;
  wire    [ 31: 0] custom_dma_burst_5_upstream_readdata_from_sa;
  wire             custom_dma_burst_5_upstream_readdatavalid;
  wire             custom_dma_burst_5_upstream_readdatavalid_from_sa;
  wire             custom_dma_burst_5_upstream_waitrequest;
  wire             custom_dma_burst_5_upstream_waitrequest_from_sa;
  wire             custom_dma_burst_5_upstream_write;
  wire    [ 31: 0] custom_dma_burst_5_upstream_writedata;
  wire    [  3: 0] custom_dma_clock_0_in_address;
  wire    [  1: 0] custom_dma_clock_0_in_byteenable;
  wire             custom_dma_clock_0_in_endofpacket;
  wire             custom_dma_clock_0_in_endofpacket_from_sa;
  wire    [  2: 0] custom_dma_clock_0_in_nativeaddress;
  wire             custom_dma_clock_0_in_read;
  wire    [ 15: 0] custom_dma_clock_0_in_readdata;
  wire    [ 15: 0] custom_dma_clock_0_in_readdata_from_sa;
  wire             custom_dma_clock_0_in_reset_n;
  wire             custom_dma_clock_0_in_waitrequest;
  wire             custom_dma_clock_0_in_waitrequest_from_sa;
  wire             custom_dma_clock_0_in_write;
  wire    [ 15: 0] custom_dma_clock_0_in_writedata;
  wire    [  3: 0] custom_dma_clock_0_out_address;
  wire    [  3: 0] custom_dma_clock_0_out_address_to_slave;
  wire    [  1: 0] custom_dma_clock_0_out_byteenable;
  wire             custom_dma_clock_0_out_endofpacket;
  wire             custom_dma_clock_0_out_granted_pll_s1;
  wire    [  2: 0] custom_dma_clock_0_out_nativeaddress;
  wire             custom_dma_clock_0_out_qualified_request_pll_s1;
  wire             custom_dma_clock_0_out_read;
  wire             custom_dma_clock_0_out_read_data_valid_pll_s1;
  wire    [ 15: 0] custom_dma_clock_0_out_readdata;
  wire             custom_dma_clock_0_out_requests_pll_s1;
  wire             custom_dma_clock_0_out_reset_n;
  wire             custom_dma_clock_0_out_waitrequest;
  wire             custom_dma_clock_0_out_write;
  wire    [ 15: 0] custom_dma_clock_0_out_writedata;
  wire             d1_cpu_jtag_debug_module_end_xfer;
  wire             d1_custom_dma_burst_0_upstream_end_xfer;
  wire             d1_custom_dma_burst_1_upstream_end_xfer;
  wire             d1_custom_dma_burst_2_upstream_end_xfer;
  wire             d1_custom_dma_burst_3_upstream_end_xfer;
  wire             d1_custom_dma_burst_4_upstream_end_xfer;
  wire             d1_custom_dma_burst_5_upstream_end_xfer;
  wire             d1_custom_dma_clock_0_in_end_xfer;
  wire             d1_ddr_sdram_s1_end_xfer;
  wire             d1_ext_ssram_bus_avalon_slave_end_xfer;
  wire             d1_fir_dma_control_end_xfer;
  wire             d1_jtag_uart_avalon_jtag_slave_end_xfer;
  wire             d1_pipeline_bridge_s1_end_xfer;
  wire             d1_pll_s1_end_xfer;
  wire             d1_sysid_control_slave_end_xfer;
  wire             d1_timestamp_timer_s1_end_xfer;
  wire    [ 12: 0] ddr_a_from_the_ddr_sdram;
  wire    [  1: 0] ddr_ba_from_the_ddr_sdram;
  wire             ddr_cas_n_from_the_ddr_sdram;
  wire             ddr_cke_from_the_ddr_sdram;
  wire             ddr_cs_n_from_the_ddr_sdram;
  wire    [  1: 0] ddr_dm_from_the_ddr_sdram;
  wire    [ 15: 0] ddr_dq_to_and_from_the_ddr_sdram;
  wire    [  1: 0] ddr_dqs_to_and_from_the_ddr_sdram;
  wire             ddr_ras_n_from_the_ddr_sdram;
  wire    [ 22: 0] ddr_sdram_s1_address;
  wire             ddr_sdram_s1_beginbursttransfer;
  wire    [  2: 0] ddr_sdram_s1_burstcount;
  wire    [  3: 0] ddr_sdram_s1_byteenable;
  wire             ddr_sdram_s1_read;
  wire    [ 31: 0] ddr_sdram_s1_readdata;
  wire    [ 31: 0] ddr_sdram_s1_readdata_from_sa;
  wire             ddr_sdram_s1_readdatavalid;
  wire             ddr_sdram_s1_reset_n;
  wire             ddr_sdram_s1_waitrequest_n;
  wire             ddr_sdram_s1_waitrequest_n_from_sa;
  wire             ddr_sdram_s1_write;
  wire    [ 31: 0] ddr_sdram_s1_writedata;
  wire             ddr_we_n_from_the_ddr_sdram;
  wire    [ 20: 0] ext_ssram_bus_address;
  wire    [ 31: 0] ext_ssram_bus_data;
  wire             external_clk_reset_n;
  wire    [  2: 0] fir_dma_control_address;
  wire    [  3: 0] fir_dma_control_byteenable;
  wire             fir_dma_control_irq;
  wire             fir_dma_control_irq_from_sa;
  wire             fir_dma_control_read;
  wire    [ 31: 0] fir_dma_control_readdata;
  wire    [ 31: 0] fir_dma_control_readdata_from_sa;
  wire             fir_dma_control_reset;
  wire             fir_dma_control_write;
  wire    [ 31: 0] fir_dma_control_writedata;
  wire    [ 31: 0] fir_dma_read_master_address;
  wire    [ 31: 0] fir_dma_read_master_address_to_slave;
  wire    [  3: 0] fir_dma_read_master_byteenable;
  wire             fir_dma_read_master_granted_ext_ssram_s1;
  wire    [  2: 0] fir_dma_read_master_latency_counter;
  wire             fir_dma_read_master_qualified_request_ext_ssram_s1;
  wire             fir_dma_read_master_read;
  wire             fir_dma_read_master_read_data_valid_ext_ssram_s1;
  wire    [ 31: 0] fir_dma_read_master_readdata;
  wire             fir_dma_read_master_readdatavalid;
  wire             fir_dma_read_master_requests_ext_ssram_s1;
  wire             fir_dma_read_master_waitrequest;
  wire    [ 31: 0] fir_dma_write_master_address;
  wire    [ 31: 0] fir_dma_write_master_address_to_slave;
  wire    [  2: 0] fir_dma_write_master_burstcount;
  wire    [  3: 0] fir_dma_write_master_byteenable;
  wire             fir_dma_write_master_granted_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_requests_custom_dma_burst_5_upstream;
  wire             fir_dma_write_master_waitrequest;
  wire             fir_dma_write_master_write;
  wire    [ 31: 0] fir_dma_write_master_writedata;
  wire    [ 31: 0] incoming_ext_ssram_bus_data;
  wire             jtag_uart_avalon_jtag_slave_address;
  wire             jtag_uart_avalon_jtag_slave_chipselect;
  wire             jtag_uart_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_irq;
  wire             jtag_uart_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_avalon_jtag_slave_reset_n;
  wire             jtag_uart_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_avalon_jtag_slave_writedata;
  wire             out_clk_pll_c0;
  wire             out_clk_pll_c1;
  wire             out_clk_pll_c2;
  wire             outputenable_n_to_the_ext_ssram;
  wire    [ 11: 0] pipeline_bridge_m1_address;
  wire    [ 11: 0] pipeline_bridge_m1_address_to_slave;
  wire             pipeline_bridge_m1_burstcount;
  wire    [  3: 0] pipeline_bridge_m1_byteenable;
  wire             pipeline_bridge_m1_chipselect;
  wire             pipeline_bridge_m1_debugaccess;
  wire             pipeline_bridge_m1_endofpacket;
  wire             pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_granted_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_granted_fir_dma_control;
  wire             pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_granted_sysid_control_slave;
  wire             pipeline_bridge_m1_granted_timestamp_timer_s1;
  wire             pipeline_bridge_m1_latency_counter;
  wire             pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_qualified_request_fir_dma_control;
  wire             pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_qualified_request_sysid_control_slave;
  wire             pipeline_bridge_m1_qualified_request_timestamp_timer_s1;
  wire             pipeline_bridge_m1_read;
  wire             pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_read_data_valid_fir_dma_control;
  wire             pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_read_data_valid_sysid_control_slave;
  wire             pipeline_bridge_m1_read_data_valid_timestamp_timer_s1;
  wire    [ 31: 0] pipeline_bridge_m1_readdata;
  wire             pipeline_bridge_m1_readdatavalid;
  wire             pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  wire             pipeline_bridge_m1_requests_custom_dma_clock_0_in;
  wire             pipeline_bridge_m1_requests_fir_dma_control;
  wire             pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  wire             pipeline_bridge_m1_requests_sysid_control_slave;
  wire             pipeline_bridge_m1_requests_timestamp_timer_s1;
  wire             pipeline_bridge_m1_waitrequest;
  wire             pipeline_bridge_m1_write;
  wire    [ 31: 0] pipeline_bridge_m1_writedata;
  wire    [  9: 0] pipeline_bridge_s1_address;
  wire             pipeline_bridge_s1_arbiterlock;
  wire             pipeline_bridge_s1_arbiterlock2;
  wire             pipeline_bridge_s1_burstcount;
  wire    [  3: 0] pipeline_bridge_s1_byteenable;
  wire             pipeline_bridge_s1_chipselect;
  wire             pipeline_bridge_s1_debugaccess;
  wire             pipeline_bridge_s1_endofpacket;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  wire    [  9: 0] pipeline_bridge_s1_nativeaddress;
  wire             pipeline_bridge_s1_read;
  wire    [ 31: 0] pipeline_bridge_s1_readdata;
  wire    [ 31: 0] pipeline_bridge_s1_readdata_from_sa;
  wire             pipeline_bridge_s1_readdatavalid;
  wire             pipeline_bridge_s1_reset_n;
  wire             pipeline_bridge_s1_waitrequest;
  wire             pipeline_bridge_s1_waitrequest_from_sa;
  wire             pipeline_bridge_s1_write;
  wire    [ 31: 0] pipeline_bridge_s1_writedata;
  wire    [  2: 0] pll_s1_address;
  wire             pll_s1_chipselect;
  wire             pll_s1_read;
  wire    [ 15: 0] pll_s1_readdata;
  wire    [ 15: 0] pll_s1_readdata_from_sa;
  wire             pll_s1_reset_n;
  wire             pll_s1_resetrequest;
  wire             pll_s1_resetrequest_from_sa;
  wire             pll_s1_write;
  wire    [ 15: 0] pll_s1_writedata;
  wire             reset_n_sources;
  wire             sdram_write_clk;
  wire             ssram_clk;
  wire             stratix_dll_control_from_the_ddr_sdram;
  wire             sysid_control_slave_address;
  wire    [ 31: 0] sysid_control_slave_readdata;
  wire    [ 31: 0] sysid_control_slave_readdata_from_sa;
  wire             system_clk;
  wire             system_clk_reset_n;
  wire    [  2: 0] timestamp_timer_s1_address;
  wire             timestamp_timer_s1_chipselect;
  wire             timestamp_timer_s1_irq;
  wire             timestamp_timer_s1_irq_from_sa;
  wire    [ 15: 0] timestamp_timer_s1_readdata;
  wire    [ 15: 0] timestamp_timer_s1_readdata_from_sa;
  wire             timestamp_timer_s1_reset_n;
  wire             timestamp_timer_s1_write_n;
  wire    [ 15: 0] timestamp_timer_s1_writedata;
  cpu_jtag_debug_module_arbitrator the_cpu_jtag_debug_module
    (
      .clk                                                        (system_clk),
      .cpu_jtag_debug_module_address                              (cpu_jtag_debug_module_address),
      .cpu_jtag_debug_module_begintransfer                        (cpu_jtag_debug_module_begintransfer),
      .cpu_jtag_debug_module_byteenable                           (cpu_jtag_debug_module_byteenable),
      .cpu_jtag_debug_module_chipselect                           (cpu_jtag_debug_module_chipselect),
      .cpu_jtag_debug_module_debugaccess                          (cpu_jtag_debug_module_debugaccess),
      .cpu_jtag_debug_module_readdata                             (cpu_jtag_debug_module_readdata),
      .cpu_jtag_debug_module_readdata_from_sa                     (cpu_jtag_debug_module_readdata_from_sa),
      .cpu_jtag_debug_module_reset_n                              (cpu_jtag_debug_module_reset_n),
      .cpu_jtag_debug_module_resetrequest                         (cpu_jtag_debug_module_resetrequest),
      .cpu_jtag_debug_module_resetrequest_from_sa                 (cpu_jtag_debug_module_resetrequest_from_sa),
      .cpu_jtag_debug_module_write                                (cpu_jtag_debug_module_write),
      .cpu_jtag_debug_module_writedata                            (cpu_jtag_debug_module_writedata),
      .d1_cpu_jtag_debug_module_end_xfer                          (d1_cpu_jtag_debug_module_end_xfer),
      .pipeline_bridge_m1_address_to_slave                        (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                              (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                              (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                              (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_debugaccess                             (pipeline_bridge_m1_debugaccess),
      .pipeline_bridge_m1_granted_cpu_jtag_debug_module           (pipeline_bridge_m1_granted_cpu_jtag_debug_module),
      .pipeline_bridge_m1_latency_counter                         (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module),
      .pipeline_bridge_m1_read                                    (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module   (pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module),
      .pipeline_bridge_m1_requests_cpu_jtag_debug_module          (pipeline_bridge_m1_requests_cpu_jtag_debug_module),
      .pipeline_bridge_m1_write                                   (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                               (pipeline_bridge_m1_writedata),
      .reset_n                                                    (system_clk_reset_n)
    );

  cpu_data_master_arbitrator the_cpu_data_master
    (
      .clk                                                                        (system_clk),
      .cpu_data_master_address                                                    (cpu_data_master_address),
      .cpu_data_master_address_to_slave                                           (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                 (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                 (cpu_data_master_byteenable),
      .cpu_data_master_granted_custom_dma_burst_0_upstream                        (cpu_data_master_granted_custom_dma_burst_0_upstream),
      .cpu_data_master_granted_custom_dma_burst_2_upstream                        (cpu_data_master_granted_custom_dma_burst_2_upstream),
      .cpu_data_master_granted_custom_dma_burst_4_upstream                        (cpu_data_master_granted_custom_dma_burst_4_upstream),
      .cpu_data_master_irq                                                        (cpu_data_master_irq),
      .cpu_data_master_latency_counter                                            (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_custom_dma_burst_0_upstream              (cpu_data_master_qualified_request_custom_dma_burst_0_upstream),
      .cpu_data_master_qualified_request_custom_dma_burst_2_upstream              (cpu_data_master_qualified_request_custom_dma_burst_2_upstream),
      .cpu_data_master_qualified_request_custom_dma_burst_4_upstream              (cpu_data_master_qualified_request_custom_dma_burst_4_upstream),
      .cpu_data_master_read                                                       (cpu_data_master_read),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register),
      .cpu_data_master_readdata                                                   (cpu_data_master_readdata),
      .cpu_data_master_readdatavalid                                              (cpu_data_master_readdatavalid),
      .cpu_data_master_requests_custom_dma_burst_0_upstream                       (cpu_data_master_requests_custom_dma_burst_0_upstream),
      .cpu_data_master_requests_custom_dma_burst_2_upstream                       (cpu_data_master_requests_custom_dma_burst_2_upstream),
      .cpu_data_master_requests_custom_dma_burst_4_upstream                       (cpu_data_master_requests_custom_dma_burst_4_upstream),
      .cpu_data_master_waitrequest                                                (cpu_data_master_waitrequest),
      .cpu_data_master_write                                                      (cpu_data_master_write),
      .cpu_data_master_writedata                                                  (cpu_data_master_writedata),
      .custom_dma_burst_0_upstream_readdata_from_sa                               (custom_dma_burst_0_upstream_readdata_from_sa),
      .custom_dma_burst_0_upstream_waitrequest_from_sa                            (custom_dma_burst_0_upstream_waitrequest_from_sa),
      .custom_dma_burst_2_upstream_readdata_from_sa                               (custom_dma_burst_2_upstream_readdata_from_sa),
      .custom_dma_burst_2_upstream_waitrequest_from_sa                            (custom_dma_burst_2_upstream_waitrequest_from_sa),
      .custom_dma_burst_4_upstream_readdata_from_sa                               (custom_dma_burst_4_upstream_readdata_from_sa),
      .custom_dma_burst_4_upstream_waitrequest_from_sa                            (custom_dma_burst_4_upstream_waitrequest_from_sa),
      .d1_custom_dma_burst_0_upstream_end_xfer                                    (d1_custom_dma_burst_0_upstream_end_xfer),
      .d1_custom_dma_burst_2_upstream_end_xfer                                    (d1_custom_dma_burst_2_upstream_end_xfer),
      .d1_custom_dma_burst_4_upstream_end_xfer                                    (d1_custom_dma_burst_4_upstream_end_xfer),
      .fir_dma_control_irq_from_sa                                                (fir_dma_control_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                                    (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .reset_n                                                                    (system_clk_reset_n),
      .timestamp_timer_s1_irq_from_sa                                             (timestamp_timer_s1_irq_from_sa)
    );

  cpu_instruction_master_arbitrator the_cpu_instruction_master
    (
      .clk                                                                               (system_clk),
      .cpu_instruction_master_address                                                    (cpu_instruction_master_address),
      .cpu_instruction_master_address_to_slave                                           (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                 (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_custom_dma_burst_1_upstream                        (cpu_instruction_master_granted_custom_dma_burst_1_upstream),
      .cpu_instruction_master_granted_custom_dma_burst_3_upstream                        (cpu_instruction_master_granted_custom_dma_burst_3_upstream),
      .cpu_instruction_master_latency_counter                                            (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream              (cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream),
      .cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream              (cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream),
      .cpu_instruction_master_read                                                       (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream                (cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream                (cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register),
      .cpu_instruction_master_readdata                                                   (cpu_instruction_master_readdata),
      .cpu_instruction_master_readdatavalid                                              (cpu_instruction_master_readdatavalid),
      .cpu_instruction_master_requests_custom_dma_burst_1_upstream                       (cpu_instruction_master_requests_custom_dma_burst_1_upstream),
      .cpu_instruction_master_requests_custom_dma_burst_3_upstream                       (cpu_instruction_master_requests_custom_dma_burst_3_upstream),
      .cpu_instruction_master_waitrequest                                                (cpu_instruction_master_waitrequest),
      .custom_dma_burst_1_upstream_readdata_from_sa                                      (custom_dma_burst_1_upstream_readdata_from_sa),
      .custom_dma_burst_1_upstream_waitrequest_from_sa                                   (custom_dma_burst_1_upstream_waitrequest_from_sa),
      .custom_dma_burst_3_upstream_readdata_from_sa                                      (custom_dma_burst_3_upstream_readdata_from_sa),
      .custom_dma_burst_3_upstream_waitrequest_from_sa                                   (custom_dma_burst_3_upstream_waitrequest_from_sa),
      .d1_custom_dma_burst_1_upstream_end_xfer                                           (d1_custom_dma_burst_1_upstream_end_xfer),
      .d1_custom_dma_burst_3_upstream_end_xfer                                           (d1_custom_dma_burst_3_upstream_end_xfer),
      .reset_n                                                                           (system_clk_reset_n)
    );

  cpu the_cpu
    (
      .clk                                   (system_clk),
      .d_address                             (cpu_data_master_address),
      .d_burstcount                          (cpu_data_master_burstcount),
      .d_byteenable                          (cpu_data_master_byteenable),
      .d_irq                                 (cpu_data_master_irq),
      .d_read                                (cpu_data_master_read),
      .d_readdata                            (cpu_data_master_readdata),
      .d_readdatavalid                       (cpu_data_master_readdatavalid),
      .d_waitrequest                         (cpu_data_master_waitrequest),
      .d_write                               (cpu_data_master_write),
      .d_writedata                           (cpu_data_master_writedata),
      .i_address                             (cpu_instruction_master_address),
      .i_burstcount                          (cpu_instruction_master_burstcount),
      .i_read                                (cpu_instruction_master_read),
      .i_readdata                            (cpu_instruction_master_readdata),
      .i_readdatavalid                       (cpu_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_jtag_debug_module_byteenable),
      .jtag_debug_module_debugaccess         (cpu_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_jtag_debug_module_readdata),
      .jtag_debug_module_resetrequest        (cpu_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_jtag_debug_module_writedata),
      .reset_n                               (cpu_jtag_debug_module_reset_n)
    );

  custom_dma_burst_0_upstream_arbitrator the_custom_dma_burst_0_upstream
    (
      .clk                                                                        (system_clk),
      .cpu_data_master_address_to_slave                                           (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                 (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                 (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                (cpu_data_master_debugaccess),
      .cpu_data_master_granted_custom_dma_burst_0_upstream                        (cpu_data_master_granted_custom_dma_burst_0_upstream),
      .cpu_data_master_latency_counter                                            (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_custom_dma_burst_0_upstream              (cpu_data_master_qualified_request_custom_dma_burst_0_upstream),
      .cpu_data_master_read                                                       (cpu_data_master_read),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register),
      .cpu_data_master_requests_custom_dma_burst_0_upstream                       (cpu_data_master_requests_custom_dma_burst_0_upstream),
      .cpu_data_master_write                                                      (cpu_data_master_write),
      .cpu_data_master_writedata                                                  (cpu_data_master_writedata),
      .custom_dma_burst_0_upstream_address                                        (custom_dma_burst_0_upstream_address),
      .custom_dma_burst_0_upstream_burstcount                                     (custom_dma_burst_0_upstream_burstcount),
      .custom_dma_burst_0_upstream_byteaddress                                    (custom_dma_burst_0_upstream_byteaddress),
      .custom_dma_burst_0_upstream_byteenable                                     (custom_dma_burst_0_upstream_byteenable),
      .custom_dma_burst_0_upstream_debugaccess                                    (custom_dma_burst_0_upstream_debugaccess),
      .custom_dma_burst_0_upstream_read                                           (custom_dma_burst_0_upstream_read),
      .custom_dma_burst_0_upstream_readdata                                       (custom_dma_burst_0_upstream_readdata),
      .custom_dma_burst_0_upstream_readdata_from_sa                               (custom_dma_burst_0_upstream_readdata_from_sa),
      .custom_dma_burst_0_upstream_readdatavalid                                  (custom_dma_burst_0_upstream_readdatavalid),
      .custom_dma_burst_0_upstream_waitrequest                                    (custom_dma_burst_0_upstream_waitrequest),
      .custom_dma_burst_0_upstream_waitrequest_from_sa                            (custom_dma_burst_0_upstream_waitrequest_from_sa),
      .custom_dma_burst_0_upstream_write                                          (custom_dma_burst_0_upstream_write),
      .custom_dma_burst_0_upstream_writedata                                      (custom_dma_burst_0_upstream_writedata),
      .d1_custom_dma_burst_0_upstream_end_xfer                                    (d1_custom_dma_burst_0_upstream_end_xfer),
      .reset_n                                                                    (system_clk_reset_n)
    );

  custom_dma_burst_0_downstream_arbitrator the_custom_dma_burst_0_downstream
    (
      .clk                                                          (system_clk),
      .custom_dma_burst_0_downstream_address                        (custom_dma_burst_0_downstream_address),
      .custom_dma_burst_0_downstream_address_to_slave               (custom_dma_burst_0_downstream_address_to_slave),
      .custom_dma_burst_0_downstream_burstcount                     (custom_dma_burst_0_downstream_burstcount),
      .custom_dma_burst_0_downstream_byteenable                     (custom_dma_burst_0_downstream_byteenable),
      .custom_dma_burst_0_downstream_granted_ext_ssram_s1           (custom_dma_burst_0_downstream_granted_ext_ssram_s1),
      .custom_dma_burst_0_downstream_latency_counter                (custom_dma_burst_0_downstream_latency_counter),
      .custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 (custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1),
      .custom_dma_burst_0_downstream_read                           (custom_dma_burst_0_downstream_read),
      .custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1   (custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1),
      .custom_dma_burst_0_downstream_readdata                       (custom_dma_burst_0_downstream_readdata),
      .custom_dma_burst_0_downstream_readdatavalid                  (custom_dma_burst_0_downstream_readdatavalid),
      .custom_dma_burst_0_downstream_requests_ext_ssram_s1          (custom_dma_burst_0_downstream_requests_ext_ssram_s1),
      .custom_dma_burst_0_downstream_reset_n                        (custom_dma_burst_0_downstream_reset_n),
      .custom_dma_burst_0_downstream_waitrequest                    (custom_dma_burst_0_downstream_waitrequest),
      .custom_dma_burst_0_downstream_write                          (custom_dma_burst_0_downstream_write),
      .custom_dma_burst_0_downstream_writedata                      (custom_dma_burst_0_downstream_writedata),
      .d1_ext_ssram_bus_avalon_slave_end_xfer                       (d1_ext_ssram_bus_avalon_slave_end_xfer),
      .incoming_ext_ssram_bus_data                                  (incoming_ext_ssram_bus_data),
      .reset_n                                                      (system_clk_reset_n)
    );

  custom_dma_burst_0 the_custom_dma_burst_0
    (
      .clk                             (system_clk),
      .downstream_readdata             (custom_dma_burst_0_downstream_readdata),
      .downstream_readdatavalid        (custom_dma_burst_0_downstream_readdatavalid),
      .downstream_waitrequest          (custom_dma_burst_0_downstream_waitrequest),
      .reg_downstream_address          (custom_dma_burst_0_downstream_address),
      .reg_downstream_arbitrationshare (custom_dma_burst_0_downstream_arbitrationshare),
      .reg_downstream_burstcount       (custom_dma_burst_0_downstream_burstcount),
      .reg_downstream_byteenable       (custom_dma_burst_0_downstream_byteenable),
      .reg_downstream_debugaccess      (custom_dma_burst_0_downstream_debugaccess),
      .reg_downstream_nativeaddress    (custom_dma_burst_0_downstream_nativeaddress),
      .reg_downstream_read             (custom_dma_burst_0_downstream_read),
      .reg_downstream_write            (custom_dma_burst_0_downstream_write),
      .reg_downstream_writedata        (custom_dma_burst_0_downstream_writedata),
      .reset_n                         (custom_dma_burst_0_downstream_reset_n),
      .upstream_address                (custom_dma_burst_0_upstream_byteaddress),
      .upstream_burstcount             (custom_dma_burst_0_upstream_burstcount),
      .upstream_byteenable             (custom_dma_burst_0_upstream_byteenable),
      .upstream_debugaccess            (custom_dma_burst_0_upstream_debugaccess),
      .upstream_nativeaddress          (custom_dma_burst_0_upstream_address),
      .upstream_read                   (custom_dma_burst_0_upstream_read),
      .upstream_readdata               (custom_dma_burst_0_upstream_readdata),
      .upstream_readdatavalid          (custom_dma_burst_0_upstream_readdatavalid),
      .upstream_waitrequest            (custom_dma_burst_0_upstream_waitrequest),
      .upstream_write                  (custom_dma_burst_0_upstream_write),
      .upstream_writedata              (custom_dma_burst_0_upstream_writedata)
    );

  custom_dma_burst_1_upstream_arbitrator the_custom_dma_burst_1_upstream
    (
      .clk                                                                               (system_clk),
      .cpu_instruction_master_address_to_slave                                           (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                 (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_custom_dma_burst_1_upstream                        (cpu_instruction_master_granted_custom_dma_burst_1_upstream),
      .cpu_instruction_master_latency_counter                                            (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream              (cpu_instruction_master_qualified_request_custom_dma_burst_1_upstream),
      .cpu_instruction_master_read                                                       (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream                (cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register),
      .cpu_instruction_master_requests_custom_dma_burst_1_upstream                       (cpu_instruction_master_requests_custom_dma_burst_1_upstream),
      .custom_dma_burst_1_upstream_address                                               (custom_dma_burst_1_upstream_address),
      .custom_dma_burst_1_upstream_byteaddress                                           (custom_dma_burst_1_upstream_byteaddress),
      .custom_dma_burst_1_upstream_byteenable                                            (custom_dma_burst_1_upstream_byteenable),
      .custom_dma_burst_1_upstream_debugaccess                                           (custom_dma_burst_1_upstream_debugaccess),
      .custom_dma_burst_1_upstream_read                                                  (custom_dma_burst_1_upstream_read),
      .custom_dma_burst_1_upstream_readdata                                              (custom_dma_burst_1_upstream_readdata),
      .custom_dma_burst_1_upstream_readdata_from_sa                                      (custom_dma_burst_1_upstream_readdata_from_sa),
      .custom_dma_burst_1_upstream_readdatavalid                                         (custom_dma_burst_1_upstream_readdatavalid),
      .custom_dma_burst_1_upstream_waitrequest                                           (custom_dma_burst_1_upstream_waitrequest),
      .custom_dma_burst_1_upstream_waitrequest_from_sa                                   (custom_dma_burst_1_upstream_waitrequest_from_sa),
      .custom_dma_burst_1_upstream_write                                                 (custom_dma_burst_1_upstream_write),
      .d1_custom_dma_burst_1_upstream_end_xfer                                           (d1_custom_dma_burst_1_upstream_end_xfer),
      .reset_n                                                                           (system_clk_reset_n)
    );

  custom_dma_burst_1_downstream_arbitrator the_custom_dma_burst_1_downstream
    (
      .clk                                                                             (system_clk),
      .custom_dma_burst_1_downstream_address                                           (custom_dma_burst_1_downstream_address),
      .custom_dma_burst_1_downstream_address_to_slave                                  (custom_dma_burst_1_downstream_address_to_slave),
      .custom_dma_burst_1_downstream_burstcount                                        (custom_dma_burst_1_downstream_burstcount),
      .custom_dma_burst_1_downstream_byteenable                                        (custom_dma_burst_1_downstream_byteenable),
      .custom_dma_burst_1_downstream_granted_pipeline_bridge_s1                        (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_latency_counter                                   (custom_dma_burst_1_downstream_latency_counter),
      .custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1              (custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_read                                              (custom_dma_burst_1_downstream_read),
      .custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1                (custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register (custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register),
      .custom_dma_burst_1_downstream_readdata                                          (custom_dma_burst_1_downstream_readdata),
      .custom_dma_burst_1_downstream_readdatavalid                                     (custom_dma_burst_1_downstream_readdatavalid),
      .custom_dma_burst_1_downstream_requests_pipeline_bridge_s1                       (custom_dma_burst_1_downstream_requests_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_reset_n                                           (custom_dma_burst_1_downstream_reset_n),
      .custom_dma_burst_1_downstream_waitrequest                                       (custom_dma_burst_1_downstream_waitrequest),
      .custom_dma_burst_1_downstream_write                                             (custom_dma_burst_1_downstream_write),
      .custom_dma_burst_1_downstream_writedata                                         (custom_dma_burst_1_downstream_writedata),
      .d1_pipeline_bridge_s1_end_xfer                                                  (d1_pipeline_bridge_s1_end_xfer),
      .pipeline_bridge_s1_readdata_from_sa                                             (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_waitrequest_from_sa                                          (pipeline_bridge_s1_waitrequest_from_sa),
      .reset_n                                                                         (system_clk_reset_n)
    );

  custom_dma_burst_1 the_custom_dma_burst_1
    (
      .clk                             (system_clk),
      .downstream_readdata             (custom_dma_burst_1_downstream_readdata),
      .downstream_readdatavalid        (custom_dma_burst_1_downstream_readdatavalid),
      .downstream_waitrequest          (custom_dma_burst_1_downstream_waitrequest),
      .reg_downstream_address          (custom_dma_burst_1_downstream_address),
      .reg_downstream_arbitrationshare (custom_dma_burst_1_downstream_arbitrationshare),
      .reg_downstream_burstcount       (custom_dma_burst_1_downstream_burstcount),
      .reg_downstream_byteenable       (custom_dma_burst_1_downstream_byteenable),
      .reg_downstream_debugaccess      (custom_dma_burst_1_downstream_debugaccess),
      .reg_downstream_nativeaddress    (custom_dma_burst_1_downstream_nativeaddress),
      .reg_downstream_read             (custom_dma_burst_1_downstream_read),
      .reg_downstream_write            (custom_dma_burst_1_downstream_write),
      .reg_downstream_writedata        (custom_dma_burst_1_downstream_writedata),
      .reset_n                         (custom_dma_burst_1_downstream_reset_n),
      .upstream_address                (custom_dma_burst_1_upstream_byteaddress),
      .upstream_byteenable             (custom_dma_burst_1_upstream_byteenable),
      .upstream_debugaccess            (custom_dma_burst_1_upstream_debugaccess),
      .upstream_nativeaddress          (custom_dma_burst_1_upstream_address),
      .upstream_read                   (custom_dma_burst_1_upstream_read),
      .upstream_readdata               (custom_dma_burst_1_upstream_readdata),
      .upstream_readdatavalid          (custom_dma_burst_1_upstream_readdatavalid),
      .upstream_waitrequest            (custom_dma_burst_1_upstream_waitrequest),
      .upstream_write                  (custom_dma_burst_1_upstream_write),
      .upstream_writedata              (custom_dma_burst_1_upstream_writedata)
    );

  custom_dma_burst_2_upstream_arbitrator the_custom_dma_burst_2_upstream
    (
      .clk                                                                        (system_clk),
      .cpu_data_master_address_to_slave                                           (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                 (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                 (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                (cpu_data_master_debugaccess),
      .cpu_data_master_granted_custom_dma_burst_2_upstream                        (cpu_data_master_granted_custom_dma_burst_2_upstream),
      .cpu_data_master_latency_counter                                            (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_custom_dma_burst_2_upstream              (cpu_data_master_qualified_request_custom_dma_burst_2_upstream),
      .cpu_data_master_read                                                       (cpu_data_master_read),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register),
      .cpu_data_master_requests_custom_dma_burst_2_upstream                       (cpu_data_master_requests_custom_dma_burst_2_upstream),
      .cpu_data_master_write                                                      (cpu_data_master_write),
      .cpu_data_master_writedata                                                  (cpu_data_master_writedata),
      .custom_dma_burst_2_upstream_address                                        (custom_dma_burst_2_upstream_address),
      .custom_dma_burst_2_upstream_burstcount                                     (custom_dma_burst_2_upstream_burstcount),
      .custom_dma_burst_2_upstream_byteaddress                                    (custom_dma_burst_2_upstream_byteaddress),
      .custom_dma_burst_2_upstream_byteenable                                     (custom_dma_burst_2_upstream_byteenable),
      .custom_dma_burst_2_upstream_debugaccess                                    (custom_dma_burst_2_upstream_debugaccess),
      .custom_dma_burst_2_upstream_read                                           (custom_dma_burst_2_upstream_read),
      .custom_dma_burst_2_upstream_readdata                                       (custom_dma_burst_2_upstream_readdata),
      .custom_dma_burst_2_upstream_readdata_from_sa                               (custom_dma_burst_2_upstream_readdata_from_sa),
      .custom_dma_burst_2_upstream_readdatavalid                                  (custom_dma_burst_2_upstream_readdatavalid),
      .custom_dma_burst_2_upstream_waitrequest                                    (custom_dma_burst_2_upstream_waitrequest),
      .custom_dma_burst_2_upstream_waitrequest_from_sa                            (custom_dma_burst_2_upstream_waitrequest_from_sa),
      .custom_dma_burst_2_upstream_write                                          (custom_dma_burst_2_upstream_write),
      .custom_dma_burst_2_upstream_writedata                                      (custom_dma_burst_2_upstream_writedata),
      .d1_custom_dma_burst_2_upstream_end_xfer                                    (d1_custom_dma_burst_2_upstream_end_xfer),
      .reset_n                                                                    (system_clk_reset_n)
    );

  custom_dma_burst_2_downstream_arbitrator the_custom_dma_burst_2_downstream
    (
      .clk                                                                             (system_clk),
      .custom_dma_burst_2_downstream_address                                           (custom_dma_burst_2_downstream_address),
      .custom_dma_burst_2_downstream_address_to_slave                                  (custom_dma_burst_2_downstream_address_to_slave),
      .custom_dma_burst_2_downstream_burstcount                                        (custom_dma_burst_2_downstream_burstcount),
      .custom_dma_burst_2_downstream_byteenable                                        (custom_dma_burst_2_downstream_byteenable),
      .custom_dma_burst_2_downstream_granted_pipeline_bridge_s1                        (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_latency_counter                                   (custom_dma_burst_2_downstream_latency_counter),
      .custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1              (custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_read                                              (custom_dma_burst_2_downstream_read),
      .custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1                (custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register (custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register),
      .custom_dma_burst_2_downstream_readdata                                          (custom_dma_burst_2_downstream_readdata),
      .custom_dma_burst_2_downstream_readdatavalid                                     (custom_dma_burst_2_downstream_readdatavalid),
      .custom_dma_burst_2_downstream_requests_pipeline_bridge_s1                       (custom_dma_burst_2_downstream_requests_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_reset_n                                           (custom_dma_burst_2_downstream_reset_n),
      .custom_dma_burst_2_downstream_waitrequest                                       (custom_dma_burst_2_downstream_waitrequest),
      .custom_dma_burst_2_downstream_write                                             (custom_dma_burst_2_downstream_write),
      .custom_dma_burst_2_downstream_writedata                                         (custom_dma_burst_2_downstream_writedata),
      .d1_pipeline_bridge_s1_end_xfer                                                  (d1_pipeline_bridge_s1_end_xfer),
      .pipeline_bridge_s1_readdata_from_sa                                             (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_waitrequest_from_sa                                          (pipeline_bridge_s1_waitrequest_from_sa),
      .reset_n                                                                         (system_clk_reset_n)
    );

  custom_dma_burst_2 the_custom_dma_burst_2
    (
      .clk                             (system_clk),
      .downstream_readdata             (custom_dma_burst_2_downstream_readdata),
      .downstream_readdatavalid        (custom_dma_burst_2_downstream_readdatavalid),
      .downstream_waitrequest          (custom_dma_burst_2_downstream_waitrequest),
      .reg_downstream_address          (custom_dma_burst_2_downstream_address),
      .reg_downstream_arbitrationshare (custom_dma_burst_2_downstream_arbitrationshare),
      .reg_downstream_burstcount       (custom_dma_burst_2_downstream_burstcount),
      .reg_downstream_byteenable       (custom_dma_burst_2_downstream_byteenable),
      .reg_downstream_debugaccess      (custom_dma_burst_2_downstream_debugaccess),
      .reg_downstream_nativeaddress    (custom_dma_burst_2_downstream_nativeaddress),
      .reg_downstream_read             (custom_dma_burst_2_downstream_read),
      .reg_downstream_write            (custom_dma_burst_2_downstream_write),
      .reg_downstream_writedata        (custom_dma_burst_2_downstream_writedata),
      .reset_n                         (custom_dma_burst_2_downstream_reset_n),
      .upstream_address                (custom_dma_burst_2_upstream_byteaddress),
      .upstream_burstcount             (custom_dma_burst_2_upstream_burstcount),
      .upstream_byteenable             (custom_dma_burst_2_upstream_byteenable),
      .upstream_debugaccess            (custom_dma_burst_2_upstream_debugaccess),
      .upstream_nativeaddress          (custom_dma_burst_2_upstream_address),
      .upstream_read                   (custom_dma_burst_2_upstream_read),
      .upstream_readdata               (custom_dma_burst_2_upstream_readdata),
      .upstream_readdatavalid          (custom_dma_burst_2_upstream_readdatavalid),
      .upstream_waitrequest            (custom_dma_burst_2_upstream_waitrequest),
      .upstream_write                  (custom_dma_burst_2_upstream_write),
      .upstream_writedata              (custom_dma_burst_2_upstream_writedata)
    );

  custom_dma_burst_3_upstream_arbitrator the_custom_dma_burst_3_upstream
    (
      .clk                                                                               (system_clk),
      .cpu_instruction_master_address_to_slave                                           (cpu_instruction_master_address_to_slave),
      .cpu_instruction_master_burstcount                                                 (cpu_instruction_master_burstcount),
      .cpu_instruction_master_granted_custom_dma_burst_3_upstream                        (cpu_instruction_master_granted_custom_dma_burst_3_upstream),
      .cpu_instruction_master_latency_counter                                            (cpu_instruction_master_latency_counter),
      .cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream              (cpu_instruction_master_qualified_request_custom_dma_burst_3_upstream),
      .cpu_instruction_master_read                                                       (cpu_instruction_master_read),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_1_upstream_shift_register),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream                (cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream),
      .cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register (cpu_instruction_master_read_data_valid_custom_dma_burst_3_upstream_shift_register),
      .cpu_instruction_master_requests_custom_dma_burst_3_upstream                       (cpu_instruction_master_requests_custom_dma_burst_3_upstream),
      .custom_dma_burst_3_upstream_address                                               (custom_dma_burst_3_upstream_address),
      .custom_dma_burst_3_upstream_byteaddress                                           (custom_dma_burst_3_upstream_byteaddress),
      .custom_dma_burst_3_upstream_byteenable                                            (custom_dma_burst_3_upstream_byteenable),
      .custom_dma_burst_3_upstream_debugaccess                                           (custom_dma_burst_3_upstream_debugaccess),
      .custom_dma_burst_3_upstream_read                                                  (custom_dma_burst_3_upstream_read),
      .custom_dma_burst_3_upstream_readdata                                              (custom_dma_burst_3_upstream_readdata),
      .custom_dma_burst_3_upstream_readdata_from_sa                                      (custom_dma_burst_3_upstream_readdata_from_sa),
      .custom_dma_burst_3_upstream_readdatavalid                                         (custom_dma_burst_3_upstream_readdatavalid),
      .custom_dma_burst_3_upstream_waitrequest                                           (custom_dma_burst_3_upstream_waitrequest),
      .custom_dma_burst_3_upstream_waitrequest_from_sa                                   (custom_dma_burst_3_upstream_waitrequest_from_sa),
      .custom_dma_burst_3_upstream_write                                                 (custom_dma_burst_3_upstream_write),
      .d1_custom_dma_burst_3_upstream_end_xfer                                           (d1_custom_dma_burst_3_upstream_end_xfer),
      .reset_n                                                                           (system_clk_reset_n)
    );

  custom_dma_burst_3_downstream_arbitrator the_custom_dma_burst_3_downstream
    (
      .clk                                                                       (system_clk),
      .custom_dma_burst_3_downstream_address                                     (custom_dma_burst_3_downstream_address),
      .custom_dma_burst_3_downstream_address_to_slave                            (custom_dma_burst_3_downstream_address_to_slave),
      .custom_dma_burst_3_downstream_burstcount                                  (custom_dma_burst_3_downstream_burstcount),
      .custom_dma_burst_3_downstream_byteenable                                  (custom_dma_burst_3_downstream_byteenable),
      .custom_dma_burst_3_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_3_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_latency_counter                             (custom_dma_burst_3_downstream_latency_counter),
      .custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_read                                        (custom_dma_burst_3_downstream_read),
      .custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_3_downstream_readdata                                    (custom_dma_burst_3_downstream_readdata),
      .custom_dma_burst_3_downstream_readdatavalid                               (custom_dma_burst_3_downstream_readdatavalid),
      .custom_dma_burst_3_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_3_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_reset_n                                     (custom_dma_burst_3_downstream_reset_n),
      .custom_dma_burst_3_downstream_waitrequest                                 (custom_dma_burst_3_downstream_waitrequest),
      .custom_dma_burst_3_downstream_write                                       (custom_dma_burst_3_downstream_write),
      .custom_dma_burst_3_downstream_writedata                                   (custom_dma_burst_3_downstream_writedata),
      .d1_ddr_sdram_s1_end_xfer                                                  (d1_ddr_sdram_s1_end_xfer),
      .ddr_sdram_s1_readdata_from_sa                                             (ddr_sdram_s1_readdata_from_sa),
      .ddr_sdram_s1_waitrequest_n_from_sa                                        (ddr_sdram_s1_waitrequest_n_from_sa),
      .reset_n                                                                   (system_clk_reset_n)
    );

  custom_dma_burst_3 the_custom_dma_burst_3
    (
      .clk                             (system_clk),
      .downstream_readdata             (custom_dma_burst_3_downstream_readdata),
      .downstream_readdatavalid        (custom_dma_burst_3_downstream_readdatavalid),
      .downstream_waitrequest          (custom_dma_burst_3_downstream_waitrequest),
      .reg_downstream_address          (custom_dma_burst_3_downstream_address),
      .reg_downstream_arbitrationshare (custom_dma_burst_3_downstream_arbitrationshare),
      .reg_downstream_burstcount       (custom_dma_burst_3_downstream_burstcount),
      .reg_downstream_byteenable       (custom_dma_burst_3_downstream_byteenable),
      .reg_downstream_debugaccess      (custom_dma_burst_3_downstream_debugaccess),
      .reg_downstream_nativeaddress    (custom_dma_burst_3_downstream_nativeaddress),
      .reg_downstream_read             (custom_dma_burst_3_downstream_read),
      .reg_downstream_write            (custom_dma_burst_3_downstream_write),
      .reg_downstream_writedata        (custom_dma_burst_3_downstream_writedata),
      .reset_n                         (custom_dma_burst_3_downstream_reset_n),
      .upstream_address                (custom_dma_burst_3_upstream_byteaddress),
      .upstream_byteenable             (custom_dma_burst_3_upstream_byteenable),
      .upstream_debugaccess            (custom_dma_burst_3_upstream_debugaccess),
      .upstream_nativeaddress          (custom_dma_burst_3_upstream_address),
      .upstream_read                   (custom_dma_burst_3_upstream_read),
      .upstream_readdata               (custom_dma_burst_3_upstream_readdata),
      .upstream_readdatavalid          (custom_dma_burst_3_upstream_readdatavalid),
      .upstream_waitrequest            (custom_dma_burst_3_upstream_waitrequest),
      .upstream_write                  (custom_dma_burst_3_upstream_write),
      .upstream_writedata              (custom_dma_burst_3_upstream_writedata)
    );

  custom_dma_burst_4_upstream_arbitrator the_custom_dma_burst_4_upstream
    (
      .clk                                                                        (system_clk),
      .cpu_data_master_address_to_slave                                           (cpu_data_master_address_to_slave),
      .cpu_data_master_burstcount                                                 (cpu_data_master_burstcount),
      .cpu_data_master_byteenable                                                 (cpu_data_master_byteenable),
      .cpu_data_master_debugaccess                                                (cpu_data_master_debugaccess),
      .cpu_data_master_granted_custom_dma_burst_4_upstream                        (cpu_data_master_granted_custom_dma_burst_4_upstream),
      .cpu_data_master_latency_counter                                            (cpu_data_master_latency_counter),
      .cpu_data_master_qualified_request_custom_dma_burst_4_upstream              (cpu_data_master_qualified_request_custom_dma_burst_4_upstream),
      .cpu_data_master_read                                                       (cpu_data_master_read),
      .cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_0_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_2_upstream_shift_register),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream                (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream),
      .cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register (cpu_data_master_read_data_valid_custom_dma_burst_4_upstream_shift_register),
      .cpu_data_master_requests_custom_dma_burst_4_upstream                       (cpu_data_master_requests_custom_dma_burst_4_upstream),
      .cpu_data_master_write                                                      (cpu_data_master_write),
      .cpu_data_master_writedata                                                  (cpu_data_master_writedata),
      .custom_dma_burst_4_upstream_address                                        (custom_dma_burst_4_upstream_address),
      .custom_dma_burst_4_upstream_burstcount                                     (custom_dma_burst_4_upstream_burstcount),
      .custom_dma_burst_4_upstream_byteaddress                                    (custom_dma_burst_4_upstream_byteaddress),
      .custom_dma_burst_4_upstream_byteenable                                     (custom_dma_burst_4_upstream_byteenable),
      .custom_dma_burst_4_upstream_debugaccess                                    (custom_dma_burst_4_upstream_debugaccess),
      .custom_dma_burst_4_upstream_read                                           (custom_dma_burst_4_upstream_read),
      .custom_dma_burst_4_upstream_readdata                                       (custom_dma_burst_4_upstream_readdata),
      .custom_dma_burst_4_upstream_readdata_from_sa                               (custom_dma_burst_4_upstream_readdata_from_sa),
      .custom_dma_burst_4_upstream_readdatavalid                                  (custom_dma_burst_4_upstream_readdatavalid),
      .custom_dma_burst_4_upstream_waitrequest                                    (custom_dma_burst_4_upstream_waitrequest),
      .custom_dma_burst_4_upstream_waitrequest_from_sa                            (custom_dma_burst_4_upstream_waitrequest_from_sa),
      .custom_dma_burst_4_upstream_write                                          (custom_dma_burst_4_upstream_write),
      .custom_dma_burst_4_upstream_writedata                                      (custom_dma_burst_4_upstream_writedata),
      .d1_custom_dma_burst_4_upstream_end_xfer                                    (d1_custom_dma_burst_4_upstream_end_xfer),
      .reset_n                                                                    (system_clk_reset_n)
    );

  custom_dma_burst_4_downstream_arbitrator the_custom_dma_burst_4_downstream
    (
      .clk                                                                       (system_clk),
      .custom_dma_burst_4_downstream_address                                     (custom_dma_burst_4_downstream_address),
      .custom_dma_burst_4_downstream_address_to_slave                            (custom_dma_burst_4_downstream_address_to_slave),
      .custom_dma_burst_4_downstream_burstcount                                  (custom_dma_burst_4_downstream_burstcount),
      .custom_dma_burst_4_downstream_byteenable                                  (custom_dma_burst_4_downstream_byteenable),
      .custom_dma_burst_4_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_4_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_latency_counter                             (custom_dma_burst_4_downstream_latency_counter),
      .custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_read                                        (custom_dma_burst_4_downstream_read),
      .custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_4_downstream_readdata                                    (custom_dma_burst_4_downstream_readdata),
      .custom_dma_burst_4_downstream_readdatavalid                               (custom_dma_burst_4_downstream_readdatavalid),
      .custom_dma_burst_4_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_4_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_reset_n                                     (custom_dma_burst_4_downstream_reset_n),
      .custom_dma_burst_4_downstream_waitrequest                                 (custom_dma_burst_4_downstream_waitrequest),
      .custom_dma_burst_4_downstream_write                                       (custom_dma_burst_4_downstream_write),
      .custom_dma_burst_4_downstream_writedata                                   (custom_dma_burst_4_downstream_writedata),
      .d1_ddr_sdram_s1_end_xfer                                                  (d1_ddr_sdram_s1_end_xfer),
      .ddr_sdram_s1_readdata_from_sa                                             (ddr_sdram_s1_readdata_from_sa),
      .ddr_sdram_s1_waitrequest_n_from_sa                                        (ddr_sdram_s1_waitrequest_n_from_sa),
      .reset_n                                                                   (system_clk_reset_n)
    );

  custom_dma_burst_4 the_custom_dma_burst_4
    (
      .clk                             (system_clk),
      .downstream_readdata             (custom_dma_burst_4_downstream_readdata),
      .downstream_readdatavalid        (custom_dma_burst_4_downstream_readdatavalid),
      .downstream_waitrequest          (custom_dma_burst_4_downstream_waitrequest),
      .reg_downstream_address          (custom_dma_burst_4_downstream_address),
      .reg_downstream_arbitrationshare (custom_dma_burst_4_downstream_arbitrationshare),
      .reg_downstream_burstcount       (custom_dma_burst_4_downstream_burstcount),
      .reg_downstream_byteenable       (custom_dma_burst_4_downstream_byteenable),
      .reg_downstream_debugaccess      (custom_dma_burst_4_downstream_debugaccess),
      .reg_downstream_nativeaddress    (custom_dma_burst_4_downstream_nativeaddress),
      .reg_downstream_read             (custom_dma_burst_4_downstream_read),
      .reg_downstream_write            (custom_dma_burst_4_downstream_write),
      .reg_downstream_writedata        (custom_dma_burst_4_downstream_writedata),
      .reset_n                         (custom_dma_burst_4_downstream_reset_n),
      .upstream_address                (custom_dma_burst_4_upstream_byteaddress),
      .upstream_burstcount             (custom_dma_burst_4_upstream_burstcount),
      .upstream_byteenable             (custom_dma_burst_4_upstream_byteenable),
      .upstream_debugaccess            (custom_dma_burst_4_upstream_debugaccess),
      .upstream_nativeaddress          (custom_dma_burst_4_upstream_address),
      .upstream_read                   (custom_dma_burst_4_upstream_read),
      .upstream_readdata               (custom_dma_burst_4_upstream_readdata),
      .upstream_readdatavalid          (custom_dma_burst_4_upstream_readdatavalid),
      .upstream_waitrequest            (custom_dma_burst_4_upstream_waitrequest),
      .upstream_write                  (custom_dma_burst_4_upstream_write),
      .upstream_writedata              (custom_dma_burst_4_upstream_writedata)
    );

  custom_dma_burst_5_upstream_arbitrator the_custom_dma_burst_5_upstream
    (
      .clk                                                                (system_clk),
      .custom_dma_burst_5_upstream_address                                (custom_dma_burst_5_upstream_address),
      .custom_dma_burst_5_upstream_burstcount                             (custom_dma_burst_5_upstream_burstcount),
      .custom_dma_burst_5_upstream_byteaddress                            (custom_dma_burst_5_upstream_byteaddress),
      .custom_dma_burst_5_upstream_byteenable                             (custom_dma_burst_5_upstream_byteenable),
      .custom_dma_burst_5_upstream_debugaccess                            (custom_dma_burst_5_upstream_debugaccess),
      .custom_dma_burst_5_upstream_read                                   (custom_dma_burst_5_upstream_read),
      .custom_dma_burst_5_upstream_readdata                               (custom_dma_burst_5_upstream_readdata),
      .custom_dma_burst_5_upstream_readdata_from_sa                       (custom_dma_burst_5_upstream_readdata_from_sa),
      .custom_dma_burst_5_upstream_readdatavalid                          (custom_dma_burst_5_upstream_readdatavalid),
      .custom_dma_burst_5_upstream_readdatavalid_from_sa                  (custom_dma_burst_5_upstream_readdatavalid_from_sa),
      .custom_dma_burst_5_upstream_waitrequest                            (custom_dma_burst_5_upstream_waitrequest),
      .custom_dma_burst_5_upstream_waitrequest_from_sa                    (custom_dma_burst_5_upstream_waitrequest_from_sa),
      .custom_dma_burst_5_upstream_write                                  (custom_dma_burst_5_upstream_write),
      .custom_dma_burst_5_upstream_writedata                              (custom_dma_burst_5_upstream_writedata),
      .d1_custom_dma_burst_5_upstream_end_xfer                            (d1_custom_dma_burst_5_upstream_end_xfer),
      .fir_dma_write_master_address_to_slave                              (fir_dma_write_master_address_to_slave),
      .fir_dma_write_master_burstcount                                    (fir_dma_write_master_burstcount),
      .fir_dma_write_master_byteenable                                    (fir_dma_write_master_byteenable),
      .fir_dma_write_master_granted_custom_dma_burst_5_upstream           (fir_dma_write_master_granted_custom_dma_burst_5_upstream),
      .fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream (fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream),
      .fir_dma_write_master_requests_custom_dma_burst_5_upstream          (fir_dma_write_master_requests_custom_dma_burst_5_upstream),
      .fir_dma_write_master_write                                         (fir_dma_write_master_write),
      .fir_dma_write_master_writedata                                     (fir_dma_write_master_writedata),
      .reset_n                                                            (system_clk_reset_n)
    );

  custom_dma_burst_5_downstream_arbitrator the_custom_dma_burst_5_downstream
    (
      .clk                                                                       (system_clk),
      .custom_dma_burst_5_downstream_address                                     (custom_dma_burst_5_downstream_address),
      .custom_dma_burst_5_downstream_address_to_slave                            (custom_dma_burst_5_downstream_address_to_slave),
      .custom_dma_burst_5_downstream_burstcount                                  (custom_dma_burst_5_downstream_burstcount),
      .custom_dma_burst_5_downstream_byteenable                                  (custom_dma_burst_5_downstream_byteenable),
      .custom_dma_burst_5_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_5_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_latency_counter                             (custom_dma_burst_5_downstream_latency_counter),
      .custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_read                                        (custom_dma_burst_5_downstream_read),
      .custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_5_downstream_readdata                                    (custom_dma_burst_5_downstream_readdata),
      .custom_dma_burst_5_downstream_readdatavalid                               (custom_dma_burst_5_downstream_readdatavalid),
      .custom_dma_burst_5_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_5_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_reset_n                                     (custom_dma_burst_5_downstream_reset_n),
      .custom_dma_burst_5_downstream_waitrequest                                 (custom_dma_burst_5_downstream_waitrequest),
      .custom_dma_burst_5_downstream_write                                       (custom_dma_burst_5_downstream_write),
      .custom_dma_burst_5_downstream_writedata                                   (custom_dma_burst_5_downstream_writedata),
      .d1_ddr_sdram_s1_end_xfer                                                  (d1_ddr_sdram_s1_end_xfer),
      .ddr_sdram_s1_readdata_from_sa                                             (ddr_sdram_s1_readdata_from_sa),
      .ddr_sdram_s1_waitrequest_n_from_sa                                        (ddr_sdram_s1_waitrequest_n_from_sa),
      .reset_n                                                                   (system_clk_reset_n)
    );

  custom_dma_burst_5 the_custom_dma_burst_5
    (
      .clk                         (system_clk),
      .downstream_address          (custom_dma_burst_5_downstream_address),
      .downstream_arbitrationshare (custom_dma_burst_5_downstream_arbitrationshare),
      .downstream_burstcount       (custom_dma_burst_5_downstream_burstcount),
      .downstream_byteenable       (custom_dma_burst_5_downstream_byteenable),
      .downstream_debugaccess      (custom_dma_burst_5_downstream_debugaccess),
      .downstream_nativeaddress    (custom_dma_burst_5_downstream_nativeaddress),
      .downstream_read             (custom_dma_burst_5_downstream_read),
      .downstream_readdata         (custom_dma_burst_5_downstream_readdata),
      .downstream_readdatavalid    (custom_dma_burst_5_downstream_readdatavalid),
      .downstream_waitrequest      (custom_dma_burst_5_downstream_waitrequest),
      .downstream_write            (custom_dma_burst_5_downstream_write),
      .downstream_writedata        (custom_dma_burst_5_downstream_writedata),
      .reset_n                     (custom_dma_burst_5_downstream_reset_n),
      .upstream_address            (custom_dma_burst_5_upstream_byteaddress),
      .upstream_burstcount         (custom_dma_burst_5_upstream_burstcount),
      .upstream_byteenable         (custom_dma_burst_5_upstream_byteenable),
      .upstream_debugaccess        (custom_dma_burst_5_upstream_debugaccess),
      .upstream_nativeaddress      (custom_dma_burst_5_upstream_address),
      .upstream_read               (custom_dma_burst_5_upstream_read),
      .upstream_readdata           (custom_dma_burst_5_upstream_readdata),
      .upstream_readdatavalid      (custom_dma_burst_5_upstream_readdatavalid),
      .upstream_waitrequest        (custom_dma_burst_5_upstream_waitrequest),
      .upstream_write              (custom_dma_burst_5_upstream_write),
      .upstream_writedata          (custom_dma_burst_5_upstream_writedata)
    );

  custom_dma_clock_0_in_arbitrator the_custom_dma_clock_0_in
    (
      .clk                                                        (system_clk),
      .custom_dma_clock_0_in_address                              (custom_dma_clock_0_in_address),
      .custom_dma_clock_0_in_byteenable                           (custom_dma_clock_0_in_byteenable),
      .custom_dma_clock_0_in_endofpacket                          (custom_dma_clock_0_in_endofpacket),
      .custom_dma_clock_0_in_endofpacket_from_sa                  (custom_dma_clock_0_in_endofpacket_from_sa),
      .custom_dma_clock_0_in_nativeaddress                        (custom_dma_clock_0_in_nativeaddress),
      .custom_dma_clock_0_in_read                                 (custom_dma_clock_0_in_read),
      .custom_dma_clock_0_in_readdata                             (custom_dma_clock_0_in_readdata),
      .custom_dma_clock_0_in_readdata_from_sa                     (custom_dma_clock_0_in_readdata_from_sa),
      .custom_dma_clock_0_in_reset_n                              (custom_dma_clock_0_in_reset_n),
      .custom_dma_clock_0_in_waitrequest                          (custom_dma_clock_0_in_waitrequest),
      .custom_dma_clock_0_in_waitrequest_from_sa                  (custom_dma_clock_0_in_waitrequest_from_sa),
      .custom_dma_clock_0_in_write                                (custom_dma_clock_0_in_write),
      .custom_dma_clock_0_in_writedata                            (custom_dma_clock_0_in_writedata),
      .d1_custom_dma_clock_0_in_end_xfer                          (d1_custom_dma_clock_0_in_end_xfer),
      .pipeline_bridge_m1_address_to_slave                        (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                              (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                              (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                              (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_custom_dma_clock_0_in           (pipeline_bridge_m1_granted_custom_dma_clock_0_in),
      .pipeline_bridge_m1_latency_counter                         (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in (pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in),
      .pipeline_bridge_m1_read                                    (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in   (pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in),
      .pipeline_bridge_m1_requests_custom_dma_clock_0_in          (pipeline_bridge_m1_requests_custom_dma_clock_0_in),
      .pipeline_bridge_m1_write                                   (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                               (pipeline_bridge_m1_writedata),
      .reset_n                                                    (system_clk_reset_n)
    );

  custom_dma_clock_0_out_arbitrator the_custom_dma_clock_0_out
    (
      .clk                                             (external_clk),
      .custom_dma_clock_0_out_address                  (custom_dma_clock_0_out_address),
      .custom_dma_clock_0_out_address_to_slave         (custom_dma_clock_0_out_address_to_slave),
      .custom_dma_clock_0_out_byteenable               (custom_dma_clock_0_out_byteenable),
      .custom_dma_clock_0_out_granted_pll_s1           (custom_dma_clock_0_out_granted_pll_s1),
      .custom_dma_clock_0_out_qualified_request_pll_s1 (custom_dma_clock_0_out_qualified_request_pll_s1),
      .custom_dma_clock_0_out_read                     (custom_dma_clock_0_out_read),
      .custom_dma_clock_0_out_read_data_valid_pll_s1   (custom_dma_clock_0_out_read_data_valid_pll_s1),
      .custom_dma_clock_0_out_readdata                 (custom_dma_clock_0_out_readdata),
      .custom_dma_clock_0_out_requests_pll_s1          (custom_dma_clock_0_out_requests_pll_s1),
      .custom_dma_clock_0_out_reset_n                  (custom_dma_clock_0_out_reset_n),
      .custom_dma_clock_0_out_waitrequest              (custom_dma_clock_0_out_waitrequest),
      .custom_dma_clock_0_out_write                    (custom_dma_clock_0_out_write),
      .custom_dma_clock_0_out_writedata                (custom_dma_clock_0_out_writedata),
      .d1_pll_s1_end_xfer                              (d1_pll_s1_end_xfer),
      .pll_s1_readdata_from_sa                         (pll_s1_readdata_from_sa),
      .reset_n                                         (external_clk_reset_n)
    );

  custom_dma_clock_0 the_custom_dma_clock_0
    (
      .master_address       (custom_dma_clock_0_out_address),
      .master_byteenable    (custom_dma_clock_0_out_byteenable),
      .master_clk           (external_clk),
      .master_endofpacket   (custom_dma_clock_0_out_endofpacket),
      .master_nativeaddress (custom_dma_clock_0_out_nativeaddress),
      .master_read          (custom_dma_clock_0_out_read),
      .master_readdata      (custom_dma_clock_0_out_readdata),
      .master_reset_n       (custom_dma_clock_0_out_reset_n),
      .master_waitrequest   (custom_dma_clock_0_out_waitrequest),
      .master_write         (custom_dma_clock_0_out_write),
      .master_writedata     (custom_dma_clock_0_out_writedata),
      .slave_address        (custom_dma_clock_0_in_address),
      .slave_byteenable     (custom_dma_clock_0_in_byteenable),
      .slave_clk            (system_clk),
      .slave_endofpacket    (custom_dma_clock_0_in_endofpacket),
      .slave_nativeaddress  (custom_dma_clock_0_in_nativeaddress),
      .slave_read           (custom_dma_clock_0_in_read),
      .slave_readdata       (custom_dma_clock_0_in_readdata),
      .slave_reset_n        (custom_dma_clock_0_in_reset_n),
      .slave_waitrequest    (custom_dma_clock_0_in_waitrequest),
      .slave_write          (custom_dma_clock_0_in_write),
      .slave_writedata      (custom_dma_clock_0_in_writedata)
    );

  ddr_sdram_s1_arbitrator the_ddr_sdram_s1
    (
      .clk                                                                       (system_clk),
      .custom_dma_burst_3_downstream_address_to_slave                            (custom_dma_burst_3_downstream_address_to_slave),
      .custom_dma_burst_3_downstream_arbitrationshare                            (custom_dma_burst_3_downstream_arbitrationshare),
      .custom_dma_burst_3_downstream_burstcount                                  (custom_dma_burst_3_downstream_burstcount),
      .custom_dma_burst_3_downstream_byteenable                                  (custom_dma_burst_3_downstream_byteenable),
      .custom_dma_burst_3_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_3_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_latency_counter                             (custom_dma_burst_3_downstream_latency_counter),
      .custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_3_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_read                                        (custom_dma_burst_3_downstream_read),
      .custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_3_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_3_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_3_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_3_downstream_write                                       (custom_dma_burst_3_downstream_write),
      .custom_dma_burst_3_downstream_writedata                                   (custom_dma_burst_3_downstream_writedata),
      .custom_dma_burst_4_downstream_address_to_slave                            (custom_dma_burst_4_downstream_address_to_slave),
      .custom_dma_burst_4_downstream_arbitrationshare                            (custom_dma_burst_4_downstream_arbitrationshare),
      .custom_dma_burst_4_downstream_burstcount                                  (custom_dma_burst_4_downstream_burstcount),
      .custom_dma_burst_4_downstream_byteenable                                  (custom_dma_burst_4_downstream_byteenable),
      .custom_dma_burst_4_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_4_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_latency_counter                             (custom_dma_burst_4_downstream_latency_counter),
      .custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_4_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_read                                        (custom_dma_burst_4_downstream_read),
      .custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_4_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_4_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_4_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_4_downstream_write                                       (custom_dma_burst_4_downstream_write),
      .custom_dma_burst_4_downstream_writedata                                   (custom_dma_burst_4_downstream_writedata),
      .custom_dma_burst_5_downstream_address_to_slave                            (custom_dma_burst_5_downstream_address_to_slave),
      .custom_dma_burst_5_downstream_arbitrationshare                            (custom_dma_burst_5_downstream_arbitrationshare),
      .custom_dma_burst_5_downstream_burstcount                                  (custom_dma_burst_5_downstream_burstcount),
      .custom_dma_burst_5_downstream_byteenable                                  (custom_dma_burst_5_downstream_byteenable),
      .custom_dma_burst_5_downstream_granted_ddr_sdram_s1                        (custom_dma_burst_5_downstream_granted_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_latency_counter                             (custom_dma_burst_5_downstream_latency_counter),
      .custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1              (custom_dma_burst_5_downstream_qualified_request_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_read                                        (custom_dma_burst_5_downstream_read),
      .custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1                (custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register (custom_dma_burst_5_downstream_read_data_valid_ddr_sdram_s1_shift_register),
      .custom_dma_burst_5_downstream_requests_ddr_sdram_s1                       (custom_dma_burst_5_downstream_requests_ddr_sdram_s1),
      .custom_dma_burst_5_downstream_write                                       (custom_dma_burst_5_downstream_write),
      .custom_dma_burst_5_downstream_writedata                                   (custom_dma_burst_5_downstream_writedata),
      .d1_ddr_sdram_s1_end_xfer                                                  (d1_ddr_sdram_s1_end_xfer),
      .ddr_sdram_s1_address                                                      (ddr_sdram_s1_address),
      .ddr_sdram_s1_beginbursttransfer                                           (ddr_sdram_s1_beginbursttransfer),
      .ddr_sdram_s1_burstcount                                                   (ddr_sdram_s1_burstcount),
      .ddr_sdram_s1_byteenable                                                   (ddr_sdram_s1_byteenable),
      .ddr_sdram_s1_read                                                         (ddr_sdram_s1_read),
      .ddr_sdram_s1_readdata                                                     (ddr_sdram_s1_readdata),
      .ddr_sdram_s1_readdata_from_sa                                             (ddr_sdram_s1_readdata_from_sa),
      .ddr_sdram_s1_readdatavalid                                                (ddr_sdram_s1_readdatavalid),
      .ddr_sdram_s1_reset_n                                                      (ddr_sdram_s1_reset_n),
      .ddr_sdram_s1_waitrequest_n                                                (ddr_sdram_s1_waitrequest_n),
      .ddr_sdram_s1_waitrequest_n_from_sa                                        (ddr_sdram_s1_waitrequest_n_from_sa),
      .ddr_sdram_s1_write                                                        (ddr_sdram_s1_write),
      .ddr_sdram_s1_writedata                                                    (ddr_sdram_s1_writedata),
      .reset_n                                                                   (system_clk_reset_n)
    );

  ddr_sdram the_ddr_sdram
    (
      .clk                 (system_clk),
      .clk_to_sdram        (clk_to_sdram_from_the_ddr_sdram),
      .clk_to_sdram_n      (clk_to_sdram_n_from_the_ddr_sdram),
      .ddr_a               (ddr_a_from_the_ddr_sdram),
      .ddr_ba              (ddr_ba_from_the_ddr_sdram),
      .ddr_cas_n           (ddr_cas_n_from_the_ddr_sdram),
      .ddr_cke             (ddr_cke_from_the_ddr_sdram),
      .ddr_cs_n            (ddr_cs_n_from_the_ddr_sdram),
      .ddr_dm              (ddr_dm_from_the_ddr_sdram),
      .ddr_dq              (ddr_dq_to_and_from_the_ddr_sdram),
      .ddr_dqs             (ddr_dqs_to_and_from_the_ddr_sdram),
      .ddr_ras_n           (ddr_ras_n_from_the_ddr_sdram),
      .ddr_we_n            (ddr_we_n_from_the_ddr_sdram),
      .dqs_delay_ctrl      (dqs_delay_ctrl_to_the_ddr_sdram),
      .dqsupdate           (dqsupdate_to_the_ddr_sdram),
      .local_addr          (ddr_sdram_s1_address),
      .local_be            (ddr_sdram_s1_byteenable),
      .local_burstbegin    (ddr_sdram_s1_beginbursttransfer),
      .local_rdata         (ddr_sdram_s1_readdata),
      .local_rdata_valid   (ddr_sdram_s1_readdatavalid),
      .local_read_req      (ddr_sdram_s1_read),
      .local_ready         (ddr_sdram_s1_waitrequest_n),
      .local_size          (ddr_sdram_s1_burstcount),
      .local_wdata         (ddr_sdram_s1_writedata),
      .local_write_req     (ddr_sdram_s1_write),
      .reset_n             (ddr_sdram_s1_reset_n),
      .stratix_dll_control (stratix_dll_control_from_the_ddr_sdram),
      .write_clk           (write_clk_to_the_ddr_sdram)
    );

  ext_ssram_bus_avalon_slave_arbitrator the_ext_ssram_bus_avalon_slave
    (
      .adsc_n_to_the_ext_ssram                                      (adsc_n_to_the_ext_ssram),
      .bw_n_to_the_ext_ssram                                        (bw_n_to_the_ext_ssram),
      .bwe_n_to_the_ext_ssram                                       (bwe_n_to_the_ext_ssram),
      .chipenable1_n_to_the_ext_ssram                               (chipenable1_n_to_the_ext_ssram),
      .clk                                                          (system_clk),
      .custom_dma_burst_0_downstream_address_to_slave               (custom_dma_burst_0_downstream_address_to_slave),
      .custom_dma_burst_0_downstream_arbitrationshare               (custom_dma_burst_0_downstream_arbitrationshare),
      .custom_dma_burst_0_downstream_burstcount                     (custom_dma_burst_0_downstream_burstcount),
      .custom_dma_burst_0_downstream_byteenable                     (custom_dma_burst_0_downstream_byteenable),
      .custom_dma_burst_0_downstream_granted_ext_ssram_s1           (custom_dma_burst_0_downstream_granted_ext_ssram_s1),
      .custom_dma_burst_0_downstream_latency_counter                (custom_dma_burst_0_downstream_latency_counter),
      .custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1 (custom_dma_burst_0_downstream_qualified_request_ext_ssram_s1),
      .custom_dma_burst_0_downstream_read                           (custom_dma_burst_0_downstream_read),
      .custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1   (custom_dma_burst_0_downstream_read_data_valid_ext_ssram_s1),
      .custom_dma_burst_0_downstream_requests_ext_ssram_s1          (custom_dma_burst_0_downstream_requests_ext_ssram_s1),
      .custom_dma_burst_0_downstream_write                          (custom_dma_burst_0_downstream_write),
      .custom_dma_burst_0_downstream_writedata                      (custom_dma_burst_0_downstream_writedata),
      .d1_ext_ssram_bus_avalon_slave_end_xfer                       (d1_ext_ssram_bus_avalon_slave_end_xfer),
      .ext_ssram_bus_address                                        (ext_ssram_bus_address),
      .ext_ssram_bus_data                                           (ext_ssram_bus_data),
      .fir_dma_read_master_address_to_slave                         (fir_dma_read_master_address_to_slave),
      .fir_dma_read_master_granted_ext_ssram_s1                     (fir_dma_read_master_granted_ext_ssram_s1),
      .fir_dma_read_master_latency_counter                          (fir_dma_read_master_latency_counter),
      .fir_dma_read_master_qualified_request_ext_ssram_s1           (fir_dma_read_master_qualified_request_ext_ssram_s1),
      .fir_dma_read_master_read                                     (fir_dma_read_master_read),
      .fir_dma_read_master_read_data_valid_ext_ssram_s1             (fir_dma_read_master_read_data_valid_ext_ssram_s1),
      .fir_dma_read_master_requests_ext_ssram_s1                    (fir_dma_read_master_requests_ext_ssram_s1),
      .incoming_ext_ssram_bus_data                                  (incoming_ext_ssram_bus_data),
      .outputenable_n_to_the_ext_ssram                              (outputenable_n_to_the_ext_ssram),
      .reset_n                                                      (system_clk_reset_n)
    );

  fir_dma_control_arbitrator the_fir_dma_control
    (
      .clk                                                  (system_clk),
      .d1_fir_dma_control_end_xfer                          (d1_fir_dma_control_end_xfer),
      .fir_dma_control_address                              (fir_dma_control_address),
      .fir_dma_control_byteenable                           (fir_dma_control_byteenable),
      .fir_dma_control_irq                                  (fir_dma_control_irq),
      .fir_dma_control_irq_from_sa                          (fir_dma_control_irq_from_sa),
      .fir_dma_control_read                                 (fir_dma_control_read),
      .fir_dma_control_readdata                             (fir_dma_control_readdata),
      .fir_dma_control_readdata_from_sa                     (fir_dma_control_readdata_from_sa),
      .fir_dma_control_reset                                (fir_dma_control_reset),
      .fir_dma_control_write                                (fir_dma_control_write),
      .fir_dma_control_writedata                            (fir_dma_control_writedata),
      .pipeline_bridge_m1_address_to_slave                  (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                        (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                        (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                        (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_fir_dma_control           (pipeline_bridge_m1_granted_fir_dma_control),
      .pipeline_bridge_m1_latency_counter                   (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_fir_dma_control (pipeline_bridge_m1_qualified_request_fir_dma_control),
      .pipeline_bridge_m1_read                              (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_fir_dma_control   (pipeline_bridge_m1_read_data_valid_fir_dma_control),
      .pipeline_bridge_m1_requests_fir_dma_control          (pipeline_bridge_m1_requests_fir_dma_control),
      .pipeline_bridge_m1_write                             (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                         (pipeline_bridge_m1_writedata),
      .reset_n                                              (system_clk_reset_n)
    );

  fir_dma_read_master_arbitrator the_fir_dma_read_master
    (
      .clk                                                (system_clk),
      .d1_ext_ssram_bus_avalon_slave_end_xfer             (d1_ext_ssram_bus_avalon_slave_end_xfer),
      .fir_dma_read_master_address                        (fir_dma_read_master_address),
      .fir_dma_read_master_address_to_slave               (fir_dma_read_master_address_to_slave),
      .fir_dma_read_master_byteenable                     (fir_dma_read_master_byteenable),
      .fir_dma_read_master_granted_ext_ssram_s1           (fir_dma_read_master_granted_ext_ssram_s1),
      .fir_dma_read_master_latency_counter                (fir_dma_read_master_latency_counter),
      .fir_dma_read_master_qualified_request_ext_ssram_s1 (fir_dma_read_master_qualified_request_ext_ssram_s1),
      .fir_dma_read_master_read                           (fir_dma_read_master_read),
      .fir_dma_read_master_read_data_valid_ext_ssram_s1   (fir_dma_read_master_read_data_valid_ext_ssram_s1),
      .fir_dma_read_master_readdata                       (fir_dma_read_master_readdata),
      .fir_dma_read_master_readdatavalid                  (fir_dma_read_master_readdatavalid),
      .fir_dma_read_master_requests_ext_ssram_s1          (fir_dma_read_master_requests_ext_ssram_s1),
      .fir_dma_read_master_waitrequest                    (fir_dma_read_master_waitrequest),
      .incoming_ext_ssram_bus_data                        (incoming_ext_ssram_bus_data),
      .reset_n                                            (system_clk_reset_n)
    );

  fir_dma_write_master_arbitrator the_fir_dma_write_master
    (
      .clk                                                                (system_clk),
      .custom_dma_burst_5_upstream_waitrequest_from_sa                    (custom_dma_burst_5_upstream_waitrequest_from_sa),
      .d1_custom_dma_burst_5_upstream_end_xfer                            (d1_custom_dma_burst_5_upstream_end_xfer),
      .fir_dma_write_master_address                                       (fir_dma_write_master_address),
      .fir_dma_write_master_address_to_slave                              (fir_dma_write_master_address_to_slave),
      .fir_dma_write_master_burstcount                                    (fir_dma_write_master_burstcount),
      .fir_dma_write_master_byteenable                                    (fir_dma_write_master_byteenable),
      .fir_dma_write_master_granted_custom_dma_burst_5_upstream           (fir_dma_write_master_granted_custom_dma_burst_5_upstream),
      .fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream (fir_dma_write_master_qualified_request_custom_dma_burst_5_upstream),
      .fir_dma_write_master_requests_custom_dma_burst_5_upstream          (fir_dma_write_master_requests_custom_dma_burst_5_upstream),
      .fir_dma_write_master_waitrequest                                   (fir_dma_write_master_waitrequest),
      .fir_dma_write_master_write                                         (fir_dma_write_master_write),
      .fir_dma_write_master_writedata                                     (fir_dma_write_master_writedata),
      .reset_n                                                            (system_clk_reset_n)
    );

  fir_dma the_fir_dma
    (
      .clk                       (system_clk),
      .read_master_address       (fir_dma_read_master_address),
      .read_master_byteenable    (fir_dma_read_master_byteenable),
      .read_master_read          (fir_dma_read_master_read),
      .read_master_readdata      (fir_dma_read_master_readdata),
      .read_master_readdatavalid (fir_dma_read_master_readdatavalid),
      .read_master_waitrequest   (fir_dma_read_master_waitrequest),
      .reset                     (fir_dma_control_reset),
      .slave_address             (fir_dma_control_address),
      .slave_byteenable          (fir_dma_control_byteenable),
      .slave_irq                 (fir_dma_control_irq),
      .slave_read                (fir_dma_control_read),
      .slave_readdata            (fir_dma_control_readdata),
      .slave_write               (fir_dma_control_write),
      .slave_writedata           (fir_dma_control_writedata),
      .write_master_address      (fir_dma_write_master_address),
      .write_master_burstcount   (fir_dma_write_master_burstcount),
      .write_master_byteenable   (fir_dma_write_master_byteenable),
      .write_master_waitrequest  (fir_dma_write_master_waitrequest),
      .write_master_write        (fir_dma_write_master_write),
      .write_master_writedata    (fir_dma_write_master_writedata)
    );

  jtag_uart_avalon_jtag_slave_arbitrator the_jtag_uart_avalon_jtag_slave
    (
      .clk                                                              (system_clk),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                          (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .jtag_uart_avalon_jtag_slave_address                              (jtag_uart_avalon_jtag_slave_address),
      .jtag_uart_avalon_jtag_slave_chipselect                           (jtag_uart_avalon_jtag_slave_chipselect),
      .jtag_uart_avalon_jtag_slave_dataavailable                        (jtag_uart_avalon_jtag_slave_dataavailable),
      .jtag_uart_avalon_jtag_slave_dataavailable_from_sa                (jtag_uart_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_avalon_jtag_slave_irq                                  (jtag_uart_avalon_jtag_slave_irq),
      .jtag_uart_avalon_jtag_slave_irq_from_sa                          (jtag_uart_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_avalon_jtag_slave_read_n                               (jtag_uart_avalon_jtag_slave_read_n),
      .jtag_uart_avalon_jtag_slave_readdata                             (jtag_uart_avalon_jtag_slave_readdata),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                     (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readyfordata                         (jtag_uart_avalon_jtag_slave_readyfordata),
      .jtag_uart_avalon_jtag_slave_readyfordata_from_sa                 (jtag_uart_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_avalon_jtag_slave_reset_n                              (jtag_uart_avalon_jtag_slave_reset_n),
      .jtag_uart_avalon_jtag_slave_waitrequest                          (jtag_uart_avalon_jtag_slave_waitrequest),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                  (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_avalon_jtag_slave_write_n                              (jtag_uart_avalon_jtag_slave_write_n),
      .jtag_uart_avalon_jtag_slave_writedata                            (jtag_uart_avalon_jtag_slave_writedata),
      .pipeline_bridge_m1_address_to_slave                              (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                    (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_chipselect                                    (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave           (pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_latency_counter                               (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave (pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_read                                          (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave          (pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_write                                         (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                     (pipeline_bridge_m1_writedata),
      .reset_n                                                          (system_clk_reset_n)
    );

  jtag_uart the_jtag_uart
    (
      .av_address     (jtag_uart_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_avalon_jtag_slave_writedata),
      .clk            (system_clk),
      .dataavailable  (jtag_uart_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_avalon_jtag_slave_reset_n)
    );

  pipeline_bridge_s1_arbitrator the_pipeline_bridge_s1
    (
      .clk                                                                             (system_clk),
      .custom_dma_burst_1_downstream_address_to_slave                                  (custom_dma_burst_1_downstream_address_to_slave),
      .custom_dma_burst_1_downstream_arbitrationshare                                  (custom_dma_burst_1_downstream_arbitrationshare),
      .custom_dma_burst_1_downstream_burstcount                                        (custom_dma_burst_1_downstream_burstcount),
      .custom_dma_burst_1_downstream_byteenable                                        (custom_dma_burst_1_downstream_byteenable),
      .custom_dma_burst_1_downstream_debugaccess                                       (custom_dma_burst_1_downstream_debugaccess),
      .custom_dma_burst_1_downstream_granted_pipeline_bridge_s1                        (custom_dma_burst_1_downstream_granted_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_latency_counter                                   (custom_dma_burst_1_downstream_latency_counter),
      .custom_dma_burst_1_downstream_nativeaddress                                     (custom_dma_burst_1_downstream_nativeaddress),
      .custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1              (custom_dma_burst_1_downstream_qualified_request_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_read                                              (custom_dma_burst_1_downstream_read),
      .custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1                (custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register (custom_dma_burst_1_downstream_read_data_valid_pipeline_bridge_s1_shift_register),
      .custom_dma_burst_1_downstream_requests_pipeline_bridge_s1                       (custom_dma_burst_1_downstream_requests_pipeline_bridge_s1),
      .custom_dma_burst_1_downstream_write                                             (custom_dma_burst_1_downstream_write),
      .custom_dma_burst_1_downstream_writedata                                         (custom_dma_burst_1_downstream_writedata),
      .custom_dma_burst_2_downstream_address_to_slave                                  (custom_dma_burst_2_downstream_address_to_slave),
      .custom_dma_burst_2_downstream_arbitrationshare                                  (custom_dma_burst_2_downstream_arbitrationshare),
      .custom_dma_burst_2_downstream_burstcount                                        (custom_dma_burst_2_downstream_burstcount),
      .custom_dma_burst_2_downstream_byteenable                                        (custom_dma_burst_2_downstream_byteenable),
      .custom_dma_burst_2_downstream_debugaccess                                       (custom_dma_burst_2_downstream_debugaccess),
      .custom_dma_burst_2_downstream_granted_pipeline_bridge_s1                        (custom_dma_burst_2_downstream_granted_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_latency_counter                                   (custom_dma_burst_2_downstream_latency_counter),
      .custom_dma_burst_2_downstream_nativeaddress                                     (custom_dma_burst_2_downstream_nativeaddress),
      .custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1              (custom_dma_burst_2_downstream_qualified_request_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_read                                              (custom_dma_burst_2_downstream_read),
      .custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1                (custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register (custom_dma_burst_2_downstream_read_data_valid_pipeline_bridge_s1_shift_register),
      .custom_dma_burst_2_downstream_requests_pipeline_bridge_s1                       (custom_dma_burst_2_downstream_requests_pipeline_bridge_s1),
      .custom_dma_burst_2_downstream_write                                             (custom_dma_burst_2_downstream_write),
      .custom_dma_burst_2_downstream_writedata                                         (custom_dma_burst_2_downstream_writedata),
      .d1_pipeline_bridge_s1_end_xfer                                                  (d1_pipeline_bridge_s1_end_xfer),
      .pipeline_bridge_s1_address                                                      (pipeline_bridge_s1_address),
      .pipeline_bridge_s1_arbiterlock                                                  (pipeline_bridge_s1_arbiterlock),
      .pipeline_bridge_s1_arbiterlock2                                                 (pipeline_bridge_s1_arbiterlock2),
      .pipeline_bridge_s1_burstcount                                                   (pipeline_bridge_s1_burstcount),
      .pipeline_bridge_s1_byteenable                                                   (pipeline_bridge_s1_byteenable),
      .pipeline_bridge_s1_chipselect                                                   (pipeline_bridge_s1_chipselect),
      .pipeline_bridge_s1_debugaccess                                                  (pipeline_bridge_s1_debugaccess),
      .pipeline_bridge_s1_endofpacket                                                  (pipeline_bridge_s1_endofpacket),
      .pipeline_bridge_s1_endofpacket_from_sa                                          (pipeline_bridge_s1_endofpacket_from_sa),
      .pipeline_bridge_s1_nativeaddress                                                (pipeline_bridge_s1_nativeaddress),
      .pipeline_bridge_s1_read                                                         (pipeline_bridge_s1_read),
      .pipeline_bridge_s1_readdata                                                     (pipeline_bridge_s1_readdata),
      .pipeline_bridge_s1_readdata_from_sa                                             (pipeline_bridge_s1_readdata_from_sa),
      .pipeline_bridge_s1_readdatavalid                                                (pipeline_bridge_s1_readdatavalid),
      .pipeline_bridge_s1_reset_n                                                      (pipeline_bridge_s1_reset_n),
      .pipeline_bridge_s1_waitrequest                                                  (pipeline_bridge_s1_waitrequest),
      .pipeline_bridge_s1_waitrequest_from_sa                                          (pipeline_bridge_s1_waitrequest_from_sa),
      .pipeline_bridge_s1_write                                                        (pipeline_bridge_s1_write),
      .pipeline_bridge_s1_writedata                                                    (pipeline_bridge_s1_writedata),
      .reset_n                                                                         (system_clk_reset_n)
    );

  pipeline_bridge_m1_arbitrator the_pipeline_bridge_m1
    (
      .clk                                                              (system_clk),
      .cpu_jtag_debug_module_readdata_from_sa                           (cpu_jtag_debug_module_readdata_from_sa),
      .custom_dma_clock_0_in_endofpacket_from_sa                        (custom_dma_clock_0_in_endofpacket_from_sa),
      .custom_dma_clock_0_in_readdata_from_sa                           (custom_dma_clock_0_in_readdata_from_sa),
      .custom_dma_clock_0_in_waitrequest_from_sa                        (custom_dma_clock_0_in_waitrequest_from_sa),
      .d1_cpu_jtag_debug_module_end_xfer                                (d1_cpu_jtag_debug_module_end_xfer),
      .d1_custom_dma_clock_0_in_end_xfer                                (d1_custom_dma_clock_0_in_end_xfer),
      .d1_fir_dma_control_end_xfer                                      (d1_fir_dma_control_end_xfer),
      .d1_jtag_uart_avalon_jtag_slave_end_xfer                          (d1_jtag_uart_avalon_jtag_slave_end_xfer),
      .d1_sysid_control_slave_end_xfer                                  (d1_sysid_control_slave_end_xfer),
      .d1_timestamp_timer_s1_end_xfer                                   (d1_timestamp_timer_s1_end_xfer),
      .fir_dma_control_readdata_from_sa                                 (fir_dma_control_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_readdata_from_sa                     (jtag_uart_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_avalon_jtag_slave_waitrequest_from_sa                  (jtag_uart_avalon_jtag_slave_waitrequest_from_sa),
      .pipeline_bridge_m1_address                                       (pipeline_bridge_m1_address),
      .pipeline_bridge_m1_address_to_slave                              (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                                    (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_byteenable                                    (pipeline_bridge_m1_byteenable),
      .pipeline_bridge_m1_chipselect                                    (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_endofpacket                                   (pipeline_bridge_m1_endofpacket),
      .pipeline_bridge_m1_granted_cpu_jtag_debug_module                 (pipeline_bridge_m1_granted_cpu_jtag_debug_module),
      .pipeline_bridge_m1_granted_custom_dma_clock_0_in                 (pipeline_bridge_m1_granted_custom_dma_clock_0_in),
      .pipeline_bridge_m1_granted_fir_dma_control                       (pipeline_bridge_m1_granted_fir_dma_control),
      .pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave           (pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_granted_sysid_control_slave                   (pipeline_bridge_m1_granted_sysid_control_slave),
      .pipeline_bridge_m1_granted_timestamp_timer_s1                    (pipeline_bridge_m1_granted_timestamp_timer_s1),
      .pipeline_bridge_m1_latency_counter                               (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module       (pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module),
      .pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in       (pipeline_bridge_m1_qualified_request_custom_dma_clock_0_in),
      .pipeline_bridge_m1_qualified_request_fir_dma_control             (pipeline_bridge_m1_qualified_request_fir_dma_control),
      .pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave (pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_qualified_request_sysid_control_slave         (pipeline_bridge_m1_qualified_request_sysid_control_slave),
      .pipeline_bridge_m1_qualified_request_timestamp_timer_s1          (pipeline_bridge_m1_qualified_request_timestamp_timer_s1),
      .pipeline_bridge_m1_read                                          (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module         (pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module),
      .pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in         (pipeline_bridge_m1_read_data_valid_custom_dma_clock_0_in),
      .pipeline_bridge_m1_read_data_valid_fir_dma_control               (pipeline_bridge_m1_read_data_valid_fir_dma_control),
      .pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave   (pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_read_data_valid_sysid_control_slave           (pipeline_bridge_m1_read_data_valid_sysid_control_slave),
      .pipeline_bridge_m1_read_data_valid_timestamp_timer_s1            (pipeline_bridge_m1_read_data_valid_timestamp_timer_s1),
      .pipeline_bridge_m1_readdata                                      (pipeline_bridge_m1_readdata),
      .pipeline_bridge_m1_readdatavalid                                 (pipeline_bridge_m1_readdatavalid),
      .pipeline_bridge_m1_requests_cpu_jtag_debug_module                (pipeline_bridge_m1_requests_cpu_jtag_debug_module),
      .pipeline_bridge_m1_requests_custom_dma_clock_0_in                (pipeline_bridge_m1_requests_custom_dma_clock_0_in),
      .pipeline_bridge_m1_requests_fir_dma_control                      (pipeline_bridge_m1_requests_fir_dma_control),
      .pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave          (pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave),
      .pipeline_bridge_m1_requests_sysid_control_slave                  (pipeline_bridge_m1_requests_sysid_control_slave),
      .pipeline_bridge_m1_requests_timestamp_timer_s1                   (pipeline_bridge_m1_requests_timestamp_timer_s1),
      .pipeline_bridge_m1_waitrequest                                   (pipeline_bridge_m1_waitrequest),
      .pipeline_bridge_m1_write                                         (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                                     (pipeline_bridge_m1_writedata),
      .reset_n                                                          (system_clk_reset_n),
      .sysid_control_slave_readdata_from_sa                             (sysid_control_slave_readdata_from_sa),
      .timestamp_timer_s1_readdata_from_sa                              (timestamp_timer_s1_readdata_from_sa)
    );

  pipeline_bridge the_pipeline_bridge
    (
      .clk              (system_clk),
      .m1_address       (pipeline_bridge_m1_address),
      .m1_burstcount    (pipeline_bridge_m1_burstcount),
      .m1_byteenable    (pipeline_bridge_m1_byteenable),
      .m1_chipselect    (pipeline_bridge_m1_chipselect),
      .m1_debugaccess   (pipeline_bridge_m1_debugaccess),
      .m1_endofpacket   (pipeline_bridge_m1_endofpacket),
      .m1_read          (pipeline_bridge_m1_read),
      .m1_readdata      (pipeline_bridge_m1_readdata),
      .m1_readdatavalid (pipeline_bridge_m1_readdatavalid),
      .m1_waitrequest   (pipeline_bridge_m1_waitrequest),
      .m1_write         (pipeline_bridge_m1_write),
      .m1_writedata     (pipeline_bridge_m1_writedata),
      .reset_n          (pipeline_bridge_s1_reset_n),
      .s1_address       (pipeline_bridge_s1_address),
      .s1_arbiterlock   (pipeline_bridge_s1_arbiterlock),
      .s1_arbiterlock2  (pipeline_bridge_s1_arbiterlock2),
      .s1_burstcount    (pipeline_bridge_s1_burstcount),
      .s1_byteenable    (pipeline_bridge_s1_byteenable),
      .s1_chipselect    (pipeline_bridge_s1_chipselect),
      .s1_debugaccess   (pipeline_bridge_s1_debugaccess),
      .s1_endofpacket   (pipeline_bridge_s1_endofpacket),
      .s1_nativeaddress (pipeline_bridge_s1_nativeaddress),
      .s1_read          (pipeline_bridge_s1_read),
      .s1_readdata      (pipeline_bridge_s1_readdata),
      .s1_readdatavalid (pipeline_bridge_s1_readdatavalid),
      .s1_waitrequest   (pipeline_bridge_s1_waitrequest),
      .s1_write         (pipeline_bridge_s1_write),
      .s1_writedata     (pipeline_bridge_s1_writedata)
    );

  pll_s1_arbitrator the_pll_s1
    (
      .clk                                             (external_clk),
      .custom_dma_clock_0_out_address_to_slave         (custom_dma_clock_0_out_address_to_slave),
      .custom_dma_clock_0_out_granted_pll_s1           (custom_dma_clock_0_out_granted_pll_s1),
      .custom_dma_clock_0_out_nativeaddress            (custom_dma_clock_0_out_nativeaddress),
      .custom_dma_clock_0_out_qualified_request_pll_s1 (custom_dma_clock_0_out_qualified_request_pll_s1),
      .custom_dma_clock_0_out_read                     (custom_dma_clock_0_out_read),
      .custom_dma_clock_0_out_read_data_valid_pll_s1   (custom_dma_clock_0_out_read_data_valid_pll_s1),
      .custom_dma_clock_0_out_requests_pll_s1          (custom_dma_clock_0_out_requests_pll_s1),
      .custom_dma_clock_0_out_write                    (custom_dma_clock_0_out_write),
      .custom_dma_clock_0_out_writedata                (custom_dma_clock_0_out_writedata),
      .d1_pll_s1_end_xfer                              (d1_pll_s1_end_xfer),
      .pll_s1_address                                  (pll_s1_address),
      .pll_s1_chipselect                               (pll_s1_chipselect),
      .pll_s1_read                                     (pll_s1_read),
      .pll_s1_readdata                                 (pll_s1_readdata),
      .pll_s1_readdata_from_sa                         (pll_s1_readdata_from_sa),
      .pll_s1_reset_n                                  (pll_s1_reset_n),
      .pll_s1_resetrequest                             (pll_s1_resetrequest),
      .pll_s1_resetrequest_from_sa                     (pll_s1_resetrequest_from_sa),
      .pll_s1_write                                    (pll_s1_write),
      .pll_s1_writedata                                (pll_s1_writedata),
      .reset_n                                         (external_clk_reset_n)
    );

  //system_clk out_clk assignment, which is an e_assign
  assign system_clk = out_clk_pll_c0;

  //ssram_clk out_clk assignment, which is an e_assign
  assign ssram_clk = out_clk_pll_c1;

  //sdram_write_clk out_clk assignment, which is an e_assign
  assign sdram_write_clk = out_clk_pll_c2;

  pll the_pll
    (
      .address      (pll_s1_address),
      .c0           (out_clk_pll_c0),
      .c1           (out_clk_pll_c1),
      .c2           (out_clk_pll_c2),
      .chipselect   (pll_s1_chipselect),
      .clk          (external_clk),
      .read         (pll_s1_read),
      .readdata     (pll_s1_readdata),
      .reset_n      (pll_s1_reset_n),
      .resetrequest (pll_s1_resetrequest),
      .write        (pll_s1_write),
      .writedata    (pll_s1_writedata)
    );

  sysid_control_slave_arbitrator the_sysid_control_slave
    (
      .clk                                                      (system_clk),
      .d1_sysid_control_slave_end_xfer                          (d1_sysid_control_slave_end_xfer),
      .pipeline_bridge_m1_address_to_slave                      (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                            (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_chipselect                            (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_sysid_control_slave           (pipeline_bridge_m1_granted_sysid_control_slave),
      .pipeline_bridge_m1_latency_counter                       (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_sysid_control_slave (pipeline_bridge_m1_qualified_request_sysid_control_slave),
      .pipeline_bridge_m1_read                                  (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_sysid_control_slave   (pipeline_bridge_m1_read_data_valid_sysid_control_slave),
      .pipeline_bridge_m1_requests_sysid_control_slave          (pipeline_bridge_m1_requests_sysid_control_slave),
      .pipeline_bridge_m1_write                                 (pipeline_bridge_m1_write),
      .reset_n                                                  (system_clk_reset_n),
      .sysid_control_slave_address                              (sysid_control_slave_address),
      .sysid_control_slave_readdata                             (sysid_control_slave_readdata),
      .sysid_control_slave_readdata_from_sa                     (sysid_control_slave_readdata_from_sa)
    );

  sysid the_sysid
    (
      .address  (sysid_control_slave_address),
      .readdata (sysid_control_slave_readdata)
    );

  timestamp_timer_s1_arbitrator the_timestamp_timer_s1
    (
      .clk                                                     (system_clk),
      .d1_timestamp_timer_s1_end_xfer                          (d1_timestamp_timer_s1_end_xfer),
      .pipeline_bridge_m1_address_to_slave                     (pipeline_bridge_m1_address_to_slave),
      .pipeline_bridge_m1_burstcount                           (pipeline_bridge_m1_burstcount),
      .pipeline_bridge_m1_chipselect                           (pipeline_bridge_m1_chipselect),
      .pipeline_bridge_m1_granted_timestamp_timer_s1           (pipeline_bridge_m1_granted_timestamp_timer_s1),
      .pipeline_bridge_m1_latency_counter                      (pipeline_bridge_m1_latency_counter),
      .pipeline_bridge_m1_qualified_request_timestamp_timer_s1 (pipeline_bridge_m1_qualified_request_timestamp_timer_s1),
      .pipeline_bridge_m1_read                                 (pipeline_bridge_m1_read),
      .pipeline_bridge_m1_read_data_valid_timestamp_timer_s1   (pipeline_bridge_m1_read_data_valid_timestamp_timer_s1),
      .pipeline_bridge_m1_requests_timestamp_timer_s1          (pipeline_bridge_m1_requests_timestamp_timer_s1),
      .pipeline_bridge_m1_write                                (pipeline_bridge_m1_write),
      .pipeline_bridge_m1_writedata                            (pipeline_bridge_m1_writedata),
      .reset_n                                                 (system_clk_reset_n),
      .timestamp_timer_s1_address                              (timestamp_timer_s1_address),
      .timestamp_timer_s1_chipselect                           (timestamp_timer_s1_chipselect),
      .timestamp_timer_s1_irq                                  (timestamp_timer_s1_irq),
      .timestamp_timer_s1_irq_from_sa                          (timestamp_timer_s1_irq_from_sa),
      .timestamp_timer_s1_readdata                             (timestamp_timer_s1_readdata),
      .timestamp_timer_s1_readdata_from_sa                     (timestamp_timer_s1_readdata_from_sa),
      .timestamp_timer_s1_reset_n                              (timestamp_timer_s1_reset_n),
      .timestamp_timer_s1_write_n                              (timestamp_timer_s1_write_n),
      .timestamp_timer_s1_writedata                            (timestamp_timer_s1_writedata)
    );

  timestamp_timer the_timestamp_timer
    (
      .address    (timestamp_timer_s1_address),
      .chipselect (timestamp_timer_s1_chipselect),
      .clk        (system_clk),
      .irq        (timestamp_timer_s1_irq),
      .readdata   (timestamp_timer_s1_readdata),
      .reset_n    (timestamp_timer_s1_reset_n),
      .write_n    (timestamp_timer_s1_write_n),
      .writedata  (timestamp_timer_s1_writedata)
    );

  //reset is asserted asynchronously and deasserted synchronously
  custom_dma_reset_system_clk_domain_synch_module custom_dma_reset_system_clk_domain_synch
    (
      .clk      (system_clk),
      .data_in  (1'b1),
      .data_out (system_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    cpu_jtag_debug_module_resetrequest_from_sa |
    cpu_jtag_debug_module_resetrequest_from_sa |
    0 |
    pll_s1_resetrequest_from_sa |
    pll_s1_resetrequest_from_sa);

  //reset is asserted asynchronously and deasserted synchronously
  custom_dma_reset_external_clk_domain_synch_module custom_dma_reset_external_clk_domain_synch
    (
      .clk      (external_clk),
      .data_in  (1'b1),
      .data_out (external_clk_reset_n),
      .reset_n  (reset_n_sources)
    );

  //custom_dma_burst_1_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign custom_dma_burst_1_upstream_writedata = 0;

  //custom_dma_burst_3_upstream_writedata of type writedata does not connect to anything so wire it to default (0)
  assign custom_dma_burst_3_upstream_writedata = 0;

  //custom_dma_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  assign custom_dma_clock_0_out_endofpacket = 0;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_lane0_module (
                                // inputs:
                                 clk,
                                 data,
                                 rdaddress,
                                 rdclken,
                                 reset_n,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 18: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 18: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 18: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [524287: 0];
  wire    [  7: 0] q;
  reg     [ 18: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ssram_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ssram_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 19,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_lane1_module (
                                // inputs:
                                 clk,
                                 data,
                                 rdaddress,
                                 rdclken,
                                 reset_n,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 18: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 18: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 18: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [524287: 0];
  wire    [  7: 0] q;
  reg     [ 18: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ssram_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ssram_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 19,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_lane2_module (
                                // inputs:
                                 clk,
                                 data,
                                 rdaddress,
                                 rdclken,
                                 reset_n,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 18: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 18: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 18: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [524287: 0];
  wire    [  7: 0] q;
  reg     [ 18: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ssram_lane2.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ssram_lane2.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 19,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram_lane3_module (
                                // inputs:
                                 clk,
                                 data,
                                 rdaddress,
                                 rdclken,
                                 reset_n,
                                 wraddress,
                                 wrclock,
                                 wren,

                                // outputs:
                                 q
                              )
;

  output  [  7: 0] q;
  input            clk;
  input   [  7: 0] data;
  input   [ 18: 0] rdaddress;
  input            rdclken;
  input            reset_n;
  input   [ 18: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 18: 0] d1_rdaddress;
  reg     [  7: 0] mem_array [524287: 0];
  wire    [  7: 0] q;
  reg     [ 18: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_rdaddress <= 0;
          read_address <= 0;
        end
      else if (rdclken)
        begin
          d1_rdaddress <= rdaddress;
          read_address <= d1_rdaddress;
        end
    end


  // Data read is synchronized through latent_rdaddress.
  assign q = mem_array[read_address];

initial
    $readmemh("ext_ssram_lane3.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .rdclock (clk),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "ext_ssram_lane3.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "REGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "REGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 19,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ext_ssram (
                   // inputs:
                    address,
                    adsc_n,
                    bw_n,
                    bwe_n,
                    chipenable1_n,
                    clk,
                    outputenable_n,
                    reset_n,

                   // outputs:
                    data
                 )
;

  inout   [ 31: 0] data;
  input   [ 18: 0] address;
  input            adsc_n;
  input   [  3: 0] bw_n;
  input            bwe_n;
  input            chipenable1_n;
  input            clk;
  input            outputenable_n;
  input            reset_n;

  wire    [ 31: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [  7: 0] data_2;
  wire    [  7: 0] data_3;
  wire    [ 31: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  wire    [  7: 0] q_2;
  wire    [  7: 0] q_3;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //ext_ssram_lane0, which is an e_ram
  ext_ssram_lane0_module ext_ssram_lane0
    (
      .clk       (clk),
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[0])
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //ext_ssram_lane1, which is an e_ram
  ext_ssram_lane1_module ext_ssram_lane1
    (
      .clk       (clk),
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[1])
    );

  assign data_2 = logic_vector_gasket[23 : 16];
  //ext_ssram_lane2, which is an e_ram
  ext_ssram_lane2_module ext_ssram_lane2
    (
      .clk       (clk),
      .data      (data_2),
      .q         (q_2),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[2])
    );

  assign data_3 = logic_vector_gasket[31 : 24];
  //ext_ssram_lane3, which is an e_ram
  ext_ssram_lane3_module ext_ssram_lane3
    (
      .clk       (clk),
      .data      (data_3),
      .q         (q_3),
      .rdaddress (address),
      .rdclken   (1'b1),
      .reset_n   (reset_n),
      .wraddress (address),
      .wrclock   (clk),
      .wren      (~chipenable1_n & ~bwe_n & ~bw_n[3])
    );

  assign data = (~chipenable1_n & ~outputenable_n)? {q_3,
    q_2,
    q_1,
    q_0}: {32{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

/* SLline 1 "ddr_sdram_auk_ddr_dqs_group.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ps / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//------------------------------------------------------------------------------
//Parameters:
//Device Family                      : Stratix II
//DQ_PER_DQS                         : 8
//NON-DQS MODE                       : false
//use Resynch clock                  : true
//Resynch clock edge                 : rising
//Postamble Clock Edge               : rising
//Postamble Clock Cycle              : 1
//Intermediate Resynch               : false
//Intermediate Postamble             : false
//Pipeline read Data                 : false
//Enable Postamble Logic             : true
//Postamble Regs Per DQS             : 1
//Stratix Insert DQS delay buffers   : 0
//------------------------------------------------------------------------------
module ddr_sdram_auk_ddr_dqs_group (
                                     // inputs:
                                      capture_clk,
                                      clk,
                                      control_be,
                                      control_doing_rd,
                                      control_doing_wr,
                                      control_dqs_burst,
                                      control_wdata,
                                      control_wdata_valid,
                                      dqs_delay_ctrl,
                                      dqsupdate,
                                      postamble_clk,
                                      reset_n,
                                      resynch_clk,
                                      write_clk,

                                     // outputs:
                                      control_rdata,
                                      ddr_dm,
                                      ddr_dq,
                                      ddr_dqs
                                   )
  /* synthesis ALTERA_ATTRIBUTE = "MESSAGE_DISABLE=14130;SUPPRESS_DA_RULE_INTERNAL=C101;SUPPRESS_DA_RULE_INTERNAL=C103;SUPPRESS_DA_RULE_INTERNAL=C105;SUPPRESS_DA_RULE_INTERNAL=C106;SUPPRESS_DA_RULE_INTERNAL=R104;SUPPRESS_DA_RULE_INTERNAL=A102;SUPPRESS_DA_RULE_INTERNAL=A103;SUPPRESS_DA_RULE_INTERNAL=C104;SUPPRESS_DA_RULE_INTERNAL=D101;SUPPRESS_DA_RULE_INTERNAL=D102;SUPPRESS_DA_RULE_INTERNAL=D103;SUPPRESS_DA_RULE_INTERNAL=R102;SUPPRESS_DA_RULE_INTERNAL=R105" */ ;

  parameter gDLL_INPUT_FREQUENCY = "10000ps";
  parameter gSTRATIXII_DQS_OUT_MODE = "delay_chain2";
  parameter gSTRATIXII_DQS_PHASE = 6000;
  parameter gSTRATIXII_DLL_DELAY_BUFFER_MODE = "low";


  output  [ 15: 0] control_rdata;
  output           ddr_dm;
  inout   [  7: 0] ddr_dq;
  inout            ddr_dqs;
  input            capture_clk;
  input            clk;
  input   [  1: 0] control_be;
  input            control_doing_rd;
  input            control_doing_wr;
  input            control_dqs_burst;
  input   [ 15: 0] control_wdata;
  input            control_wdata_valid;
  input   [  5: 0] dqs_delay_ctrl;
  input            dqsupdate;
  input            postamble_clk;
  input            reset_n;
  input            resynch_clk;
  input            write_clk;

  wire             ZERO;
  wire    [  7: 0] ZEROS;
  wire    [ 13: 0] ZEROS_14;
  wire    [  1: 0] be;
  wire    [ 15: 0] control_rdata;
  wire             ddr_dm;
  wire    [  7: 0] ddr_dq;
  wire             ddr_dqs;
  wire    [ 15: 0] delayed_dq_captured;
  reg     [  1: 0] dm_out;
  wire             doing_rd;
  reg              doing_rd_delayed;
  reg     [  2: 0] doing_rd_pipe;
  wire             doing_wr;
  reg              doing_wr_r;
  wire             dq_capture_clk;
  wire    [ 15: 0] dq_captured_0;
  wire    [  7: 0] dq_captured_falling;
  wire    [  7: 0] dq_captured_rising;
  reg     [  0: 0] dq_enable_reset;
  reg              dq_oe;
  wire             dqs_burst;
  wire    [  0: 0] dqs_clk;
  wire             dqs_oe;
  reg     [  0: 0] dqs_oe_r;
  wire    [ 15: 0] inter_rdata;
  wire    [  0: 0] not_dqs_clk;
  wire    [ 15: 0] rdata;
  wire             reset;
  reg     [ 15: 0] resynched_data;
  wire             tmp_dmout0;
  wire             tmp_dmout1;
  wire    [  0: 0] undelayed_dqs;
  wire    [ 15: 0] wdata;
  reg     [ 15: 0] wdata_r;
  wire             wdata_valid;
  //


  assign ZERO = 1'b0;
  assign ZEROS = 0;
  assign ZEROS_14 = 0;
  assign reset = ~reset_n;
  assign not_dqs_clk = ~dqs_clk;
  // rename user i/f signals, outputs
  assign control_rdata = rdata;

  // rename user i/f signals, inputs
  assign wdata = control_wdata;

  assign wdata_valid = control_wdata_valid;
  assign doing_wr = control_doing_wr;
  assign doing_rd = control_doing_rd;
  assign be = control_be;
  assign dqs_burst = control_dqs_burst;
  //-----------------------------------------------------------------------------
  //DQS pin and its logic
  //Generate the output enable for DQS from the signal that indicates we're
  //doing a write. The DQS burst signal is generated by the controller to keep
  //the DQS toggling for the required burst length.
  //-----------------------------------------------------------------------------

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          dqs_oe_r <= 1'b0;
          doing_wr_r <= 1'b0;
        end
      else 
        begin
          dqs_oe_r <= dqs_oe;
          doing_wr_r <= doing_wr;
        end
    end


  assign dqs_oe = doing_wr | dqs_burst;
  //-----------------------------------------------------------------------------
  //DM pins and their logic
  //Although these don't get tristated like DQ, they do share the same IO timing.
  //-----------------------------------------------------------------------------
  assign tmp_dmout0 = dm_out[0];
  assign tmp_dmout1 = dm_out[1];
  altddio_out dm_pin
    (
      .aclr (reset),
      .aset (),
      .datain_h (tmp_dmout0),
      .datain_l (tmp_dmout1),
      .dataout (ddr_dm),
      .oe (1'b1),
      .outclock (write_clk),
      .outclocken (1'b1)
    );

  defparam dm_pin.extend_oe_disable = "UNUSED",
           dm_pin.intended_device_family = "Stratix II",
           dm_pin.invert_output = "OFF",
           dm_pin.lpm_hint = "UNUSED",
           dm_pin.lpm_type = "altddio_out",
           dm_pin.oe_reg = "UNUSED",
           dm_pin.power_up_high = "OFF",
           dm_pin.width = 1;

  //-----------------------------------------------------------------------------
  //Data mask registers
  //These are the last registers before the registers in the altddio_out. They
  //are clocked off the system clock but feed registers which are clocked off the
  //write clock, so their output is the beginning of 3/4 cycle path.
  //-----------------------------------------------------------------------------
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dm_out <= {2{1'b1}};
      else if (doing_wr)
          // don't latch in data unless it's valid
          dm_out <= ~be;

      else 
        dm_out <= {2{1'b1}};
    end


  //-----------------------------------------------------------------------------
  //Logic to disable the capture registers (particularly during DQS postamble)
  //The output of the dq_enable_reset register holds the dq_enable register in
  //reset (which *enables* the dq capture registers). The controller releases
  //the dq_enable register so that it is clocked by the last falling edge of the
  //read dqs signal. This disables the dq capture registers during and after the
  //dqs postamble so that the output of the dq capture registers can be safely
  //resynchronised.
  //Postamble Clock Cycle  : 1
  //Postamble Clock Edge   : rising
  //Postamble Regs Per DQS : 1
  //-----------------------------------------------------------------------------

  //Use a rising edge for postamble
  //The registers which generate the reset signal to the above registers
  //Can be clocked off the resynch or system clock
  always @(posedge postamble_clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dq_enable_reset <= 1'b0;
      else 
        dq_enable_reset <= doing_rd_delayed;
    end


  //pipeline the doing_rd signal to enable and disable the DQ capture regs at the right time
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          doing_rd_pipe <= 0;
      else 
        //shift bits up
        doing_rd_pipe <= {doing_rd_pipe[1 : 0], doing_rd};

    end


  //It's safe to clock from falling edge of clk to postamble_clk, so use falling edge clock
  always @(negedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          doing_rd_delayed <= 1'b0;
      else 
        doing_rd_delayed <= doing_rd_pipe[1];
    end


  //-----------------------------------------------------------------------------
  //Decide which clock to use for capturing the DQ data
  //-----------------------------------------------------------------------------
  //Use DQS to capture DQ read data
  assign dq_capture_clk = ~dqs_clk;

  //-----------------------------------------------------------------------------
  //DQ pins and their logic
  //-----------------------------------------------------------------------------
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dq_oe <= 1'b0;
      else 
        dq_oe <= doing_wr;
    end


  stratixii_io ^^^$_g_dq_io:0:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[0]),
      .ddiodatain (wdata_r[8]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[0]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[0]),
      .regout (dq_captured_falling[0]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:0:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:0:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:0:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:0:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:0:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:0:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:0:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:0:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:0:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:0:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:0:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:0:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:0:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:0:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:0:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:0:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:0:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:0:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:0:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:0:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:1:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[1]),
      .ddiodatain (wdata_r[9]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[1]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[1]),
      .regout (dq_captured_falling[1]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:1:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:1:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:1:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:1:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:1:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:1:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:1:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:1:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:1:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:1:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:1:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:1:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:1:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:1:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:1:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:1:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:1:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:1:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:1:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:1:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:2:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[2]),
      .ddiodatain (wdata_r[10]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[2]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[2]),
      .regout (dq_captured_falling[2]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:2:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:2:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:2:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:2:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:2:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:2:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:2:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:2:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:2:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:2:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:2:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:2:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:2:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:2:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:2:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:2:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:2:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:2:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:2:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:2:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:3:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[3]),
      .ddiodatain (wdata_r[11]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[3]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[3]),
      .regout (dq_captured_falling[3]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:3:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:3:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:3:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:3:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:3:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:3:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:3:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:3:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:3:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:3:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:3:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:3:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:3:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:3:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:3:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:3:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:3:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:3:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:3:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:3:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:4:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[4]),
      .ddiodatain (wdata_r[12]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[4]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[4]),
      .regout (dq_captured_falling[4]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:4:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:4:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:4:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:4:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:4:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:4:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:4:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:4:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:4:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:4:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:4:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:4:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:4:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:4:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:4:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:4:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:4:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:4:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:4:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:4:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:5:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[5]),
      .ddiodatain (wdata_r[13]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[5]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[5]),
      .regout (dq_captured_falling[5]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:5:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:5:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:5:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:5:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:5:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:5:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:5:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:5:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:5:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:5:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:5:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:5:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:5:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:5:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:5:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:5:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:5:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:5:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:5:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:5:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:6:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[6]),
      .ddiodatain (wdata_r[14]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[6]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[6]),
      .regout (dq_captured_falling[6]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:6:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:6:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:6:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:6:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:6:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:6:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:6:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:6:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:6:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:6:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:6:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:6:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:6:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:6:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:6:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:6:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:6:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:6:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:6:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:6:dq_io_$^^^.tie_off_output_clock_enable = "false";

  stratixii_io ^^^$_g_dq_io:7:dq_io_$^^^
    (
      .areset (reset),
      .combout (),
      .datain (wdata_r[7]),
      .ddiodatain (wdata_r[15]),
      .ddioinclk (ZEROS[0]),
      .ddioregout (dq_captured_rising[7]),
      .delayctrlin (),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (),
      .dqsupdateen (),
      .inclk (dq_capture_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dq_oe),
      .offsetctrlin (),
      .outclk (write_clk),
      .outclkena (1'b1),
      .padio (ddr_dq[7]),
      .regout (dq_captured_falling[7]),
      .sreset (),
      .terminationcontrol ()
    );

  defparam ^^^$_g_dq_io:7:dq_io_$^^^.bus_hold = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.ddio_mode = "bidir",
           ^^^$_g_dq_io:7:dq_io_$^^^.ddioinclk_input = "negated_inclk",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_ctrl_latches_enable = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_delay_buffer_mode = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_edge_detect_enable = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_input_frequency = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_offsetctrl_enable = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_out_mode = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.dqs_phase_shift = 0,
           ^^^$_g_dq_io:7:dq_io_$^^^.extend_oe_disable = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.gated_dqs = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.inclk_input = "dqs_bus",
           ^^^$_g_dq_io:7:dq_io_$^^^.input_async_reset = "clear",
           ^^^$_g_dq_io:7:dq_io_$^^^.input_power_up = "low",
           ^^^$_g_dq_io:7:dq_io_$^^^.input_register_mode = "register",
           ^^^$_g_dq_io:7:dq_io_$^^^.input_sync_reset = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.lpm_type = "stratixii_io",
           ^^^$_g_dq_io:7:dq_io_$^^^.oe_async_reset = "clear",
           ^^^$_g_dq_io:7:dq_io_$^^^.oe_power_up = "low",
           ^^^$_g_dq_io:7:dq_io_$^^^.oe_register_mode = "register",
           ^^^$_g_dq_io:7:dq_io_$^^^.oe_sync_reset = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.open_drain_output = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.operation_mode = "bidir",
           ^^^$_g_dq_io:7:dq_io_$^^^.output_async_reset = "clear",
           ^^^$_g_dq_io:7:dq_io_$^^^.output_power_up = "low",
           ^^^$_g_dq_io:7:dq_io_$^^^.output_register_mode = "register",
           ^^^$_g_dq_io:7:dq_io_$^^^.output_sync_reset = "none",
           ^^^$_g_dq_io:7:dq_io_$^^^.sim_dqs_delay_increment = 0,
           ^^^$_g_dq_io:7:dq_io_$^^^.sim_dqs_intrinsic_delay = 0,
           ^^^$_g_dq_io:7:dq_io_$^^^.sim_dqs_offset_increment = 0,
           ^^^$_g_dq_io:7:dq_io_$^^^.tie_off_oe_clock_enable = "false",
           ^^^$_g_dq_io:7:dq_io_$^^^.tie_off_output_clock_enable = "false";

  //-----------------------------------------------------------------------------
  //Write data registers
  //These are the last registers before the registers in the altddio_bidir. They
  //are clocked off the system clock but feed registers which are clocked off the
  //write clock, so their output is the beginning of 3/4 cycle path.
  //-----------------------------------------------------------------------------
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          wdata_r <= 0;
      else if (wdata_valid)
          //don't latch in data unless it's valid
          wdata_r <= wdata;

    end


  //Concatenate the rising and falling edge data to make a single bus
  assign dq_captured_0 = {dq_captured_falling, dq_captured_rising};

  //Apply delays in 1 chunks to avoid having to use transport delays
  assign #2500 delayed_dq_captured = dq_captured_0;

  //-----------------------------------------------------------------------------
  //Resynchronisation registers
  //These registers resychronise the captured read data from the DQS clock
  //domain back into an internal PLL clock domain. 
  //-----------------------------------------------------------------------------
  //Use a rising edge for resynch
  always @(posedge resynch_clk or negedge reset_n)
    begin
      if (reset_n == 0)
          resynched_data <= 0;
      else 
        resynched_data <= delayed_dq_captured;
    end


  //don't insert pipeline registers
  assign inter_rdata = resynched_data;

  //don't insert pipeline registers
  assign rdata = inter_rdata;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  stratixii_io dqs_io
    (
      .areset (1'b1),
      .combout (undelayed_dqs),
      .datain (dqs_oe_r),
      .ddiodatain (ZEROS[0]),
      .ddioinclk (),
      .ddioregout (),
      .delayctrlin (dqs_delay_ctrl),
      .devclrn (),
      .devoe (),
      .devpor (),
      .dqsbusout (dqs_clk),
      .dqsupdateen (dqsupdate),
      .inclk (not_dqs_clk),
      .inclkena (1'b1),
      .linkin (),
      .linkout (),
      .oe (dqs_oe),
      .offsetctrlin (),
      .outclk (clk),
      .outclkena (1'b1),
      .padio (ddr_dqs),
      .regout (),
      .sreset (),
      .terminationcontrol ()
    );

  defparam dqs_io.bus_hold = "false",
           dqs_io.ddio_mode = "output",
           dqs_io.ddioinclk_input = "inclk",
           dqs_io.dqs_ctrl_latches_enable = "true",
           dqs_io.dqs_delay_buffer_mode = gSTRATIXII_DLL_DELAY_BUFFER_MODE,
           dqs_io.dqs_edge_detect_enable = "false",
           dqs_io.dqs_input_frequency = gDLL_INPUT_FREQUENCY,
           dqs_io.dqs_offsetctrl_enable = "false",
           dqs_io.dqs_out_mode = gSTRATIXII_DQS_OUT_MODE,
           dqs_io.dqs_phase_shift = 6000,
           dqs_io.extend_oe_disable = "true",
           dqs_io.gated_dqs = "true",
           dqs_io.inclk_input = "dqs_bus",
           dqs_io.input_async_reset = "preset",
           dqs_io.input_power_up = "high",
           dqs_io.input_register_mode = "register",
           dqs_io.input_sync_reset = "clear",
           dqs_io.lpm_type = "stratixii_io",
           dqs_io.oe_async_reset = "none",
           dqs_io.oe_power_up = "low",
           dqs_io.oe_register_mode = "register",
           dqs_io.oe_sync_reset = "none",
           dqs_io.open_drain_output = "false",
           dqs_io.operation_mode = "bidir",
           dqs_io.output_async_reset = "none",
           dqs_io.output_power_up = "low",
           dqs_io.output_register_mode = "register",
           dqs_io.output_sync_reset = "none",
           dqs_io.sim_dqs_delay_increment = 36,
           dqs_io.sim_dqs_intrinsic_delay = 900,
           dqs_io.sim_dqs_offset_increment = 0,
           dqs_io.tie_off_oe_clock_enable = "false",
           dqs_io.tie_off_output_clock_enable = "false";


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  stratixii_io dqs_io
//    (
//      .areset (dq_enable_reset),
//      .combout (undelayed_dqs),
//      .datain (dqs_oe_r),
//      .ddiodatain (ZEROS[0]),
//      .ddioinclk (),
//      .ddioregout (),
//      .delayctrlin (dqs_delay_ctrl),
//      .devclrn (),
//      .devoe (),
//      .devpor (),
//      .dqsbusout (dqs_clk),
//      .dqsupdateen (dqsupdate),
//      .inclk (not_dqs_clk),
//      .inclkena (1'b1),
//      .linkin (),
//      .linkout (),
//      .oe (dqs_oe),
//      .offsetctrlin (),
//      .outclk (clk),
//      .outclkena (1'b1),
//      .padio (ddr_dqs),
//      .regout (),
//      .sreset (1'b1),
//      .terminationcontrol ()
//    );
//
//  defparam dqs_io.bus_hold = "false",
//           dqs_io.ddio_mode = "output",
//           dqs_io.ddioinclk_input = "negated_inclk",
//           dqs_io.dqs_ctrl_latches_enable = "true",
//           dqs_io.dqs_delay_buffer_mode = gSTRATIXII_DLL_DELAY_BUFFER_MODE,
//           dqs_io.dqs_edge_detect_enable = "false",
//           dqs_io.dqs_input_frequency = gDLL_INPUT_FREQUENCY,
//           dqs_io.dqs_offsetctrl_enable = "false",
//           dqs_io.dqs_out_mode = gSTRATIXII_DQS_OUT_MODE,
//           dqs_io.dqs_phase_shift = 6000,
//           dqs_io.extend_oe_disable = "true",
//           dqs_io.gated_dqs = "true",
//           dqs_io.inclk_input = "dqs_bus",
//           dqs_io.input_async_reset = "preset",
//           dqs_io.input_power_up = "high",
//           dqs_io.input_register_mode = "register",
//           dqs_io.input_sync_reset = "clear",
//           dqs_io.lpm_type = "stratixii_io",
//           dqs_io.oe_async_reset = "none",
//           dqs_io.oe_power_up = "low",
//           dqs_io.oe_register_mode = "register",
//           dqs_io.oe_sync_reset = "none",
//           dqs_io.open_drain_output = "false",
//           dqs_io.operation_mode = "bidir",
//           dqs_io.output_async_reset = "none",
//           dqs_io.output_power_up = "low",
//           dqs_io.output_register_mode = "register",
//           dqs_io.output_sync_reset = "none",
//           dqs_io.sim_dqs_delay_increment = 36,
//           dqs_io.sim_dqs_intrinsic_delay = 900,
//           dqs_io.sim_dqs_offset_increment = 0,
//           dqs_io.tie_off_oe_clock_enable = "false",
//           dqs_io.tie_off_output_clock_enable = "false";
//
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20471 "custom_dma.v" 2 */
/* SLline 1 "ddr_sdram_auk_ddr_clk_gen.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ps / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//----------------------------------------------------------------------------------
//Parameters:
//Number of memory clock output pairs    : 1
//----------------------------------------------------------------------------------

module ddr_sdram_auk_ddr_clk_gen (
                                   // inputs:
                                    clk,
                                    reset_n,

                                   // outputs:
                                    clk_to_sdram,
                                    clk_to_sdram_n
                                 )
;

  output           clk_to_sdram;
  output           clk_to_sdram_n;
  input            clk;
  input            reset_n;

  wire             clk_n;
  wire             clk_to_sdram;
  wire             clk_to_sdram_n;
  wire             gnd_signal;
  wire             vcc_signal;
  assign clk_n = ~clk;
  assign vcc_signal = {1{1'b1}};
  assign gnd_signal = 0;
  //------------------------------------------------------------
  //Stratix/Cyclone can drive clocks out on normal pins using
  //ALTDDIO_OUT megafunction
  //------------------------------------------------------------
  //Instantiate DDR IOs for driving the SDRAM clock off-chip

  altddio_out ddr_clk_out_p
    (
      .aclr (),
      .aset (),
      .datain_h (gnd_signal),
      .datain_l (vcc_signal),
      .dataout (clk_to_sdram),
      .oe (),
      .outclock (clk_n),
      .outclocken ()
    );

  defparam ddr_clk_out_p.extend_oe_disable = "UNUSED",
           ddr_clk_out_p.intended_device_family = "Stratix II",
           ddr_clk_out_p.invert_output = "OFF",
           ddr_clk_out_p.lpm_hint = "UNUSED",
           ddr_clk_out_p.lpm_type = "altddio_out",
           ddr_clk_out_p.oe_reg = "UNUSED",
           ddr_clk_out_p.power_up_high = "OFF",
           ddr_clk_out_p.width = 1;

  altddio_out ddr_clk_out_n
    (
      .aclr (),
      .aset (),
      .datain_h (gnd_signal),
      .datain_l (vcc_signal),
      .dataout (clk_to_sdram_n),
      .oe (),
      .outclock (clk),
      .outclocken ()
    );

  defparam ddr_clk_out_n.extend_oe_disable = "UNUSED",
           ddr_clk_out_n.intended_device_family = "Stratix II",
           ddr_clk_out_n.invert_output = "OFF",
           ddr_clk_out_n.lpm_hint = "UNUSED",
           ddr_clk_out_n.lpm_type = "altddio_out",
           ddr_clk_out_n.oe_reg = "UNUSED",
           ddr_clk_out_n.power_up_high = "OFF",
           ddr_clk_out_n.width = 1;


endmodule


/* SLline 20472 "custom_dma.v" 2 */
/* SLline 1 "ddr_sdram_auk_ddr_datapath.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ps / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_auk_ddr_datapath (
                                    // inputs:
                                     capture_clk,
                                     clk,
                                     control_be,
                                     control_doing_rd,
                                     control_doing_wr,
                                     control_dqs_burst,
                                     control_wdata,
                                     control_wdata_valid,
                                     dqs_delay_ctrl,
                                     dqsupdate,
                                     postamble_clk,
                                     reset_n,
                                     resynch_clk,
                                     write_clk,

                                    // outputs:
                                     clk_to_sdram,
                                     clk_to_sdram_n,
                                     control_rdata,
                                     ddr_dm,
                                     ddr_dq,
                                     ddr_dqs
                                  )
;

  parameter gstratixii_dqs_phase = 6000;
  parameter gstratixii_dqs_out_mode = "delay_chain2";
  parameter gstratixii_dll_delay_buffer_mode = "low";


  output           clk_to_sdram;
  output           clk_to_sdram_n;
  output  [ 31: 0] control_rdata;
  output  [  1: 0] ddr_dm;
  inout   [ 15: 0] ddr_dq;
  inout   [  1: 0] ddr_dqs;
  input            capture_clk;
  input            clk;
  input   [  3: 0] control_be;
  input            control_doing_rd;
  input            control_doing_wr;
  input            control_dqs_burst;
  input   [ 31: 0] control_wdata;
  input            control_wdata_valid;
  input   [  5: 0] dqs_delay_ctrl;
  input            dqsupdate;
  input            postamble_clk;
  input            reset_n;
  input            resynch_clk;
  input            write_clk;

  wire    [  3: 0] be_temp;
  wire             capture_clk_int;
  wire             clk_to_sdram;
  wire             clk_to_sdram_n;
  wire    [ 31: 0] control_rdata;
  wire    [  1: 0] ddr_dm;
  wire    [ 15: 0] ddr_dq;
  wire    [  1: 0] ddr_dqs;
  wire             postamble_clk_int;
  wire    [ 31: 0] rdata_temp;
  wire             resynch_clk_int;
  wire    [ 31: 0] wdata_temp;
  wire             write_clk_int;
  //
  //************************
  // Clock generator module 
  ddr_sdram_auk_ddr_clk_gen ddr_clk_gen
    (
      .clk (clk),
      .clk_to_sdram (clk_to_sdram),
      .clk_to_sdram_n (clk_to_sdram_n),
      .reset_n (reset_n)
    );


  //
  //**********************************
  // DQS group instantiation for dqs[0] 
  assign wdata_temp[15 : 0] = {control_wdata[23 : 16],control_wdata[7 : 0]};
  assign control_rdata[23 : 16] = rdata_temp[15 : 8];
  assign control_rdata[7 : 0] = rdata_temp[7 : 0];
  assign be_temp[1 : 0] = {control_be[2], control_be[0]};
  ddr_sdram_auk_ddr_dqs_group ^^^$_g_datapath:0:g_ddr_io_$^^^
    (
      .capture_clk (capture_clk_int),
      .clk (clk),
      .control_be (be_temp[1 : 0]),
      .control_doing_rd (control_doing_rd),
      .control_doing_wr (control_doing_wr),
      .control_dqs_burst (control_dqs_burst),
      .control_rdata (rdata_temp[15 : 0]),
      .control_wdata (wdata_temp[15 : 0]),
      .control_wdata_valid (control_wdata_valid),
      .ddr_dm (ddr_dm[0]),
      .ddr_dq (ddr_dq[7 : 0]),
      .ddr_dqs (ddr_dqs[0]),
      .dqs_delay_ctrl (dqs_delay_ctrl),
      .dqsupdate (dqsupdate),
      .postamble_clk (postamble_clk_int),
      .reset_n (reset_n),
      .resynch_clk (resynch_clk_int),
      .write_clk (write_clk_int)
    );

  defparam ^^^$_g_datapath:0:g_ddr_io_$^^^.gDLL_INPUT_FREQUENCY = "10000ps",
           ^^^$_g_datapath:0:g_ddr_io_$^^^.gSTRATIXII_DLL_DELAY_BUFFER_MODE = "low",
           ^^^$_g_datapath:0:g_ddr_io_$^^^.gSTRATIXII_DQS_OUT_MODE = "delay_chain2";

  //
  //**********************************
  // DQS group instantiation for dqs[1] 
  assign wdata_temp[31 : 16] = {control_wdata[31 : 24],control_wdata[15 : 8]};
  assign control_rdata[31 : 24] = rdata_temp[31 : 24];
  assign control_rdata[15 : 8] = rdata_temp[23 : 16];
  assign be_temp[3 : 2] = {control_be[3], control_be[1]};
  ddr_sdram_auk_ddr_dqs_group ^^^$_g_datapath:1:g_ddr_io_$^^^
    (
      .capture_clk (capture_clk_int),
      .clk (clk),
      .control_be (be_temp[3 : 2]),
      .control_doing_rd (control_doing_rd),
      .control_doing_wr (control_doing_wr),
      .control_dqs_burst (control_dqs_burst),
      .control_rdata (rdata_temp[31 : 16]),
      .control_wdata (wdata_temp[31 : 16]),
      .control_wdata_valid (control_wdata_valid),
      .ddr_dm (ddr_dm[1]),
      .ddr_dq (ddr_dq[15 : 8]),
      .ddr_dqs (ddr_dqs[1]),
      .dqs_delay_ctrl (dqs_delay_ctrl),
      .dqsupdate (dqsupdate),
      .postamble_clk (postamble_clk_int),
      .reset_n (reset_n),
      .resynch_clk (resynch_clk_int),
      .write_clk (write_clk_int)
    );

  defparam ^^^$_g_datapath:1:g_ddr_io_$^^^.gDLL_INPUT_FREQUENCY = "10000ps",
           ^^^$_g_datapath:1:g_ddr_io_$^^^.gSTRATIXII_DLL_DELAY_BUFFER_MODE = "low",
           ^^^$_g_datapath:1:g_ddr_io_$^^^.gSTRATIXII_DQS_OUT_MODE = "delay_chain2";


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign #2500 write_clk_int = ~clk;
  assign resynch_clk_int = resynch_clk;
  assign postamble_clk_int = postamble_clk;
  assign capture_clk_int = capture_clk;

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  assign write_clk_int = write_clk;
//  assign resynch_clk_int = resynch_clk;
//  assign postamble_clk_int = postamble_clk;
//  assign capture_clk_int = capture_clk;
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20473 "custom_dma.v" 2 */
/* SLline 1 "pll.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pll (
             // inputs:
              address,
              chipselect,
              clk,
              read,
              reset_n,
              write,
              writedata,

             // outputs:
              c0,
              c1,
              c2,
              readdata,
              resetrequest
           )
;

  output           c0;
  output           c1;
  output           c2;
  output  [ 15: 0] readdata;
  output           resetrequest;
  input   [  2: 0] address;
  input            chipselect;
  input            clk;
  input            read;
  input            reset_n;
  input            write;
  input   [ 15: 0] writedata;

  wire             always_one;
  wire             areset_n;
  wire             c0;
  wire             c1;
  wire             c2;
  wire             control_reg_en;
  wire    [ 15: 0] control_reg_in;
  reg     [ 15: 0] control_reg_out;
  reg              count_done;
  reg     [  5: 0] countup;
  wire             inclk0;
  reg              not_areset /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  wire    [ 15: 0] readdata;
  wire             resetrequest;
  wire    [ 15: 0] status_reg_in;
  reg     [ 15: 0] status_reg_out;
initial
  begin
    countup = 1'b0;
    count_done = 1'b0;
    not_areset = 1'b0;
  end
  assign status_reg_in[15 : 1] = 15'b000000000000000;
  assign resetrequest = ~count_done;
  //Up counter that stops counting when it reaches max value
  always @(posedge clk or negedge areset_n)
    begin
      if (areset_n == 0)
          countup <= 0;
      else if (count_done != 1'b1)
          countup <= countup + 1;
    end


  //Count_done signal, which is also the resetrequest_n
  always @(posedge clk or negedge areset_n)
    begin
      if (areset_n == 0)
          count_done <= 0;
      else if (countup == 6'b111111)
          count_done <= 1'b1;
    end


  //Creates a reset generator that will reset internal counters that are independent of global system reset
  always @(posedge clk or negedge 1'b1)
    begin
      if (1'b1 == 0)
          not_areset <= 0;
      else 
        not_areset <= always_one;
    end


  assign always_one = 1'b1;
  assign status_reg_in[0] = 1'b0;
  assign areset_n = not_areset;
  assign inclk0 = clk;
  //Mux status and control registers to the readdata output using address as select
  assign readdata = (address[0] == 0)? status_reg_out :
    ({control_reg_out[15 : 2], ~control_reg_out[1], control_reg_out[0]} );

  //Status register - Read-Only
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          status_reg_out <= 0;
      else 
        status_reg_out <= status_reg_in;
    end


  //Control register - R/W
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          control_reg_out <= 0;
      else if (control_reg_en)
          control_reg_out <= {control_reg_in[15 : 2], ~control_reg_in[1], control_reg_in[0]};
    end


  assign control_reg_in = writedata;
  assign control_reg_en = (address == 3'b001) && write && chipselect;
  //s1, which is an e_avalon_slave
  altpllpll the_pll
    (
      .c0 (c0),
      .c1 (c1),
      .c2 (c2),
      .inclk0 (inclk0)
    );



endmodule


/* SLline 20476 "custom_dma.v" 2 */
/* SLline 1 "altpllpll.v" 1 */
// megafunction wizard: %ALTPLL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altpll 

// ============================================================
// File Name: altpllpll.v
// Megafunction Name(s):
// 			altpll
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 345 02/24/2010 SP 2 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpllpll (
	inclk0,
	c0,
	c1,
	c2);

	input	  inclk0;
	output	  c0;
	output	  c1;
	output	  c2;

	wire [5:0] sub_wire0;
	wire [0:0] sub_wire6 = 1'h0;
	wire [2:2] sub_wire3 = sub_wire0[2:2];
	wire [1:1] sub_wire2 = sub_wire0[1:1];
	wire [0:0] sub_wire1 = sub_wire0[0:0];
	wire  c0 = sub_wire1;
	wire  c1 = sub_wire2;
	wire  c2 = sub_wire3;
	wire  sub_wire4 = inclk0;
	wire [1:0] sub_wire5 = {sub_wire6, sub_wire4};

	altpll	altpll_component (
				.inclk (sub_wire5),
				.clk (sub_wire0),
				.activeclock (),
				.areset (1'b0),
				.clkbad (),
				.clkena ({6{1'b1}}),
				.clkloss (),
				.clkswitch (1'b0),
				.configupdate (1'b0),
				.enable0 (),
				.enable1 (),
				.extclk (),
				.extclkena ({4{1'b1}}),
				.fbin (1'b1),
				.fbmimicbidir (),
				.fbout (),
				.fref (),
				.icdrclk (),
				.locked (),
				.pfdena (1'b1),
				.phasecounterselect ({4{1'b1}}),
				.phasedone (),
				.phasestep (1'b1),
				.phaseupdown (1'b1),
				.pllena (1'b1),
				.scanaclr (1'b0),
				.scanclk (1'b0),
				.scanclkena (1'b1),
				.scandata (1'b0),
				.scandataout (),
				.scandone (),
				.scanread (1'b0),
				.scanwrite (1'b0),
				.sclkout0 (),
				.sclkout1 (),
				.vcooverrange (),
				.vcounderrange ());
	defparam
		altpll_component.bandwidth_type = "AUTO",
		altpll_component.clk0_divide_by = 1,
		altpll_component.clk0_duty_cycle = 50,
		altpll_component.clk0_multiply_by = 2,
		altpll_component.clk0_phase_shift = "0",
		altpll_component.clk1_divide_by = 1,
		altpll_component.clk1_duty_cycle = 50,
		altpll_component.clk1_multiply_by = 2,
		altpll_component.clk1_phase_shift = "-3380",
		altpll_component.clk2_divide_by = 1,
		altpll_component.clk2_duty_cycle = 50,
		altpll_component.clk2_multiply_by = 2,
		altpll_component.clk2_phase_shift = "7500",
		altpll_component.compensate_clock = "CLK0",
		altpll_component.inclk0_input_frequency = 20000,
		altpll_component.intended_device_family = "Stratix II",
		altpll_component.lpm_type = "altpll",
		altpll_component.operation_mode = "NORMAL",
		altpll_component.pll_type = "AUTO",
		altpll_component.port_activeclock = "PORT_UNUSED",
		altpll_component.port_areset = "PORT_UNUSED",
		altpll_component.port_clkbad0 = "PORT_UNUSED",
		altpll_component.port_clkbad1 = "PORT_UNUSED",
		altpll_component.port_clkloss = "PORT_UNUSED",
		altpll_component.port_clkswitch = "PORT_UNUSED",
		altpll_component.port_configupdate = "PORT_UNUSED",
		altpll_component.port_fbin = "PORT_UNUSED",
		altpll_component.port_inclk0 = "PORT_USED",
		altpll_component.port_inclk1 = "PORT_UNUSED",
		altpll_component.port_locked = "PORT_UNUSED",
		altpll_component.port_pfdena = "PORT_UNUSED",
		altpll_component.port_phasecounterselect = "PORT_UNUSED",
		altpll_component.port_phasedone = "PORT_UNUSED",
		altpll_component.port_phasestep = "PORT_UNUSED",
		altpll_component.port_phaseupdown = "PORT_UNUSED",
		altpll_component.port_pllena = "PORT_UNUSED",
		altpll_component.port_scanaclr = "PORT_UNUSED",
		altpll_component.port_scanclk = "PORT_UNUSED",
		altpll_component.port_scanclkena = "PORT_UNUSED",
		altpll_component.port_scandata = "PORT_UNUSED",
		altpll_component.port_scandataout = "PORT_UNUSED",
		altpll_component.port_scandone = "PORT_UNUSED",
		altpll_component.port_scanread = "PORT_UNUSED",
		altpll_component.port_scanwrite = "PORT_UNUSED",
		altpll_component.port_clk0 = "PORT_USED",
		altpll_component.port_clk1 = "PORT_USED",
		altpll_component.port_clk2 = "PORT_USED",
		altpll_component.port_clk3 = "PORT_UNUSED",
		altpll_component.port_clk4 = "PORT_UNUSED",
		altpll_component.port_clk5 = "PORT_UNUSED",
		altpll_component.port_clkena0 = "PORT_UNUSED",
		altpll_component.port_clkena1 = "PORT_UNUSED",
		altpll_component.port_clkena2 = "PORT_UNUSED",
		altpll_component.port_clkena3 = "PORT_UNUSED",
		altpll_component.port_clkena4 = "PORT_UNUSED",
		altpll_component.port_clkena5 = "PORT_UNUSED",
		altpll_component.port_enable0 = "PORT_UNUSED",
		altpll_component.port_enable1 = "PORT_UNUSED",
		altpll_component.port_extclk0 = "PORT_UNUSED",
		altpll_component.port_extclk1 = "PORT_UNUSED",
		altpll_component.port_extclk2 = "PORT_UNUSED",
		altpll_component.port_extclk3 = "PORT_UNUSED",
		altpll_component.port_sclkout0 = "PORT_UNUSED",
		altpll_component.port_sclkout1 = "PORT_UNUSED",
		altpll_component.spread_frequency = 0;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACTIVECLK_CHECK STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH STRING "1.000"
// Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT STRING "MHz"
// Retrieval info: PRIVATE: BANDWIDTH_PRESET STRING "Low"
// Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO STRING "1"
// Retrieval info: PRIVATE: BANDWIDTH_USE_CUSTOM STRING "0"
// Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET STRING "0"
// Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKLOSS_CHECK STRING "0"
// Retrieval info: PRIVATE: CLKSWITCH_CHECK STRING "0"
// Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO STRING "0"
// Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK STRING "0"
// Retrieval info: PRIVATE: CREATE_INCLK1_CHECK STRING "0"
// Retrieval info: PRIVATE: CUR_DEDICATED_CLK STRING "c0"
// Retrieval info: PRIVATE: CUR_FBIN_CLK STRING "e0"
// Retrieval info: PRIVATE: DEVICE_SPEED_GRADE STRING "3"
// Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "1"
// Retrieval info: PRIVATE: DIV_FACTOR1 NUMERIC "1"
// Retrieval info: PRIVATE: DIV_FACTOR2 NUMERIC "1"
// Retrieval info: PRIVATE: DUTY_CYCLE0 STRING "50.00000000"
// Retrieval info: PRIVATE: DUTY_CYCLE1 STRING "50.00000000"
// Retrieval info: PRIVATE: DUTY_CYCLE2 STRING "50.00000000"
// Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE0 STRING "100.000000"
// Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE1 STRING "100.000000"
// Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE2 STRING "100.000000"
// Retrieval info: PRIVATE: EXPLICIT_SWITCHOVER_COUNTER STRING "0"
// Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO STRING "0"
// Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: GLOCKED_MODE_CHECK STRING "0"
// Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "1048575"
// Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER STRING "1"
// Retrieval info: PRIVATE: INCLK0_FREQ_EDIT STRING "50.000"
// Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT STRING "100.000"
// Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED STRING "1"
// Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO STRING "MHz"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK STRING "0"
// Retrieval info: PRIVATE: LONG_SCAN_RADIO STRING "1"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE STRING "150.000"
// Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
// Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 STRING "ps"
// Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT1 STRING "ps"
// Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT2 STRING "ps"
// Retrieval info: PRIVATE: MIG_DEVICE_SPEED_GRADE STRING "Any"
// Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "2"
// Retrieval info: PRIVATE: MULT_FACTOR1 NUMERIC "2"
// Retrieval info: PRIVATE: MULT_FACTOR2 NUMERIC "2"
// Retrieval info: PRIVATE: NORMAL_MODE_RADIO STRING "1"
// Retrieval info: PRIVATE: OUTPUT_FREQ0 STRING "100.00000000"
// Retrieval info: PRIVATE: OUTPUT_FREQ1 STRING "100.00000000"
// Retrieval info: PRIVATE: OUTPUT_FREQ2 STRING "100.00000000"
// Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 STRING "0"
// Retrieval info: PRIVATE: OUTPUT_FREQ_MODE1 STRING "0"
// Retrieval info: PRIVATE: OUTPUT_FREQ_MODE2 STRING "0"
// Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 STRING "MHz"
// Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT1 STRING "MHz"
// Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT2 STRING "MHz"
// Retrieval info: PRIVATE: PHASE_RECONFIG_FEATURE_ENABLED STRING "0"
// Retrieval info: PRIVATE: PHASE_RECONFIG_INPUTS_CHECK STRING "0"
// Retrieval info: PRIVATE: PHASE_SHIFT0 STRING "0.00000000"
// Retrieval info: PRIVATE: PHASE_SHIFT1 STRING "-3.38000000"
// Retrieval info: PRIVATE: PHASE_SHIFT2 STRING "270.00000000"
// Retrieval info: PRIVATE: PHASE_SHIFT_STEP_ENABLED_CHECK STRING "0"
// Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 STRING "ps"
// Retrieval info: PRIVATE: PHASE_SHIFT_UNIT1 STRING "ns"
// Retrieval info: PRIVATE: PHASE_SHIFT_UNIT2 STRING "deg"
// Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ARESET_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "1"
// Retrieval info: PRIVATE: PLL_ENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_FBMIMIC_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PLL_PFDENA_CHECK STRING "0"
// Retrieval info: PRIVATE: PLL_TARGET_HARCOPY_CHECK NUMERIC "0"
// Retrieval info: PRIVATE: PRIMARY_CLK_COMBO STRING "inclk0"
// Retrieval info: PRIVATE: RECONFIG_FILE STRING "altpllpll.mif"
// Retrieval info: PRIVATE: SACN_INPUTS_CHECK STRING "0"
// Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SELF_RESET_LOCK_LOSS STRING "0"
// Retrieval info: PRIVATE: SHORT_SCAN_RADIO STRING "0"
// Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SPREAD_FREQ STRING "50.000"
// Retrieval info: PRIVATE: SPREAD_FREQ_UNIT STRING "KHz"
// Retrieval info: PRIVATE: SPREAD_PERCENT STRING "0.500"
// Retrieval info: PRIVATE: SPREAD_USE STRING "0"
// Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO STRING "0"
// Retrieval info: PRIVATE: STICKY_CLK0 STRING "1"
// Retrieval info: PRIVATE: STICKY_CLK1 STRING "1"
// Retrieval info: PRIVATE: STICKY_CLK2 STRING "1"
// Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
// Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED STRING "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USE_CLK0 STRING "1"
// Retrieval info: PRIVATE: USE_CLK1 STRING "1"
// Retrieval info: PRIVATE: USE_CLK2 STRING "1"
// Retrieval info: PRIVATE: USE_MIL_SPEED_GRADE NUMERIC "0"
// Retrieval info: PRIVATE: ZERO_DELAY_RADIO STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: BANDWIDTH_TYPE STRING "AUTO"
// Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
// Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "2"
// Retrieval info: CONSTANT: CLK0_PHASE_SHIFT STRING "0"
// Retrieval info: CONSTANT: CLK1_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: CLK1_DUTY_CYCLE NUMERIC "50"
// Retrieval info: CONSTANT: CLK1_MULTIPLY_BY NUMERIC "2"
// Retrieval info: CONSTANT: CLK1_PHASE_SHIFT STRING "-3380"
// Retrieval info: CONSTANT: CLK2_DIVIDE_BY NUMERIC "1"
// Retrieval info: CONSTANT: CLK2_DUTY_CYCLE NUMERIC "50"
// Retrieval info: CONSTANT: CLK2_MULTIPLY_BY NUMERIC "2"
// Retrieval info: CONSTANT: CLK2_PHASE_SHIFT STRING "7500"
// Retrieval info: CONSTANT: COMPENSATE_CLOCK STRING "CLK0"
// Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "20000"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altpll"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "NORMAL"
// Retrieval info: CONSTANT: PLL_TYPE STRING "AUTO"
// Retrieval info: CONSTANT: PORT_ACTIVECLOCK STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_ARESET STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_CLKBAD0 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_CLKBAD1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_CLKLOSS STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_CLKSWITCH STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_CONFIGUPDATE STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_FBIN STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_INCLK0 STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_INCLK1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_LOCKED STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PFDENA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PHASECOUNTERSELECT STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PHASEDONE STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PHASESTEP STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PHASEUPDOWN STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_PLLENA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANACLR STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANCLK STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANCLKENA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANDATA STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANDATAOUT STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANDONE STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANREAD STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_SCANWRITE STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clk0 STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_clk1 STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_clk2 STRING "PORT_USED"
// Retrieval info: CONSTANT: PORT_clk3 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clk4 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clk5 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena0 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena2 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena3 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena4 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_clkena5 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_enable0 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_enable1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_extclk0 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_extclk1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_extclk2 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_extclk3 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_sclkout0 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_sclkout1 STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: SPREAD_FREQUENCY NUMERIC "0"
// Retrieval info: USED_PORT: @clk 0 0 6 0 OUTPUT_CLK_EXT VCC "@clk[5..0]"
// Retrieval info: USED_PORT: @extclk 0 0 4 0 OUTPUT_CLK_EXT VCC "@extclk[3..0]"
// Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT_CLK_EXT VCC "c0"
// Retrieval info: USED_PORT: c1 0 0 0 0 OUTPUT_CLK_EXT VCC "c1"
// Retrieval info: USED_PORT: c2 0 0 0 0 OUTPUT_CLK_EXT VCC "c2"
// Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT_CLK_EXT GND "inclk0"
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
// Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
// Retrieval info: CONNECT: c1 0 0 0 0 @clk 0 0 1 1
// Retrieval info: CONNECT: c2 0 0 0 0 @clk 0 0 1 2
// Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpllpll_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf

/* SLline 20477 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_2.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: cpu/data_master
//adapter masters: pipeline_bridge/s1
//asp_debug: 0
//byteaddr_width: 14
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 4
//downstream_addr_shift: 2
//downstream_burstcount_width: 1
//downstream_max_burstcount: 1
//downstream_pipeline: 1
//dynamic_slave: 1
//master_always_burst_max_burst: 0
//master_burst_on_burst_boundaries_only: 1
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 0
//nativeaddr_width: 12
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 0
//upstream_burstcount: upstream_burstcount
//upstream_burstcount_width: 4
//upstream_max_burstcount: 8
//zero_address_width: 0


module custom_dma_burst_2 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_burstcount,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             reg_downstream_address,
                             reg_downstream_arbitrationshare,
                             reg_downstream_burstcount,
                             reg_downstream_byteenable,
                             reg_downstream_debugaccess,
                             reg_downstream_nativeaddress,
                             reg_downstream_read,
                             reg_downstream_write,
                             reg_downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 11: 0] reg_downstream_address;
  output  [  3: 0] reg_downstream_arbitrationshare;
  output           reg_downstream_burstcount;
  output  [  3: 0] reg_downstream_byteenable;
  output           reg_downstream_debugaccess;
  output  [ 11: 0] reg_downstream_nativeaddress;
  output           reg_downstream_read;
  output           reg_downstream_write;
  output  [ 31: 0] reg_downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 13: 0] upstream_address;
  input   [  3: 0] upstream_burstcount;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 11: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  2: 0] address_offset;
  reg              atomic_counter;
  wire    [ 13: 0] current_upstream_address;
  wire    [  3: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  3: 0] data_counter;
  wire    [  3: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 11: 0] downstream_address;
  wire    [ 13: 0] downstream_address_base;
  wire    [  3: 0] downstream_arbitrationshare;
  wire             downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 11: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire             max_burst_size;
  wire             p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  2: 0] read_address_offset;
  wire             read_update_count;
  wire    [  3: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 11: 0] reg_downstream_address;
  reg     [  3: 0] reg_downstream_arbitrationshare;
  reg              reg_downstream_burstcount;
  reg     [  3: 0] reg_downstream_byteenable;
  reg              reg_downstream_debugaccess;
  reg     [ 11: 0] reg_downstream_nativeaddress;
  reg              reg_downstream_read;
  reg              reg_downstream_write;
  reg     [ 31: 0] reg_downstream_writedata;
  reg     [  3: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 13: 0] registered_upstream_address;
  reg     [  3: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 11: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  3: 0] transactions_remaining;
  reg     [  3: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  2: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= upstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? upstream_burstcount : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 1;
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign downstream_arbitrationshare = current_upstream_read ? (dbs_adjusted_upstream_burstcount) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign downstream_address = downstream_address_base + {address_offset, 2'b00};
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_address <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_address <= downstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_arbitrationshare <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_arbitrationshare <= downstream_arbitrationshare;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_burstcount <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_burstcount <= downstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_byteenable <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_byteenable <= downstream_byteenable;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_debugaccess <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_debugaccess <= downstream_debugaccess;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_nativeaddress <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_nativeaddress <= downstream_nativeaddress;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_read <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_read <= downstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_write <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_write <= downstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_writedata <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_writedata <= downstream_writedata;
    end



endmodule


/* SLline 20478 "custom_dma.v" 2 */
/* SLline 1 "sysid.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sysid (
               // inputs:
                address,

               // outputs:
                readdata
             )
;

  output  [ 31: 0] readdata;
  input            address;

  wire    [ 31: 0] readdata;
  //control_slave, which is an e_avalon_slave
  assign readdata = address ? 1271845543 : 2057062574;

endmodule


/* SLline 20479 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_5.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: fir_dma/write_master
//adapter masters: ddr_sdram/s1
//asp_debug: 0
//byteaddr_width: 27
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 3
//downstream_addr_shift: 2
//downstream_burstcount_width: 3
//downstream_max_burstcount: 4
//downstream_pipeline: 0
//dynamic_slave: 1
//master_always_burst_max_burst: 0
//master_burst_on_burst_boundaries_only: 0
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 0
//nativeaddr_width: 25
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 1
//upstream_burstcount: upstream_burstcount
//upstream_burstcount_width: 3
//upstream_max_burstcount: 4
//zero_address_width: 0


module custom_dma_burst_5 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_burstcount,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             downstream_address,
                             downstream_arbitrationshare,
                             downstream_burstcount,
                             downstream_byteenable,
                             downstream_debugaccess,
                             downstream_nativeaddress,
                             downstream_read,
                             downstream_write,
                             downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 24: 0] downstream_address;
  output  [  2: 0] downstream_arbitrationshare;
  output  [  2: 0] downstream_burstcount;
  output  [  3: 0] downstream_byteenable;
  output           downstream_debugaccess;
  output  [ 24: 0] downstream_nativeaddress;
  output           downstream_read;
  output           downstream_write;
  output  [ 31: 0] downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 26: 0] upstream_address;
  input   [  2: 0] upstream_burstcount;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 24: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  1: 0] address_offset;
  reg     [  2: 0] atomic_counter;
  wire    [ 26: 0] current_upstream_address;
  wire    [  2: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  2: 0] data_counter;
  wire    [  2: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 24: 0] downstream_address;
  wire    [ 26: 0] downstream_address_base;
  wire    [  2: 0] downstream_arbitrationshare;
  wire    [  2: 0] downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 24: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire    [  2: 0] interleave_end;
  wire    [  2: 0] max_burst_size;
  wire    [  2: 0] p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  1: 0] read_address_offset;
  wire             read_update_count;
  wire    [  2: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [  2: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 26: 0] registered_upstream_address;
  reg     [  2: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 24: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  2: 0] transactions_remaining;
  reg     [  2: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  1: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= upstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? upstream_burstcount : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 4;
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign interleave_end = (dbs_adjusted_upstream_burstcount > 0) ? (dbs_adjusted_upstream_burstcount - 0) : 0;
  assign downstream_arbitrationshare = current_upstream_read ? (0 + (interleave_end >> 2) + |(interleave_end[1 : 0])) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign downstream_address = downstream_address_base + {address_offset, 2'b00};
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;

endmodule


/* SLline 20480 "custom_dma.v" 2 */
/* SLline 1 "jtag_uart.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_log_module (
                              // inputs:
                               clk,
                               data,
                               strobe,
                               valid
                            )
;

  input            clk;
  input   [  7: 0] data;
  input            strobe;
  input            valid;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
   reg [31:0] text_handle; // for $fopen
   initial text_handle = $fopen ("C:/Projects/10/accelerated_fir_dma_cleanup/Custom_FIR_DMA/StratixII/custom_dma_sim/jtag_uart_output_stream.dat");

   always @(posedge clk) begin
      if (valid && strobe) begin
	 $fwrite (text_handle, "%b\n", data);
          // echo raw binary strings to file as ascii to screen
         $write("%s", ((data == 8'hd) ? 8'ha : data));
                     
	 // non-standard; poorly documented; required to get real data stream.
	 $fflush (text_handle);
      end
   end // clk


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_sim_scfifo_w (
                                // inputs:
                                 clk,
                                 fifo_wdata,
                                 fifo_wr,

                                // outputs:
                                 fifo_FF,
                                 r_dat,
                                 wfifo_empty,
                                 wfifo_used
                              )
;

  output           fifo_FF;
  output  [  7: 0] r_dat;
  output           wfifo_empty;
  output  [  5: 0] wfifo_used;
  input            clk;
  input   [  7: 0] fifo_wdata;
  input            fifo_wr;

  wire             fifo_FF;
  wire    [  7: 0] r_dat;
  wire             wfifo_empty;
  wire    [  5: 0] wfifo_used;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_log, which is an e_log
  jtag_uart_log_module jtag_uart_log
    (
      .clk    (clk),
      .data   (fifo_wdata),
      .strobe (fifo_wr),
      .valid  (fifo_wr)
    );

  assign wfifo_used = {6{1'b0}};
  assign r_dat = {8{1'b0}};
  assign fifo_FF = 1'b0;
  assign wfifo_empty = 1'b1;

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_scfifo_w (
                            // inputs:
                             clk,
                             fifo_clear,
                             fifo_wdata,
                             fifo_wr,
                             rd_wfifo,

                            // outputs:
                             fifo_FF,
                             r_dat,
                             wfifo_empty,
                             wfifo_used
                          )
;

  output           fifo_FF;
  output  [  7: 0] r_dat;
  output           wfifo_empty;
  output  [  5: 0] wfifo_used;
  input            clk;
  input            fifo_clear;
  input   [  7: 0] fifo_wdata;
  input            fifo_wr;
  input            rd_wfifo;

  wire             fifo_FF;
  wire    [  7: 0] r_dat;
  wire             wfifo_empty;
  wire    [  5: 0] wfifo_used;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  jtag_uart_sim_scfifo_w the_jtag_uart_sim_scfifo_w
    (
      .clk         (clk),
      .fifo_FF     (fifo_FF),
      .fifo_wdata  (fifo_wdata),
      .fifo_wr     (fifo_wr),
      .r_dat       (r_dat),
      .wfifo_empty (wfifo_empty),
      .wfifo_used  (wfifo_used)
    );


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  scfifo wfifo
//    (
//      .aclr (fifo_clear),
//      .clock (clk),
//      .data (fifo_wdata),
//      .empty (wfifo_empty),
//      .full (fifo_FF),
//      .q (r_dat),
//      .rdreq (rd_wfifo),
//      .usedw (wfifo_used),
//      .wrreq (fifo_wr)
//    );
//
//  defparam wfifo.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
//           wfifo.lpm_numwords = 64,
//           wfifo.lpm_showahead = "OFF",
//           wfifo.lpm_type = "scfifo",
//           wfifo.lpm_width = 8,
//           wfifo.lpm_widthu = 6,
//           wfifo.overflow_checking = "OFF",
//           wfifo.underflow_checking = "OFF",
//           wfifo.use_eab = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_drom_module (
                               // inputs:
                                clk,
                                incr_addr,
                                reset_n,

                               // outputs:
                                new_rom,
                                num_bytes,
                                q,
                                safe
                             )
;

  parameter POLL_RATE = 100;


  output           new_rom;
  output  [ 31: 0] num_bytes;
  output  [  7: 0] q;
  output           safe;
  input            clk;
  input            incr_addr;
  input            reset_n;

  reg     [ 11: 0] address;
  reg              d1_pre;
  reg              d2_pre;
  reg              d3_pre;
  reg              d4_pre;
  reg              d5_pre;
  reg              d6_pre;
  reg              d7_pre;
  reg              d8_pre;
  reg              d9_pre;
  reg     [  7: 0] mem_array [2047: 0];
  reg     [ 31: 0] mutex [  1: 0];
  reg              new_rom;
  wire    [ 31: 0] num_bytes;
  reg              pre;
  wire    [  7: 0] q;
  wire             safe;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign q = mem_array[address];
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
          d1_pre <= 0;
          d2_pre <= 0;
          d3_pre <= 0;
          d4_pre <= 0;
          d5_pre <= 0;
          d6_pre <= 0;
          d7_pre <= 0;
          d8_pre <= 0;
          d9_pre <= 0;
          new_rom <= 0;
        end
      else 
        begin
          d1_pre <= pre;
          d2_pre <= d1_pre;
          d3_pre <= d2_pre;
          d4_pre <= d3_pre;
          d5_pre <= d4_pre;
          d6_pre <= d5_pre;
          d7_pre <= d6_pre;
          d8_pre <= d7_pre;
          d9_pre <= d8_pre;
          new_rom <= d9_pre;
        end
    end



   assign     num_bytes = mutex[1];
                   reg        safe_delay;
   reg [31:0] poll_count;
   reg [31:0] mutex_handle;
   wire       interactive = 1'b0 ; // '
   assign     safe = (address < mutex[1]);

   initial poll_count = POLL_RATE;

   always @(posedge clk or negedge reset_n) begin
      if (reset_n !== 1) begin
         safe_delay <= 0;
      end else begin
         safe_delay <= safe;
      end
   end // safe_delay

   always @(posedge clk or negedge reset_n) begin
      if (reset_n !== 1) begin  // dont worry about null _stream.dat file
         address <= 0;
         mem_array[0] <= 0;
         mutex[0] <= 0;
         mutex[1] <= 0;
         pre <= 0;
      end else begin            // deal with the non-reset case
         pre <= 0;
         if (incr_addr && safe) address <= address + 1;
         if (mutex[0] && !safe && safe_delay) begin
            // and blast the mutex after falling edge of safe if interactive
            if (interactive) begin
               mutex_handle = $fopen ("C:/Projects/10/accelerated_fir_dma_cleanup/Custom_FIR_DMA/StratixII/custom_dma_sim/jtag_uart_input_mutex.dat");
               $fdisplay (mutex_handle, "0");
               $fclose (mutex_handle);
               // $display ($stime, "\t%m:\n\t\tMutex cleared!");
            end else begin
               // sleep until next reset, do not bash mutex.
               wait (!reset_n);
            end
         end // OK to bash mutex.
         if (poll_count < POLL_RATE) begin // wait
            poll_count = poll_count + 1;
         end else begin         // do the interesting stuff.
            poll_count = 0;
            $readmemh ("C:/Projects/10/accelerated_fir_dma_cleanup/Custom_FIR_DMA/StratixII/custom_dma_sim/jtag_uart_input_mutex.dat", mutex);
            if (mutex[0] && !safe) begin
            // read stream into mem_array after current characters are gone!
               // save mutex[0] value to compare to address (generates 'safe')
               mutex[1] <= mutex[0];
               // $display ($stime, "\t%m:\n\t\tMutex hit: Trying to read %d bytes...", mutex[0]);
               $readmemb("C:/Projects/10/accelerated_fir_dma_cleanup/Custom_FIR_DMA/StratixII/custom_dma_sim/jtag_uart_input_stream.dat", mem_array);
               // bash address and send pulse outside to send the char:
               address <= 0;
               pre <= -1;
            end // else mutex miss...
         end // poll_count
      end // reset
   end // posedge clk


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_sim_scfifo_r (
                                // inputs:
                                 clk,
                                 fifo_rd,
                                 rst_n,

                                // outputs:
                                 fifo_EF,
                                 fifo_rdata,
                                 rfifo_full,
                                 rfifo_used
                              )
;

  output           fifo_EF;
  output  [  7: 0] fifo_rdata;
  output           rfifo_full;
  output  [  5: 0] rfifo_used;
  input            clk;
  input            fifo_rd;
  input            rst_n;

  reg     [ 31: 0] bytes_left;
  wire             fifo_EF;
  reg              fifo_rd_d;
  wire    [  7: 0] fifo_rdata;
  wire             new_rom;
  wire    [ 31: 0] num_bytes;
  wire    [  6: 0] rfifo_entries;
  wire             rfifo_full;
  wire    [  5: 0] rfifo_used;
  wire             safe;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_drom, which is an e_drom
  jtag_uart_drom_module jtag_uart_drom
    (
      .clk       (clk),
      .incr_addr (fifo_rd_d),
      .new_rom   (new_rom),
      .num_bytes (num_bytes),
      .q         (fifo_rdata),
      .reset_n   (rst_n),
      .safe      (safe)
    );

  // Generate rfifo_entries for simulation
  always @(posedge clk or negedge rst_n)
    begin
      if (rst_n == 0)
        begin
          bytes_left <= 32'h0;
          fifo_rd_d <= 1'b0;
        end
      else 
        begin
          fifo_rd_d <= fifo_rd;
          // decrement on read
          if (fifo_rd_d)
              bytes_left <= bytes_left - 1'b1;
          // catch new contents
          if (new_rom)
              bytes_left <= num_bytes;
        end
    end


  assign fifo_EF = bytes_left == 32'b0;
  assign rfifo_full = bytes_left > 7'h40;
  assign rfifo_entries = (rfifo_full) ? 7'h40 : bytes_left;
  assign rfifo_used = rfifo_entries[5 : 0];

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_scfifo_r (
                            // inputs:
                             clk,
                             fifo_clear,
                             fifo_rd,
                             rst_n,
                             t_dat,
                             wr_rfifo,

                            // outputs:
                             fifo_EF,
                             fifo_rdata,
                             rfifo_full,
                             rfifo_used
                          )
;

  output           fifo_EF;
  output  [  7: 0] fifo_rdata;
  output           rfifo_full;
  output  [  5: 0] rfifo_used;
  input            clk;
  input            fifo_clear;
  input            fifo_rd;
  input            rst_n;
  input   [  7: 0] t_dat;
  input            wr_rfifo;

  wire             fifo_EF;
  wire    [  7: 0] fifo_rdata;
  wire             rfifo_full;
  wire    [  5: 0] rfifo_used;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  jtag_uart_sim_scfifo_r the_jtag_uart_sim_scfifo_r
    (
      .clk        (clk),
      .fifo_EF    (fifo_EF),
      .fifo_rd    (fifo_rd),
      .fifo_rdata (fifo_rdata),
      .rfifo_full (rfifo_full),
      .rfifo_used (rfifo_used),
      .rst_n      (rst_n)
    );


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  scfifo rfifo
//    (
//      .aclr (fifo_clear),
//      .clock (clk),
//      .data (t_dat),
//      .empty (fifo_EF),
//      .full (rfifo_full),
//      .q (fifo_rdata),
//      .rdreq (fifo_rd),
//      .usedw (rfifo_used),
//      .wrreq (wr_rfifo)
//    );
//
//  defparam rfifo.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
//           rfifo.lpm_numwords = 64,
//           rfifo.lpm_showahead = "OFF",
//           rfifo.lpm_type = "scfifo",
//           rfifo.lpm_width = 8,
//           rfifo.lpm_widthu = 6,
//           rfifo.overflow_checking = "OFF",
//           rfifo.underflow_checking = "OFF",
//           rfifo.use_eab = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart (
                   // inputs:
                    av_address,
                    av_chipselect,
                    av_read_n,
                    av_write_n,
                    av_writedata,
                    clk,
                    rst_n,

                   // outputs:
                    av_irq,
                    av_readdata,
                    av_waitrequest,
                    dataavailable,
                    readyfordata
                 )
  /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"R101,C106,D101,D103\"" */ ;

  output           av_irq;
  output  [ 31: 0] av_readdata;
  output           av_waitrequest;
  output           dataavailable;
  output           readyfordata;
  input            av_address;
  input            av_chipselect;
  input            av_read_n;
  input            av_write_n;
  input   [ 31: 0] av_writedata;
  input            clk;
  input            rst_n;

  reg              ac;
  wire             activity;
  wire             av_irq;
  wire    [ 31: 0] av_readdata;
  reg              av_waitrequest;
  reg              dataavailable;
  reg              fifo_AE;
  reg              fifo_AF;
  wire             fifo_EF;
  wire             fifo_FF;
  wire             fifo_clear;
  wire             fifo_rd;
  wire    [  7: 0] fifo_rdata;
  wire    [  7: 0] fifo_wdata;
  reg              fifo_wr;
  reg              ien_AE;
  reg              ien_AF;
  wire             ipen_AE;
  wire             ipen_AF;
  reg              pause_irq;
  wire    [  7: 0] r_dat;
  wire             r_ena;
  reg              r_val;
  wire             rd_wfifo;
  reg              read_0;
  reg              readyfordata;
  wire             rfifo_full;
  wire    [  5: 0] rfifo_used;
  reg              rvalid;
  reg              sim_r_ena;
  reg              sim_t_dat;
  reg              sim_t_ena;
  reg              sim_t_pause;
  wire    [  7: 0] t_dat;
  reg              t_dav;
  wire             t_ena;
  wire             t_pause;
  wire             wfifo_empty;
  wire    [  5: 0] wfifo_used;
  reg              woverflow;
  wire             wr_rfifo;
  //avalon_jtag_slave, which is an e_avalon_slave
  assign rd_wfifo = r_ena & ~wfifo_empty;
  assign wr_rfifo = t_ena & ~rfifo_full;
  assign fifo_clear = ~rst_n;
  jtag_uart_scfifo_w the_jtag_uart_scfifo_w
    (
      .clk         (clk),
      .fifo_FF     (fifo_FF),
      .fifo_clear  (fifo_clear),
      .fifo_wdata  (fifo_wdata),
      .fifo_wr     (fifo_wr),
      .r_dat       (r_dat),
      .rd_wfifo    (rd_wfifo),
      .wfifo_empty (wfifo_empty),
      .wfifo_used  (wfifo_used)
    );

  jtag_uart_scfifo_r the_jtag_uart_scfifo_r
    (
      .clk        (clk),
      .fifo_EF    (fifo_EF),
      .fifo_clear (fifo_clear),
      .fifo_rd    (fifo_rd),
      .fifo_rdata (fifo_rdata),
      .rfifo_full (rfifo_full),
      .rfifo_used (rfifo_used),
      .rst_n      (rst_n),
      .t_dat      (t_dat),
      .wr_rfifo   (wr_rfifo)
    );

  assign ipen_AE = ien_AE & fifo_AE;
  assign ipen_AF = ien_AF & (pause_irq | fifo_AF);
  assign av_irq = ipen_AE | ipen_AF;
  assign activity = t_pause | t_ena;
  always @(posedge clk or negedge rst_n)
    begin
      if (rst_n == 0)
          pause_irq <= 1'b0;
      else // only if fifo is not empty...
      if (t_pause & ~fifo_EF)
          pause_irq <= 1'b1;
      else if (read_0)
          pause_irq <= 1'b0;
    end


  always @(posedge clk or negedge rst_n)
    begin
      if (rst_n == 0)
        begin
          r_val <= 1'b0;
          t_dav <= 1'b1;
        end
      else 
        begin
          r_val <= r_ena & ~wfifo_empty;
          t_dav <= ~rfifo_full;
        end
    end


  always @(posedge clk or negedge rst_n)
    begin
      if (rst_n == 0)
        begin
          fifo_AE <= 1'b0;
          fifo_AF <= 1'b0;
          fifo_wr <= 1'b0;
          rvalid <= 1'b0;
          read_0 <= 1'b0;
          ien_AE <= 1'b0;
          ien_AF <= 1'b0;
          ac <= 1'b0;
          woverflow <= 1'b0;
          av_waitrequest <= 1'b1;
        end
      else 
        begin
          fifo_AE <= {fifo_FF,wfifo_used} <= 8;
          fifo_AF <= (7'h40 - {rfifo_full,rfifo_used}) <= 8;
          fifo_wr <= 1'b0;
          read_0 <= 1'b0;
          av_waitrequest <= ~(av_chipselect & (~av_write_n | ~av_read_n) & av_waitrequest);
          if (activity)
              ac <= 1'b1;
          // write
          if (av_chipselect & ~av_write_n & av_waitrequest)
              // addr 1 is control; addr 0 is data
              if (av_address)
                begin
                  ien_AF <= av_writedata[0];
                  ien_AE <= av_writedata[1];
                  if (av_writedata[10] & ~activity)
                      ac <= 1'b0;
                end
              else 
                begin
                  fifo_wr <= ~fifo_FF;
                  woverflow <= fifo_FF;
                end
          // read
          if (av_chipselect & ~av_read_n & av_waitrequest)
            begin
              // addr 1 is interrupt; addr 0 is data
              if (~av_address)
                  rvalid <= ~fifo_EF;
              read_0 <= ~av_address;
            end
        end
    end


  assign fifo_wdata = av_writedata[7 : 0];
  assign fifo_rd = (av_chipselect & ~av_read_n & av_waitrequest & ~av_address) ? ~fifo_EF : 1'b0;
  assign av_readdata = read_0 ? { {9{1'b0}},rfifo_full,rfifo_used,rvalid,woverflow,~fifo_FF,~fifo_EF,1'b0,ac,ipen_AE,ipen_AF,fifo_rdata } : { {9{1'b0}},(7'h40 - {fifo_FF,wfifo_used}),rvalid,woverflow,~fifo_FF,~fifo_EF,1'b0,ac,ipen_AE,ipen_AF,{6{1'b0}},ien_AE,ien_AF };
  always @(posedge clk or negedge rst_n)
    begin
      if (rst_n == 0)
          readyfordata <= 0;
      else 
        readyfordata <= ~fifo_FF;
    end



//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  // Tie off Atlantic Interface signals not used for simulation
  always @(posedge clk)
    begin
      sim_t_pause <= 1'b0;
      sim_t_ena <= 1'b0;
      sim_t_dat <= t_dav ? r_dat : {8{r_val}};
      sim_r_ena <= 1'b0;
    end


  assign r_ena = sim_r_ena;
  assign t_ena = sim_t_ena;
  assign t_dat = sim_t_dat;
  assign t_pause = sim_t_pause;
  always @(fifo_EF)
    begin
      dataavailable = ~fifo_EF;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  alt_jtag_atlantic jtag_uart_alt_jtag_atlantic
//    (
//      .clk (clk),
//      .r_dat (r_dat),
//      .r_ena (r_ena),
//      .r_val (r_val),
//      .rst_n (rst_n),
//      .t_dat (t_dat),
//      .t_dav (t_dav),
//      .t_ena (t_ena),
//      .t_pause (t_pause)
//    );
//
//  defparam jtag_uart_alt_jtag_atlantic.INSTANCE_ID = 0,
//           jtag_uart_alt_jtag_atlantic.LOG2_RXFIFO_DEPTH = 6,
//           jtag_uart_alt_jtag_atlantic.LOG2_TXFIFO_DEPTH = 6,
//           jtag_uart_alt_jtag_atlantic.SLD_AUTO_INSTANCE_INDEX = "YES";
//
//  always @(posedge clk or negedge rst_n)
//    begin
//      if (rst_n == 0)
//          dataavailable <= 0;
//      else 
//        dataavailable <= ~fifo_EF;
//    end
//
//
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20481 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_0.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: cpu/data_master
//adapter masters: ext_ssram/s1
//asp_debug: 0
//byteaddr_width: 23
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 4
//downstream_addr_shift: 2
//downstream_burstcount_width: 1
//downstream_max_burstcount: 1
//downstream_pipeline: 1
//dynamic_slave: 1
//master_always_burst_max_burst: 0
//master_burst_on_burst_boundaries_only: 1
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 0
//nativeaddr_width: 21
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 0
//upstream_burstcount: upstream_burstcount
//upstream_burstcount_width: 4
//upstream_max_burstcount: 8
//zero_address_width: 0


module custom_dma_burst_0 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_burstcount,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             reg_downstream_address,
                             reg_downstream_arbitrationshare,
                             reg_downstream_burstcount,
                             reg_downstream_byteenable,
                             reg_downstream_debugaccess,
                             reg_downstream_nativeaddress,
                             reg_downstream_read,
                             reg_downstream_write,
                             reg_downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 20: 0] reg_downstream_address;
  output  [  3: 0] reg_downstream_arbitrationshare;
  output           reg_downstream_burstcount;
  output  [  3: 0] reg_downstream_byteenable;
  output           reg_downstream_debugaccess;
  output  [ 20: 0] reg_downstream_nativeaddress;
  output           reg_downstream_read;
  output           reg_downstream_write;
  output  [ 31: 0] reg_downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 22: 0] upstream_address;
  input   [  3: 0] upstream_burstcount;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 20: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  2: 0] address_offset;
  reg              atomic_counter;
  wire    [ 22: 0] current_upstream_address;
  wire    [  3: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  3: 0] data_counter;
  wire    [  3: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 20: 0] downstream_address;
  wire    [ 22: 0] downstream_address_base;
  wire    [  3: 0] downstream_arbitrationshare;
  wire             downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 20: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire             max_burst_size;
  wire             p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  2: 0] read_address_offset;
  wire             read_update_count;
  wire    [  3: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 20: 0] reg_downstream_address;
  reg     [  3: 0] reg_downstream_arbitrationshare;
  reg              reg_downstream_burstcount;
  reg     [  3: 0] reg_downstream_byteenable;
  reg              reg_downstream_debugaccess;
  reg     [ 20: 0] reg_downstream_nativeaddress;
  reg              reg_downstream_read;
  reg              reg_downstream_write;
  reg     [ 31: 0] reg_downstream_writedata;
  reg     [  3: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 22: 0] registered_upstream_address;
  reg     [  3: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 20: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  3: 0] transactions_remaining;
  reg     [  3: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  2: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= upstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? upstream_burstcount : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 1;
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign downstream_arbitrationshare = current_upstream_read ? (dbs_adjusted_upstream_burstcount) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign downstream_address = downstream_address_base + {address_offset, 2'b00};
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_address <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_address <= downstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_arbitrationshare <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_arbitrationshare <= downstream_arbitrationshare;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_burstcount <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_burstcount <= downstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_byteenable <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_byteenable <= downstream_byteenable;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_debugaccess <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_debugaccess <= downstream_debugaccess;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_nativeaddress <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_nativeaddress <= downstream_nativeaddress;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_read <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_read <= downstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_write <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_write <= downstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_writedata <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_writedata <= downstream_writedata;
    end



endmodule


/* SLline 20482 "custom_dma.v" 2 */
/* SLline 1 "pipeline_bridge.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_downstream_adapter (
                                            // inputs:
                                             m1_clk,
                                             m1_endofpacket,
                                             m1_readdata,
                                             m1_readdatavalid,
                                             m1_reset_n,
                                             m1_waitrequest,
                                             s1_address,
                                             s1_arbiterlock,
                                             s1_arbiterlock2,
                                             s1_burstcount,
                                             s1_byteenable,
                                             s1_chipselect,
                                             s1_debugaccess,
                                             s1_nativeaddress,
                                             s1_read,
                                             s1_write,
                                             s1_writedata,

                                            // outputs:
                                             m1_address,
                                             m1_arbiterlock,
                                             m1_arbiterlock2,
                                             m1_burstcount,
                                             m1_byteenable,
                                             m1_chipselect,
                                             m1_debugaccess,
                                             m1_nativeaddress,
                                             m1_read,
                                             m1_write,
                                             m1_writedata,
                                             s1_endofpacket,
                                             s1_readdata,
                                             s1_readdatavalid,
                                             s1_waitrequest
                                          )
;

  output  [ 11: 0] m1_address;
  output           m1_arbiterlock;
  output           m1_arbiterlock2;
  output           m1_burstcount;
  output  [  3: 0] m1_byteenable;
  output           m1_chipselect;
  output           m1_debugaccess;
  output  [  9: 0] m1_nativeaddress;
  output           m1_read;
  output           m1_write;
  output  [ 31: 0] m1_writedata;
  output           s1_endofpacket;
  output  [ 31: 0] s1_readdata;
  output           s1_readdatavalid;
  output           s1_waitrequest;
  input            m1_clk;
  input            m1_endofpacket;
  input   [ 31: 0] m1_readdata;
  input            m1_readdatavalid;
  input            m1_reset_n;
  input            m1_waitrequest;
  input   [ 11: 0] s1_address;
  input            s1_arbiterlock;
  input            s1_arbiterlock2;
  input            s1_burstcount;
  input   [  3: 0] s1_byteenable;
  input            s1_chipselect;
  input            s1_debugaccess;
  input   [  9: 0] s1_nativeaddress;
  input            s1_read;
  input            s1_write;
  input   [ 31: 0] s1_writedata;

  reg     [ 11: 0] m1_address;
  reg              m1_arbiterlock;
  reg              m1_arbiterlock2;
  reg              m1_burstcount;
  reg     [  3: 0] m1_byteenable;
  reg              m1_chipselect;
  reg              m1_debugaccess;
  reg     [  9: 0] m1_nativeaddress;
  reg              m1_read;
  reg              m1_write;
  reg     [ 31: 0] m1_writedata;
  wire             s1_endofpacket;
  wire    [ 31: 0] s1_readdata;
  wire             s1_readdatavalid;
  wire             s1_waitrequest;
  //s1, which is an e_avalon_adapter_slave
  //m1, which is an e_avalon_adapter_master
  assign s1_endofpacket = m1_endofpacket;
  assign s1_readdata = m1_readdata;
  assign s1_readdatavalid = m1_readdatavalid;
  assign s1_waitrequest = m1_waitrequest;
  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_address <= 0;
      else if (~m1_waitrequest)
          m1_address <= s1_address;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_arbiterlock <= 0;
      else if (~m1_waitrequest)
          m1_arbiterlock <= s1_arbiterlock;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_arbiterlock2 <= 0;
      else if (~m1_waitrequest)
          m1_arbiterlock2 <= s1_arbiterlock2;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_burstcount <= 0;
      else if (~m1_waitrequest)
          m1_burstcount <= s1_burstcount;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_byteenable <= 0;
      else if (~m1_waitrequest)
          m1_byteenable <= s1_byteenable;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_chipselect <= 0;
      else if (~m1_waitrequest)
          m1_chipselect <= s1_chipselect;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_debugaccess <= 0;
      else if (~m1_waitrequest)
          m1_debugaccess <= s1_debugaccess;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_nativeaddress <= 0;
      else if (~m1_waitrequest)
          m1_nativeaddress <= s1_nativeaddress;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_read <= 0;
      else if (~m1_waitrequest)
          m1_read <= s1_read;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_write <= 0;
      else if (~m1_waitrequest)
          m1_write <= s1_write;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          m1_writedata <= 0;
      else if (~m1_waitrequest)
          m1_writedata <= s1_writedata;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_upstream_adapter (
                                          // inputs:
                                           m1_clk,
                                           m1_endofpacket,
                                           m1_readdata,
                                           m1_readdatavalid,
                                           m1_reset_n,
                                           m1_waitrequest,
                                           s1_address,
                                           s1_arbiterlock,
                                           s1_arbiterlock2,
                                           s1_burstcount,
                                           s1_byteenable,
                                           s1_chipselect,
                                           s1_clk,
                                           s1_debugaccess,
                                           s1_flush,
                                           s1_nativeaddress,
                                           s1_read,
                                           s1_reset_n,
                                           s1_write,
                                           s1_writedata,

                                          // outputs:
                                           m1_address,
                                           m1_arbiterlock,
                                           m1_arbiterlock2,
                                           m1_burstcount,
                                           m1_byteenable,
                                           m1_chipselect,
                                           m1_debugaccess,
                                           m1_nativeaddress,
                                           m1_read,
                                           m1_write,
                                           m1_writedata,
                                           s1_endofpacket,
                                           s1_readdata,
                                           s1_readdatavalid,
                                           s1_waitrequest
                                        )
;

  output  [ 11: 0] m1_address;
  output           m1_arbiterlock;
  output           m1_arbiterlock2;
  output           m1_burstcount;
  output  [  3: 0] m1_byteenable;
  output           m1_chipselect;
  output           m1_debugaccess;
  output  [  9: 0] m1_nativeaddress;
  output           m1_read;
  output           m1_write;
  output  [ 31: 0] m1_writedata;
  output           s1_endofpacket;
  output  [ 31: 0] s1_readdata;
  output           s1_readdatavalid;
  output           s1_waitrequest;
  input            m1_clk;
  input            m1_endofpacket;
  input   [ 31: 0] m1_readdata;
  input            m1_readdatavalid;
  input            m1_reset_n;
  input            m1_waitrequest;
  input   [ 11: 0] s1_address;
  input            s1_arbiterlock;
  input            s1_arbiterlock2;
  input            s1_burstcount;
  input   [  3: 0] s1_byteenable;
  input            s1_chipselect;
  input            s1_clk;
  input            s1_debugaccess;
  input            s1_flush;
  input   [  9: 0] s1_nativeaddress;
  input            s1_read;
  input            s1_reset_n;
  input            s1_write;
  input   [ 31: 0] s1_writedata;

  wire    [ 11: 0] m1_address;
  wire             m1_arbiterlock;
  wire             m1_arbiterlock2;
  wire             m1_burstcount;
  wire    [  3: 0] m1_byteenable;
  wire             m1_chipselect;
  wire             m1_debugaccess;
  wire    [  9: 0] m1_nativeaddress;
  wire             m1_read;
  wire             m1_write;
  wire    [ 31: 0] m1_writedata;
  reg              s1_endofpacket;
  reg     [ 31: 0] s1_readdata;
  reg              s1_readdatavalid;
  wire             s1_waitrequest;
  //s1, which is an e_avalon_adapter_slave
  //m1, which is an e_avalon_adapter_master
  always @(posedge s1_clk or negedge s1_reset_n)
    begin
      if (s1_reset_n == 0)
          s1_readdatavalid <= 0;
      else if (s1_flush)
          s1_readdatavalid <= 0;
      else 
        s1_readdatavalid <= m1_readdatavalid;
    end


  assign s1_waitrequest = m1_waitrequest;
  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          s1_endofpacket <= 0;
      else if (m1_readdatavalid)
          s1_endofpacket <= m1_endofpacket;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          s1_readdata <= 0;
      else if (m1_readdatavalid)
          s1_readdata <= m1_readdata;
    end


  assign m1_address = s1_address;
  assign m1_arbiterlock = s1_arbiterlock;
  assign m1_arbiterlock2 = s1_arbiterlock2;
  assign m1_burstcount = s1_burstcount;
  assign m1_byteenable = s1_byteenable;
  assign m1_chipselect = s1_chipselect;
  assign m1_debugaccess = s1_debugaccess;
  assign m1_nativeaddress = s1_nativeaddress;
  assign m1_read = s1_read;
  assign m1_write = s1_write;
  assign m1_writedata = s1_writedata;

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge_waitrequest_adapter (
                                             // inputs:
                                              m1_clk,
                                              m1_endofpacket,
                                              m1_readdata,
                                              m1_readdatavalid,
                                              m1_reset_n,
                                              m1_waitrequest,
                                              reset_n,
                                              s1_address,
                                              s1_arbiterlock,
                                              s1_arbiterlock2,
                                              s1_burstcount,
                                              s1_byteenable,
                                              s1_chipselect,
                                              s1_debugaccess,
                                              s1_nativeaddress,
                                              s1_read,
                                              s1_write,
                                              s1_writedata,

                                             // outputs:
                                              m1_address,
                                              m1_arbiterlock,
                                              m1_arbiterlock2,
                                              m1_burstcount,
                                              m1_byteenable,
                                              m1_chipselect,
                                              m1_debugaccess,
                                              m1_nativeaddress,
                                              m1_read,
                                              m1_write,
                                              m1_writedata,
                                              s1_endofpacket,
                                              s1_readdata,
                                              s1_readdatavalid,
                                              s1_waitrequest
                                           )
;

  output  [ 11: 0] m1_address;
  output           m1_arbiterlock;
  output           m1_arbiterlock2;
  output           m1_burstcount;
  output  [  3: 0] m1_byteenable;
  output           m1_chipselect;
  output           m1_debugaccess;
  output  [  9: 0] m1_nativeaddress;
  output           m1_read;
  output           m1_write;
  output  [ 31: 0] m1_writedata;
  output           s1_endofpacket;
  output  [ 31: 0] s1_readdata;
  output           s1_readdatavalid;
  output           s1_waitrequest;
  input            m1_clk;
  input            m1_endofpacket;
  input   [ 31: 0] m1_readdata;
  input            m1_readdatavalid;
  input            m1_reset_n;
  input            m1_waitrequest;
  input            reset_n;
  input   [ 11: 0] s1_address;
  input            s1_arbiterlock;
  input            s1_arbiterlock2;
  input            s1_burstcount;
  input   [  3: 0] s1_byteenable;
  input            s1_chipselect;
  input            s1_debugaccess;
  input   [  9: 0] s1_nativeaddress;
  input            s1_read;
  input            s1_write;
  input   [ 31: 0] s1_writedata;

  reg     [ 11: 0] d1_s1_address;
  reg              d1_s1_arbiterlock;
  reg              d1_s1_arbiterlock2;
  reg              d1_s1_burstcount;
  reg     [  3: 0] d1_s1_byteenable;
  reg              d1_s1_chipselect;
  reg              d1_s1_debugaccess;
  reg     [  9: 0] d1_s1_nativeaddress;
  reg              d1_s1_read;
  reg              d1_s1_write;
  reg     [ 31: 0] d1_s1_writedata;
  wire    [ 11: 0] m1_address;
  wire             m1_arbiterlock;
  wire             m1_arbiterlock2;
  wire             m1_burstcount;
  wire    [  3: 0] m1_byteenable;
  wire             m1_chipselect;
  wire             m1_debugaccess;
  wire    [  9: 0] m1_nativeaddress;
  wire             m1_read;
  wire             m1_write;
  wire    [ 31: 0] m1_writedata;
  wire             s1_endofpacket;
  wire    [ 31: 0] s1_readdata;
  wire             s1_readdatavalid;
  reg              s1_waitrequest;
  wire             set_use_registered;
  reg              use_registered;
  //s1, which is an e_avalon_adapter_slave
  //m1, which is an e_avalon_adapter_master
  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          s1_waitrequest <= 0;
      else 
        s1_waitrequest <= m1_waitrequest;
    end


  assign s1_endofpacket = m1_endofpacket;
  assign s1_readdata = m1_readdata;
  assign s1_readdatavalid = m1_readdatavalid;
  //set use registered, which is an e_assign
  assign set_use_registered = m1_waitrequest & ~s1_waitrequest;

  //use registered, which is an e_register
  always @(posedge m1_clk or negedge reset_n)
    begin
      if (reset_n == 0)
          use_registered <= 0;
      else if (~m1_waitrequest & s1_waitrequest)
          use_registered <= 0;
      else if (set_use_registered)
          use_registered <= -1;
    end


  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_address <= 0;
      else if (set_use_registered)
          d1_s1_address <= s1_address;
    end


  assign m1_address = (use_registered)? d1_s1_address :
    s1_address;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_arbiterlock <= 0;
      else if (set_use_registered)
          d1_s1_arbiterlock <= s1_arbiterlock;
    end


  assign m1_arbiterlock = (use_registered)? d1_s1_arbiterlock :
    s1_arbiterlock;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_arbiterlock2 <= 0;
      else if (set_use_registered)
          d1_s1_arbiterlock2 <= s1_arbiterlock2;
    end


  assign m1_arbiterlock2 = (use_registered)? d1_s1_arbiterlock2 :
    s1_arbiterlock2;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_burstcount <= 0;
      else if (set_use_registered)
          d1_s1_burstcount <= s1_burstcount;
    end


  assign m1_burstcount = (use_registered)? d1_s1_burstcount :
    s1_burstcount;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_byteenable <= 0;
      else if (set_use_registered)
          d1_s1_byteenable <= s1_byteenable;
    end


  assign m1_byteenable = (use_registered)? d1_s1_byteenable :
    s1_byteenable;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_chipselect <= 0;
      else if (set_use_registered)
          d1_s1_chipselect <= s1_chipselect;
    end


  assign m1_chipselect = (use_registered)? d1_s1_chipselect :
    s1_chipselect;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_debugaccess <= 0;
      else if (set_use_registered)
          d1_s1_debugaccess <= s1_debugaccess;
    end


  assign m1_debugaccess = (use_registered)? d1_s1_debugaccess :
    s1_debugaccess;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_nativeaddress <= 0;
      else if (set_use_registered)
          d1_s1_nativeaddress <= s1_nativeaddress;
    end


  assign m1_nativeaddress = (use_registered)? d1_s1_nativeaddress :
    s1_nativeaddress;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_read <= 0;
      else if (set_use_registered)
          d1_s1_read <= s1_read;
    end


  assign m1_read = (use_registered)? d1_s1_read :
    s1_read;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_write <= 0;
      else if (set_use_registered)
          d1_s1_write <= s1_write;
    end


  assign m1_write = (use_registered)? d1_s1_write :
    s1_write;

  always @(posedge m1_clk or negedge m1_reset_n)
    begin
      if (m1_reset_n == 0)
          d1_s1_writedata <= 0;
      else if (set_use_registered)
          d1_s1_writedata <= s1_writedata;
    end


  assign m1_writedata = (use_registered)? d1_s1_writedata :
    s1_writedata;


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module pipeline_bridge (
                         // inputs:
                          clk,
                          m1_endofpacket,
                          m1_readdata,
                          m1_readdatavalid,
                          m1_waitrequest,
                          reset_n,
                          s1_address,
                          s1_arbiterlock,
                          s1_arbiterlock2,
                          s1_burstcount,
                          s1_byteenable,
                          s1_chipselect,
                          s1_debugaccess,
                          s1_nativeaddress,
                          s1_read,
                          s1_write,
                          s1_writedata,

                         // outputs:
                          m1_address,
                          m1_burstcount,
                          m1_byteenable,
                          m1_chipselect,
                          m1_debugaccess,
                          m1_read,
                          m1_write,
                          m1_writedata,
                          s1_endofpacket,
                          s1_readdata,
                          s1_readdatavalid,
                          s1_waitrequest
                       )
;

  output  [ 11: 0] m1_address;
  output           m1_burstcount;
  output  [  3: 0] m1_byteenable;
  output           m1_chipselect;
  output           m1_debugaccess;
  output           m1_read;
  output           m1_write;
  output  [ 31: 0] m1_writedata;
  output           s1_endofpacket;
  output  [ 31: 0] s1_readdata;
  output           s1_readdatavalid;
  output           s1_waitrequest;
  input            clk;
  input            m1_endofpacket;
  input   [ 31: 0] m1_readdata;
  input            m1_readdatavalid;
  input            m1_waitrequest;
  input            reset_n;
  input   [  9: 0] s1_address;
  input            s1_arbiterlock;
  input            s1_arbiterlock2;
  input            s1_burstcount;
  input   [  3: 0] s1_byteenable;
  input            s1_chipselect;
  input            s1_debugaccess;
  input   [  9: 0] s1_nativeaddress;
  input            s1_read;
  input            s1_write;
  input   [ 31: 0] s1_writedata;

  wire    [ 11: 0] downstream_m1_address;
  wire             downstream_m1_arbiterlock;
  wire             downstream_m1_arbiterlock2;
  wire             downstream_m1_burstcount;
  wire    [  3: 0] downstream_m1_byteenable;
  wire             downstream_m1_chipselect;
  wire             downstream_m1_debugaccess;
  wire             downstream_m1_endofpacket;
  wire    [  9: 0] downstream_m1_nativeaddress;
  wire             downstream_m1_read;
  wire    [ 31: 0] downstream_m1_readdata;
  wire             downstream_m1_readdatavalid;
  wire             downstream_m1_waitrequest;
  wire             downstream_m1_write;
  wire    [ 31: 0] downstream_m1_writedata;
  wire    [ 11: 0] downstream_s1_address;
  wire             downstream_s1_arbiterlock;
  wire             downstream_s1_arbiterlock2;
  wire             downstream_s1_burstcount;
  wire    [  3: 0] downstream_s1_byteenable;
  wire             downstream_s1_chipselect;
  wire             downstream_s1_debugaccess;
  wire             downstream_s1_endofpacket;
  wire    [  9: 0] downstream_s1_nativeaddress;
  wire             downstream_s1_read;
  wire    [ 31: 0] downstream_s1_readdata;
  wire             downstream_s1_readdatavalid;
  wire             downstream_s1_waitrequest;
  wire             downstream_s1_write;
  wire    [ 31: 0] downstream_s1_writedata;
  wire    [ 11: 0] m1_address;
  wire             m1_arbiterlock;
  wire             m1_arbiterlock2;
  wire             m1_burstcount;
  wire    [  3: 0] m1_byteenable;
  wire             m1_chipselect;
  wire             m1_debugaccess;
  wire    [  9: 0] m1_nativeaddress;
  wire             m1_read;
  wire             m1_write;
  wire    [ 31: 0] m1_writedata;
  wire             s1_endofpacket;
  wire    [ 31: 0] s1_readdata;
  wire             s1_readdatavalid;
  wire             s1_waitrequest;
  wire    [ 11: 0] upstream_m1_address;
  wire             upstream_m1_arbiterlock;
  wire             upstream_m1_arbiterlock2;
  wire             upstream_m1_burstcount;
  wire    [  3: 0] upstream_m1_byteenable;
  wire             upstream_m1_chipselect;
  wire             upstream_m1_debugaccess;
  wire             upstream_m1_endofpacket;
  wire    [  9: 0] upstream_m1_nativeaddress;
  wire             upstream_m1_read;
  wire    [ 31: 0] upstream_m1_readdata;
  wire             upstream_m1_readdatavalid;
  wire             upstream_m1_waitrequest;
  wire             upstream_m1_write;
  wire    [ 31: 0] upstream_m1_writedata;
  wire    [ 11: 0] upstream_s1_address;
  wire             upstream_s1_arbiterlock;
  wire             upstream_s1_arbiterlock2;
  wire             upstream_s1_burstcount;
  wire    [  3: 0] upstream_s1_byteenable;
  wire             upstream_s1_chipselect;
  wire             upstream_s1_debugaccess;
  wire             upstream_s1_endofpacket;
  wire    [  9: 0] upstream_s1_nativeaddress;
  wire             upstream_s1_read;
  wire    [ 31: 0] upstream_s1_readdata;
  wire             upstream_s1_readdatavalid;
  wire             upstream_s1_waitrequest;
  wire             upstream_s1_write;
  wire    [ 31: 0] upstream_s1_writedata;
  wire    [ 11: 0] waitrequest_m1_address;
  wire             waitrequest_m1_arbiterlock;
  wire             waitrequest_m1_arbiterlock2;
  wire             waitrequest_m1_burstcount;
  wire    [  3: 0] waitrequest_m1_byteenable;
  wire             waitrequest_m1_chipselect;
  wire             waitrequest_m1_debugaccess;
  wire             waitrequest_m1_endofpacket;
  wire    [  9: 0] waitrequest_m1_nativeaddress;
  wire             waitrequest_m1_read;
  wire    [ 31: 0] waitrequest_m1_readdata;
  wire             waitrequest_m1_readdatavalid;
  wire             waitrequest_m1_waitrequest;
  wire             waitrequest_m1_write;
  wire    [ 31: 0] waitrequest_m1_writedata;
  wire    [ 11: 0] waitrequest_s1_address;
  wire             waitrequest_s1_arbiterlock;
  wire             waitrequest_s1_arbiterlock2;
  wire             waitrequest_s1_burstcount;
  wire    [  3: 0] waitrequest_s1_byteenable;
  wire             waitrequest_s1_chipselect;
  wire             waitrequest_s1_debugaccess;
  wire             waitrequest_s1_endofpacket;
  wire    [  9: 0] waitrequest_s1_nativeaddress;
  wire             waitrequest_s1_read;
  wire    [ 31: 0] waitrequest_s1_readdata;
  wire             waitrequest_s1_readdatavalid;
  wire             waitrequest_s1_waitrequest;
  wire             waitrequest_s1_write;
  wire    [ 31: 0] waitrequest_s1_writedata;
  pipeline_bridge_downstream_adapter the_pipeline_bridge_downstream_adapter
    (
      .m1_address       (downstream_m1_address),
      .m1_arbiterlock   (downstream_m1_arbiterlock),
      .m1_arbiterlock2  (downstream_m1_arbiterlock2),
      .m1_burstcount    (downstream_m1_burstcount),
      .m1_byteenable    (downstream_m1_byteenable),
      .m1_chipselect    (downstream_m1_chipselect),
      .m1_clk           (clk),
      .m1_debugaccess   (downstream_m1_debugaccess),
      .m1_endofpacket   (downstream_m1_endofpacket),
      .m1_nativeaddress (downstream_m1_nativeaddress),
      .m1_read          (downstream_m1_read),
      .m1_readdata      (downstream_m1_readdata),
      .m1_readdatavalid (downstream_m1_readdatavalid),
      .m1_reset_n       (reset_n),
      .m1_waitrequest   (downstream_m1_waitrequest),
      .m1_write         (downstream_m1_write),
      .m1_writedata     (downstream_m1_writedata),
      .s1_address       (downstream_s1_address),
      .s1_arbiterlock   (downstream_s1_arbiterlock),
      .s1_arbiterlock2  (downstream_s1_arbiterlock2),
      .s1_burstcount    (downstream_s1_burstcount),
      .s1_byteenable    (downstream_s1_byteenable),
      .s1_chipselect    (downstream_s1_chipselect),
      .s1_debugaccess   (downstream_s1_debugaccess),
      .s1_endofpacket   (downstream_s1_endofpacket),
      .s1_nativeaddress (downstream_s1_nativeaddress),
      .s1_read          (downstream_s1_read),
      .s1_readdata      (downstream_s1_readdata),
      .s1_readdatavalid (downstream_s1_readdatavalid),
      .s1_waitrequest   (downstream_s1_waitrequest),
      .s1_write         (downstream_s1_write),
      .s1_writedata     (downstream_s1_writedata)
    );

  pipeline_bridge_upstream_adapter the_pipeline_bridge_upstream_adapter
    (
      .m1_address       (upstream_m1_address),
      .m1_arbiterlock   (upstream_m1_arbiterlock),
      .m1_arbiterlock2  (upstream_m1_arbiterlock2),
      .m1_burstcount    (upstream_m1_burstcount),
      .m1_byteenable    (upstream_m1_byteenable),
      .m1_chipselect    (upstream_m1_chipselect),
      .m1_clk           (clk),
      .m1_debugaccess   (upstream_m1_debugaccess),
      .m1_endofpacket   (upstream_m1_endofpacket),
      .m1_nativeaddress (upstream_m1_nativeaddress),
      .m1_read          (upstream_m1_read),
      .m1_readdata      (upstream_m1_readdata),
      .m1_readdatavalid (upstream_m1_readdatavalid),
      .m1_reset_n       (reset_n),
      .m1_waitrequest   (upstream_m1_waitrequest),
      .m1_write         (upstream_m1_write),
      .m1_writedata     (upstream_m1_writedata),
      .s1_address       (upstream_s1_address),
      .s1_arbiterlock   (upstream_s1_arbiterlock),
      .s1_arbiterlock2  (upstream_s1_arbiterlock2),
      .s1_burstcount    (upstream_s1_burstcount),
      .s1_byteenable    (upstream_s1_byteenable),
      .s1_chipselect    (upstream_s1_chipselect),
      .s1_clk           (clk),
      .s1_debugaccess   (upstream_s1_debugaccess),
      .s1_endofpacket   (upstream_s1_endofpacket),
      .s1_flush         (1'b0),
      .s1_nativeaddress (upstream_s1_nativeaddress),
      .s1_read          (upstream_s1_read),
      .s1_readdata      (upstream_s1_readdata),
      .s1_readdatavalid (upstream_s1_readdatavalid),
      .s1_reset_n       (reset_n),
      .s1_waitrequest   (upstream_s1_waitrequest),
      .s1_write         (upstream_s1_write),
      .s1_writedata     (upstream_s1_writedata)
    );

  pipeline_bridge_waitrequest_adapter the_pipeline_bridge_waitrequest_adapter
    (
      .m1_address       (waitrequest_m1_address),
      .m1_arbiterlock   (waitrequest_m1_arbiterlock),
      .m1_arbiterlock2  (waitrequest_m1_arbiterlock2),
      .m1_burstcount    (waitrequest_m1_burstcount),
      .m1_byteenable    (waitrequest_m1_byteenable),
      .m1_chipselect    (waitrequest_m1_chipselect),
      .m1_clk           (clk),
      .m1_debugaccess   (waitrequest_m1_debugaccess),
      .m1_endofpacket   (waitrequest_m1_endofpacket),
      .m1_nativeaddress (waitrequest_m1_nativeaddress),
      .m1_read          (waitrequest_m1_read),
      .m1_readdata      (waitrequest_m1_readdata),
      .m1_readdatavalid (waitrequest_m1_readdatavalid),
      .m1_reset_n       (reset_n),
      .m1_waitrequest   (waitrequest_m1_waitrequest),
      .m1_write         (waitrequest_m1_write),
      .m1_writedata     (waitrequest_m1_writedata),
      .reset_n          (reset_n),
      .s1_address       (waitrequest_s1_address),
      .s1_arbiterlock   (waitrequest_s1_arbiterlock),
      .s1_arbiterlock2  (waitrequest_s1_arbiterlock2),
      .s1_burstcount    (waitrequest_s1_burstcount),
      .s1_byteenable    (waitrequest_s1_byteenable),
      .s1_chipselect    (waitrequest_s1_chipselect),
      .s1_debugaccess   (waitrequest_s1_debugaccess),
      .s1_endofpacket   (waitrequest_s1_endofpacket),
      .s1_nativeaddress (waitrequest_s1_nativeaddress),
      .s1_read          (waitrequest_s1_read),
      .s1_readdata      (waitrequest_s1_readdata),
      .s1_readdatavalid (waitrequest_s1_readdatavalid),
      .s1_waitrequest   (waitrequest_s1_waitrequest),
      .s1_write         (waitrequest_s1_write),
      .s1_writedata     (waitrequest_s1_writedata)
    );

  assign m1_nativeaddress = downstream_m1_nativeaddress;
  assign downstream_s1_nativeaddress = upstream_m1_nativeaddress;
  assign upstream_s1_nativeaddress = waitrequest_m1_nativeaddress;
  assign waitrequest_s1_nativeaddress = s1_nativeaddress;
  assign m1_debugaccess = downstream_m1_debugaccess;
  assign downstream_s1_debugaccess = upstream_m1_debugaccess;
  assign upstream_s1_debugaccess = waitrequest_m1_debugaccess;
  assign waitrequest_s1_debugaccess = s1_debugaccess;
  assign m1_arbiterlock = downstream_m1_arbiterlock;
  assign downstream_s1_arbiterlock = upstream_m1_arbiterlock;
  assign upstream_s1_arbiterlock = waitrequest_m1_arbiterlock;
  assign waitrequest_s1_arbiterlock = s1_arbiterlock;
  assign m1_writedata = downstream_m1_writedata;
  assign downstream_s1_writedata = upstream_m1_writedata;
  assign upstream_s1_writedata = waitrequest_m1_writedata;
  assign waitrequest_s1_writedata = s1_writedata;
  assign m1_chipselect = downstream_m1_chipselect;
  assign downstream_s1_chipselect = upstream_m1_chipselect;
  assign upstream_s1_chipselect = waitrequest_m1_chipselect;
  assign waitrequest_s1_chipselect = s1_chipselect;
  assign m1_burstcount = downstream_m1_burstcount;
  assign downstream_s1_burstcount = upstream_m1_burstcount;
  assign upstream_s1_burstcount = waitrequest_m1_burstcount;
  assign waitrequest_s1_burstcount = s1_burstcount;
  assign m1_byteenable = downstream_m1_byteenable;
  assign downstream_s1_byteenable = upstream_m1_byteenable;
  assign upstream_s1_byteenable = waitrequest_m1_byteenable;
  assign waitrequest_s1_byteenable = s1_byteenable;
  assign m1_arbiterlock2 = downstream_m1_arbiterlock2;
  assign downstream_s1_arbiterlock2 = upstream_m1_arbiterlock2;
  assign upstream_s1_arbiterlock2 = waitrequest_m1_arbiterlock2;
  assign waitrequest_s1_arbiterlock2 = s1_arbiterlock2;
  assign m1_read = downstream_m1_read;
  assign downstream_s1_read = upstream_m1_read;
  assign upstream_s1_read = waitrequest_m1_read;
  assign waitrequest_s1_read = s1_read;
  assign m1_write = downstream_m1_write;
  assign downstream_s1_write = upstream_m1_write;
  assign upstream_s1_write = waitrequest_m1_write;
  assign waitrequest_s1_write = s1_write;
  assign waitrequest_s1_address = {s1_address, 2'b0};
  assign upstream_s1_address = waitrequest_m1_address;
  assign downstream_s1_address = upstream_m1_address;
  assign m1_address = downstream_m1_address;
  assign downstream_m1_readdatavalid = m1_readdatavalid;
  assign upstream_m1_readdatavalid = downstream_s1_readdatavalid;
  assign waitrequest_m1_readdatavalid = upstream_s1_readdatavalid;
  assign s1_readdatavalid = waitrequest_s1_readdatavalid;
  assign downstream_m1_waitrequest = m1_waitrequest;
  assign upstream_m1_waitrequest = downstream_s1_waitrequest;
  assign waitrequest_m1_waitrequest = upstream_s1_waitrequest;
  assign s1_waitrequest = waitrequest_s1_waitrequest;
  assign downstream_m1_endofpacket = m1_endofpacket;
  assign upstream_m1_endofpacket = downstream_s1_endofpacket;
  assign waitrequest_m1_endofpacket = upstream_s1_endofpacket;
  assign s1_endofpacket = waitrequest_s1_endofpacket;
  assign downstream_m1_readdata = m1_readdata;
  assign upstream_m1_readdata = downstream_s1_readdata;
  assign waitrequest_m1_readdata = upstream_s1_readdata;
  assign s1_readdata = waitrequest_s1_readdata;
  //s1, which is an e_avalon_slave
  //m1, which is an e_avalon_master

endmodule


/* SLline 20483 "custom_dma.v" 2 */
/* SLline 1 "ddr_sdram_test_component.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_test_component_ram_module (
                                             // inputs:
                                              data,
                                              rdaddress,
                                              rdclken,
                                              wraddress,
                                              wrclock,
                                              wren,

                                             // outputs:
                                              q
                                           )
;

  output  [ 31: 0] q;
  input   [ 31: 0] data;
  input   [ 23: 0] rdaddress;
  input            rdclken;
  input   [ 23: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [ 31: 0] mem_array [16777215: 0];
  wire    [ 31: 0] q;
  reg     [ 23: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("ddr_sdram.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "UNUSED",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 32,
//           lpm_ram_dp_component.lpm_widthad = 24,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module ddr_sdram_test_component (
                                  // inputs:
                                   clk,
                                   ddr_a,
                                   ddr_ba,
                                   ddr_cas_n,
                                   ddr_cke,
                                   ddr_cs_n,
                                   ddr_dm,
                                   ddr_ras_n,
                                   ddr_we_n,

                                  // outputs:
                                   ddr_dq,
                                   ddr_dqs
                                )
;

  inout   [ 15: 0] ddr_dq;
  inout   [  1: 0] ddr_dqs;
  input            clk;
  input   [ 12: 0] ddr_a;
  input   [  1: 0] ddr_ba;
  input            ddr_cas_n;
  input            ddr_cke;
  input            ddr_cs_n;
  input   [  1: 0] ddr_dm;
  input            ddr_ras_n;
  input            ddr_we_n;

  wire    [ 23: 0] CODE;
  wire    [ 12: 0] a;
  wire    [  7: 0] addr_col;
  wire    [  1: 0] ba;
  reg     [  2: 0] burstlength;
  reg              burstmode;
  reg              cas2;
  reg              cas25;
  reg              cas3;
  wire             cas_n;
  wire             cke;
  wire    [  2: 0] cmd_code;
  wire             cs_n;
  wire    [  2: 0] current_row;
  wire    [ 15: 0] ddr_dq;
  wire    [  1: 0] ddr_dqs;
  wire    [  1: 0] dm;
  reg     [  3: 0] dm_captured;
  reg     [ 31: 0] dq_captured;
  wire    [ 15: 0] dq_out_0;
  wire    [ 15: 0] dq_temp;
  wire             dq_valid;
  wire    [  1: 0] dqs_out_0;
  wire    [  1: 0] dqs_temp;
  wire             dqs_valid;
  reg              dqs_valid_temp;
  reg     [ 15: 0] first_half_dq;
  reg     [  2: 0] index;
  wire    [ 31: 0] mem_bytes;
  reg     [ 12: 0] open_rows [  7: 0];
  wire             ras_n;
  reg     [ 23: 0] rd_addr_pipe_0;
  reg     [ 23: 0] rd_addr_pipe_1;
  reg     [ 23: 0] rd_addr_pipe_2;
  reg     [ 23: 0] rd_addr_pipe_3;
  reg     [ 23: 0] rd_addr_pipe_4;
  reg     [ 23: 0] rd_addr_pipe_5;
  reg     [ 23: 0] rd_burst_counter;
  reg     [  5: 0] rd_valid_pipe;
  wire    [ 23: 0] read_addr_delayed;
  reg              read_cmd;
  wire    [ 31: 0] read_data;
  wire    [ 15: 0] read_dq;
  wire             read_valid;
  reg              read_valid_r;
  reg              read_valid_r2;
  reg              read_valid_r3;
  reg              read_valid_r4;
  wire    [ 23: 0] rmw_address;
  reg     [ 31: 0] rmw_temp;
  reg     [ 15: 0] second_half_dq;
  wire    [ 23: 0] txt_code;
  wire             we_n;
  wire    [ 23: 0] wr_addr_delayed;
  reg     [ 23: 0] wr_addr_pipe_0;
  reg     [ 23: 0] wr_addr_pipe_1;
  reg     [ 23: 0] wr_addr_pipe_2;
  reg     [ 23: 0] wr_addr_pipe_3;
  reg     [ 23: 0] wr_burst_counter;
  reg              write_cmd;
  wire             write_to_ram;
  reg              write_to_ram_r;
  reg              write_valid;
  reg              write_valid_r;
  reg              write_valid_r2;
  reg              write_valid_r3;
initial
  begin
    $write("\n");
    $write("**********************************************************************\n");
    $write("This testbench includes an SOPC Builder generated Altera memory model:\n");
    $write("'ddr_sdram_test_component.v', to simulate accesses to the DDR SDRAM memory.\n");
    $write(" \n");
    $write("Initial contents are loaded from the file: 'ddr_sdram.dat'.\n");
    $write("**********************************************************************\n");
  end
  //Synchronous write when (CODE == 24'h205752 (write))
  ddr_sdram_test_component_ram_module ddr_sdram_test_component_ram
    (
      .data      (rmw_temp),
      .q         (read_data),
      .rdaddress (rmw_address),
      .rdclken   (1'b1),
      .wraddress (wr_addr_delayed),
      .wrclock   (clk),
      .wren      (write_to_ram_r)
    );

  assign cke = ddr_cke;
  assign cs_n = ddr_cs_n;
  assign ras_n = ddr_ras_n;
  assign cas_n = ddr_cas_n;
  assign we_n = ddr_we_n;
  assign dm = ddr_dm;
  assign ba = ddr_ba;
  assign a = ddr_a;
  assign cmd_code = {ras_n, cas_n, we_n};
  assign CODE = (&cs_n) ? 24'h494e48 : txt_code;
  assign addr_col = a[8 : 1];
  assign current_row = {cs_n,ba};
  // Decode commands into their actions
  always @(posedge clk)
    begin
      // No Activity if the clock is
      if (cke)
        begin
          // This is a read command
          if (cmd_code == 3'b101)
              read_cmd <= 1'b1;
          else 
            read_cmd <= 1'b0;
          // This is a write command
          if (cmd_code == 3'b100)
              write_cmd <= 1'b1;
          else 
            write_cmd <= 1'b0;
          // This is an activate - store the chip/row/bank address in the same order as the DDR controller
          if (cmd_code == 3'b011)
              open_rows[current_row] <= a;
          //Load mode register - set CAS latency, burst mode and length
          if (cmd_code == 3'b000 && ba == 2'b00)
            begin
              burstmode <= a[3];
              burstlength <= a[2 : 0] << 1;
              //Decode CAS Latency from bits a[6..4]
              if (a[6 : 4] == 3'b010)
                begin
                  cas2 <= 1'b1;
                  index <= 3'b001;
                end
              else //CAS Latency = 2.5 
              if (a[6 : 4] == 3'b110)
                begin
                  cas25 <= 1'b1;
                  index <= 3'b001;
                end
              else 
                begin
                  cas3 <= 1'b1;
                  index <= 3'b010;
                end
            end
          rd_valid_pipe[5 : 1] <= rd_valid_pipe[4 : 0];
          rd_addr_pipe_5 <= rd_addr_pipe_4;
          rd_addr_pipe_4 <= rd_addr_pipe_3;
          rd_addr_pipe_3 <= rd_addr_pipe_2;
          rd_addr_pipe_2 <= rd_addr_pipe_1;
          rd_addr_pipe_1 <= rd_addr_pipe_0;
          rd_valid_pipe[0] <= cmd_code == 3'b101;
          wr_addr_pipe_3 <= wr_addr_pipe_2;
          wr_addr_pipe_2 <= wr_addr_pipe_1;
          wr_addr_pipe_1 <= wr_addr_pipe_0;
        end
    end


  // Burst support - make the wr_addr & rd_addr keep counting
  always @(posedge clk)
    begin
      // Reset write address otherwise if the first write is partial it breaks!
      if (cmd_code == 3'b000 && ba == 2'b00)
        begin
          wr_addr_pipe_0 <= 0;
          wr_burst_counter <= 0;
        end
      else if (cmd_code == 3'b100)
        begin
          wr_addr_pipe_0 <= {ba,open_rows[current_row],addr_col};
          wr_burst_counter[23 : 2] <= {ba,open_rows[current_row],addr_col[7 : 2]};
          wr_burst_counter[1 : 0] <= addr_col[1 : 0] + 1;
        end
      else if (write_cmd || write_to_ram)
        begin
          wr_addr_pipe_0 <= wr_burst_counter;
          wr_burst_counter[1 : 0] <= wr_burst_counter[1 : 0] + 1;
        end
      else 
        wr_addr_pipe_0 <= 0;
      // Reset read address otherwise if the first write is partial it breaks!
      if (cmd_code == 3'b000 && ba == 2'b00)
          rd_addr_pipe_0 <= 0;
      else if (cmd_code == 3'b101)
        begin
          rd_addr_pipe_0 <= {ba,open_rows[current_row],addr_col};
          rd_burst_counter[23 : 2] <= {ba,open_rows[current_row],addr_col[7 : 2]};
          rd_burst_counter[1 : 0] <= addr_col[1 : 0] + 1;
        end
      else if (read_cmd || dq_valid || read_valid)
        begin
          rd_addr_pipe_0 <= rd_burst_counter;
          rd_burst_counter[1 : 0] <= rd_burst_counter[1 : 0] + 1;
        end
      else 
        rd_addr_pipe_0 <= 0;
    end


  // read data transition from single to double clock rate
  always @(posedge clk)
    begin
      first_half_dq <= read_data[31 : 16];
      second_half_dq <= read_data[15 : 0];
    end


  assign read_dq = clk  ? second_half_dq : first_half_dq;
  assign dqs_temp = dqs_valid ? {2{clk}} : {2{1'bz}};
  assign dq_temp = dq_valid  ? read_dq : {16{1'bz}};
  assign #2.5 dqs_out_0 = dqs_temp;
  assign #2.5 dq_out_0 = dq_temp;
  assign #2.5 ddr_dqs = dqs_out_0;
  assign #2.5 ddr_dq = dq_out_0;
  //Pipelining registers for burst counting
  always @(posedge clk)
    begin
      write_valid <= write_cmd;
      write_valid_r <= write_valid;
      read_valid_r <= read_valid;
      write_valid_r2 <= write_valid_r;
      write_valid_r3 <= write_valid_r2;
      write_to_ram_r <= write_to_ram;
      read_valid_r2 <= read_valid_r;
      read_valid_r3 <= read_valid_r2;
      read_valid_r4 <= read_valid_r3;
    end


  assign write_to_ram = write_valid || write_valid_r || write_valid_r2 || write_valid_r3;
  assign dq_valid = read_valid_r || read_valid_r2 || read_valid_r3 || read_valid_r4;
  assign dqs_valid = dq_valid || dqs_valid_temp;
  // 
  always @(negedge clk)
    begin
      dqs_valid_temp <= read_valid;
    end


  //capture first half of write data with rising edge of DQS, for simulation use only 1 DQS pin
  always @(posedge ddr_dqs[0])
    begin
      dq_captured[15 : 0] <= ddr_dq[15 : 0];
      dm_captured[1 : 0] <= ddr_dm[1 : 0];
    end


  //capture second half of write data with falling edge of DQS, for simulation use only 1 DQS pin
  always @(negedge ddr_dqs[0])
    begin
      dq_captured[31 : 16] <= ddr_dq[15 : 0];
      dm_captured[3 : 2] <= ddr_dm[1 : 0];
    end


  //Support for incomplete writes, do a read-modify-write with mem_bytes and the write data
  always @(posedge clk)
    begin
      if (write_to_ram)
          rmw_temp[7 : 0] <= dm_captured[0] ? mem_bytes[7 : 0] : dq_captured[7 : 0];
    end


  always @(posedge clk)
    begin
      if (write_to_ram)
          rmw_temp[15 : 8] <= dm_captured[1] ? mem_bytes[15 : 8] : dq_captured[15 : 8];
    end


  always @(posedge clk)
    begin
      if (write_to_ram)
          rmw_temp[23 : 16] <= dm_captured[2] ? mem_bytes[23 : 16] : dq_captured[23 : 16];
    end


  always @(posedge clk)
    begin
      if (write_to_ram)
          rmw_temp[31 : 24] <= dm_captured[3] ? mem_bytes[31 : 24] : dq_captured[31 : 24];
    end


  assign mem_bytes = (rmw_address == wr_addr_delayed && write_to_ram_r) ? rmw_temp : read_data;
  assign rmw_address = (write_to_ram) ? wr_addr_pipe_1 : read_addr_delayed;
  assign wr_addr_delayed = wr_addr_pipe_2;
  //use index to select which pipeline stage drives addr
  assign read_addr_delayed = (index == 0)? rd_addr_pipe_0 :
    (index == 1)? rd_addr_pipe_1 :
    (index == 2)? rd_addr_pipe_2 :
    (index == 3)? rd_addr_pipe_3 :
    (index == 4)? rd_addr_pipe_4 :
    rd_addr_pipe_5;

  //use index to select which pipeline stage drives valid
  assign read_valid = (index == 0)? rd_valid_pipe[0] :
    (index == 1)? rd_valid_pipe[1] :
    (index == 2)? rd_valid_pipe[2] :
    (index == 3)? rd_valid_pipe[3] :
    (index == 4)? rd_valid_pipe[4] :
    rd_valid_pipe[5];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign txt_code = (cmd_code == 3'h0)? 24'h4c4d52 :
    (cmd_code == 3'h1)? 24'h415246 :
    (cmd_code == 3'h2)? 24'h505245 :
    (cmd_code == 3'h3)? 24'h414354 :
    (cmd_code == 3'h4)? 24'h205752 :
    (cmd_code == 3'h5)? 24'h205244 :
    (cmd_code == 3'h6)? 24'h425354 :
    (cmd_code == 3'h7)? 24'h4e4f50 :
    24'h424144;


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


/* SLline 20484 "custom_dma.v" 2 */
/* SLline 1 "cpu_test_bench.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_test_bench (
                        // inputs:
                         A_bstatus_reg,
                         A_cmp_result,
                         A_ctrl_exception,
                         A_ctrl_ld_non_bypass,
                         A_dst_regnum,
                         A_en,
                         A_estatus_reg,
                         A_ienable_reg,
                         A_ipending_reg,
                         A_iw,
                         A_mem_byte_en,
                         A_op_hbreak,
                         A_op_intr,
                         A_pcb,
                         A_st_data,
                         A_status_reg,
                         A_valid,
                         A_wr_data_unfiltered,
                         A_wr_dst_reg,
                         E_add_br_to_taken_history_unfiltered,
                         E_logic_result,
                         E_valid,
                         M_bht_ptr_unfiltered,
                         M_bht_wr_data_unfiltered,
                         M_bht_wr_en_unfiltered,
                         M_mem_baddr,
                         M_target_pcb,
                         M_valid,
                         W_dst_regnum,
                         W_iw,
                         W_iw_op,
                         W_iw_opx,
                         W_pcb,
                         W_valid,
                         W_vinst,
                         W_wr_dst_reg,
                         clk,
                         d_address,
                         d_byteenable,
                         d_read,
                         d_write,
                         i_address,
                         i_read,
                         i_readdatavalid,
                         reset_n,

                        // outputs:
                         A_wr_data_filtered,
                         E_add_br_to_taken_history_filtered,
                         E_src1_eq_src2,
                         M_bht_ptr_filtered,
                         M_bht_wr_data_filtered,
                         M_bht_wr_en_filtered,
                         test_has_ended
                      )
;

  output  [ 31: 0] A_wr_data_filtered;
  output           E_add_br_to_taken_history_filtered;
  output           E_src1_eq_src2;
  output  [  7: 0] M_bht_ptr_filtered;
  output  [  1: 0] M_bht_wr_data_filtered;
  output           M_bht_wr_en_filtered;
  output           test_has_ended;
  input   [ 31: 0] A_bstatus_reg;
  input            A_cmp_result;
  input            A_ctrl_exception;
  input            A_ctrl_ld_non_bypass;
  input   [  4: 0] A_dst_regnum;
  input            A_en;
  input   [ 31: 0] A_estatus_reg;
  input   [ 31: 0] A_ienable_reg;
  input   [ 31: 0] A_ipending_reg;
  input   [ 31: 0] A_iw;
  input   [  3: 0] A_mem_byte_en;
  input            A_op_hbreak;
  input            A_op_intr;
  input   [ 26: 0] A_pcb;
  input   [ 31: 0] A_st_data;
  input   [ 31: 0] A_status_reg;
  input            A_valid;
  input   [ 31: 0] A_wr_data_unfiltered;
  input            A_wr_dst_reg;
  input            E_add_br_to_taken_history_unfiltered;
  input   [ 31: 0] E_logic_result;
  input            E_valid;
  input   [  7: 0] M_bht_ptr_unfiltered;
  input   [  1: 0] M_bht_wr_data_unfiltered;
  input            M_bht_wr_en_unfiltered;
  input   [ 26: 0] M_mem_baddr;
  input   [ 26: 0] M_target_pcb;
  input            M_valid;
  input   [  4: 0] W_dst_regnum;
  input   [ 31: 0] W_iw;
  input   [  5: 0] W_iw_op;
  input   [  5: 0] W_iw_opx;
  input   [ 26: 0] W_pcb;
  input            W_valid;
  input   [ 55: 0] W_vinst;
  input            W_wr_dst_reg;
  input            clk;
  input   [ 26: 0] d_address;
  input   [  3: 0] d_byteenable;
  input            d_read;
  input            d_write;
  input   [ 26: 0] i_address;
  input            i_read;
  input            i_readdatavalid;
  input            reset_n;

  reg     [ 26: 0] A_mem_baddr;
  reg     [ 26: 0] A_target_pcb;
  wire    [ 31: 0] A_wr_data_filtered;
  wire             A_wr_data_unfiltered_0_is_x;
  wire             A_wr_data_unfiltered_10_is_x;
  wire             A_wr_data_unfiltered_11_is_x;
  wire             A_wr_data_unfiltered_12_is_x;
  wire             A_wr_data_unfiltered_13_is_x;
  wire             A_wr_data_unfiltered_14_is_x;
  wire             A_wr_data_unfiltered_15_is_x;
  wire             A_wr_data_unfiltered_16_is_x;
  wire             A_wr_data_unfiltered_17_is_x;
  wire             A_wr_data_unfiltered_18_is_x;
  wire             A_wr_data_unfiltered_19_is_x;
  wire             A_wr_data_unfiltered_1_is_x;
  wire             A_wr_data_unfiltered_20_is_x;
  wire             A_wr_data_unfiltered_21_is_x;
  wire             A_wr_data_unfiltered_22_is_x;
  wire             A_wr_data_unfiltered_23_is_x;
  wire             A_wr_data_unfiltered_24_is_x;
  wire             A_wr_data_unfiltered_25_is_x;
  wire             A_wr_data_unfiltered_26_is_x;
  wire             A_wr_data_unfiltered_27_is_x;
  wire             A_wr_data_unfiltered_28_is_x;
  wire             A_wr_data_unfiltered_29_is_x;
  wire             A_wr_data_unfiltered_2_is_x;
  wire             A_wr_data_unfiltered_30_is_x;
  wire             A_wr_data_unfiltered_31_is_x;
  wire             A_wr_data_unfiltered_3_is_x;
  wire             A_wr_data_unfiltered_4_is_x;
  wire             A_wr_data_unfiltered_5_is_x;
  wire             A_wr_data_unfiltered_6_is_x;
  wire             A_wr_data_unfiltered_7_is_x;
  wire             A_wr_data_unfiltered_8_is_x;
  wire             A_wr_data_unfiltered_9_is_x;
  wire             E_add_br_to_taken_history_filtered;
  wire             E_src1_eq_src2;
  wire    [  7: 0] M_bht_ptr_filtered;
  wire    [  1: 0] M_bht_wr_data_filtered;
  wire             M_bht_wr_en_filtered;
  wire             W_op_add;
  wire             W_op_addi;
  wire             W_op_and;
  wire             W_op_andhi;
  wire             W_op_andi;
  wire             W_op_beq;
  wire             W_op_bge;
  wire             W_op_bgeu;
  wire             W_op_blt;
  wire             W_op_bltu;
  wire             W_op_bne;
  wire             W_op_br;
  wire             W_op_break;
  wire             W_op_bret;
  wire             W_op_call;
  wire             W_op_callr;
  wire             W_op_cmpeq;
  wire             W_op_cmpeqi;
  wire             W_op_cmpge;
  wire             W_op_cmpgei;
  wire             W_op_cmpgeu;
  wire             W_op_cmpgeui;
  wire             W_op_cmplt;
  wire             W_op_cmplti;
  wire             W_op_cmpltu;
  wire             W_op_cmpltui;
  wire             W_op_cmpne;
  wire             W_op_cmpnei;
  wire             W_op_crst;
  wire             W_op_custom;
  wire             W_op_div;
  wire             W_op_divu;
  wire             W_op_eret;
  wire             W_op_flushd;
  wire             W_op_flushda;
  wire             W_op_flushi;
  wire             W_op_flushp;
  wire             W_op_hbreak;
  wire             W_op_initd;
  wire             W_op_initda;
  wire             W_op_initi;
  wire             W_op_intr;
  wire             W_op_jmp;
  wire             W_op_jmpi;
  wire             W_op_ldb;
  wire             W_op_ldbio;
  wire             W_op_ldbu;
  wire             W_op_ldbuio;
  wire             W_op_ldh;
  wire             W_op_ldhio;
  wire             W_op_ldhu;
  wire             W_op_ldhuio;
  wire             W_op_ldl;
  wire             W_op_ldw;
  wire             W_op_ldwio;
  wire             W_op_mul;
  wire             W_op_muli;
  wire             W_op_mulxss;
  wire             W_op_mulxsu;
  wire             W_op_mulxuu;
  wire             W_op_nextpc;
  wire             W_op_nor;
  wire             W_op_opx;
  wire             W_op_or;
  wire             W_op_orhi;
  wire             W_op_ori;
  wire             W_op_rdctl;
  wire             W_op_rdprs;
  wire             W_op_ret;
  wire             W_op_rol;
  wire             W_op_roli;
  wire             W_op_ror;
  wire             W_op_rsv02;
  wire             W_op_rsv09;
  wire             W_op_rsv10;
  wire             W_op_rsv17;
  wire             W_op_rsv18;
  wire             W_op_rsv25;
  wire             W_op_rsv26;
  wire             W_op_rsv33;
  wire             W_op_rsv34;
  wire             W_op_rsv41;
  wire             W_op_rsv42;
  wire             W_op_rsv49;
  wire             W_op_rsv57;
  wire             W_op_rsv61;
  wire             W_op_rsv62;
  wire             W_op_rsv63;
  wire             W_op_rsvx00;
  wire             W_op_rsvx10;
  wire             W_op_rsvx15;
  wire             W_op_rsvx17;
  wire             W_op_rsvx21;
  wire             W_op_rsvx25;
  wire             W_op_rsvx33;
  wire             W_op_rsvx34;
  wire             W_op_rsvx35;
  wire             W_op_rsvx42;
  wire             W_op_rsvx43;
  wire             W_op_rsvx44;
  wire             W_op_rsvx47;
  wire             W_op_rsvx50;
  wire             W_op_rsvx51;
  wire             W_op_rsvx55;
  wire             W_op_rsvx56;
  wire             W_op_rsvx60;
  wire             W_op_rsvx63;
  wire             W_op_sll;
  wire             W_op_slli;
  wire             W_op_sra;
  wire             W_op_srai;
  wire             W_op_srl;
  wire             W_op_srli;
  wire             W_op_stb;
  wire             W_op_stbio;
  wire             W_op_stc;
  wire             W_op_sth;
  wire             W_op_sthio;
  wire             W_op_stw;
  wire             W_op_stwio;
  wire             W_op_sub;
  wire             W_op_sync;
  wire             W_op_trap;
  wire             W_op_wrctl;
  wire             W_op_wrprs;
  wire             W_op_xor;
  wire             W_op_xorhi;
  wire             W_op_xori;
  wire             test_has_ended;
  assign W_op_call = W_iw_op == 0;
  assign W_op_jmpi = W_iw_op == 1;
  assign W_op_ldbu = W_iw_op == 3;
  assign W_op_addi = W_iw_op == 4;
  assign W_op_stb = W_iw_op == 5;
  assign W_op_br = W_iw_op == 6;
  assign W_op_ldb = W_iw_op == 7;
  assign W_op_cmpgei = W_iw_op == 8;
  assign W_op_ldhu = W_iw_op == 11;
  assign W_op_andi = W_iw_op == 12;
  assign W_op_sth = W_iw_op == 13;
  assign W_op_bge = W_iw_op == 14;
  assign W_op_ldh = W_iw_op == 15;
  assign W_op_cmplti = W_iw_op == 16;
  assign W_op_initda = W_iw_op == 19;
  assign W_op_ori = W_iw_op == 20;
  assign W_op_stw = W_iw_op == 21;
  assign W_op_blt = W_iw_op == 22;
  assign W_op_ldw = W_iw_op == 23;
  assign W_op_cmpnei = W_iw_op == 24;
  assign W_op_flushda = W_iw_op == 27;
  assign W_op_xori = W_iw_op == 28;
  assign W_op_stc = W_iw_op == 29;
  assign W_op_bne = W_iw_op == 30;
  assign W_op_ldl = W_iw_op == 31;
  assign W_op_cmpeqi = W_iw_op == 32;
  assign W_op_ldbuio = W_iw_op == 35;
  assign W_op_muli = W_iw_op == 36;
  assign W_op_stbio = W_iw_op == 37;
  assign W_op_beq = W_iw_op == 38;
  assign W_op_ldbio = W_iw_op == 39;
  assign W_op_cmpgeui = W_iw_op == 40;
  assign W_op_ldhuio = W_iw_op == 43;
  assign W_op_andhi = W_iw_op == 44;
  assign W_op_sthio = W_iw_op == 45;
  assign W_op_bgeu = W_iw_op == 46;
  assign W_op_ldhio = W_iw_op == 47;
  assign W_op_cmpltui = W_iw_op == 48;
  assign W_op_initd = W_iw_op == 51;
  assign W_op_orhi = W_iw_op == 52;
  assign W_op_stwio = W_iw_op == 53;
  assign W_op_bltu = W_iw_op == 54;
  assign W_op_ldwio = W_iw_op == 55;
  assign W_op_rdprs = W_iw_op == 56;
  assign W_op_flushd = W_iw_op == 59;
  assign W_op_xorhi = W_iw_op == 60;
  assign W_op_rsv02 = W_iw_op == 2;
  assign W_op_rsv09 = W_iw_op == 9;
  assign W_op_rsv10 = W_iw_op == 10;
  assign W_op_rsv17 = W_iw_op == 17;
  assign W_op_rsv18 = W_iw_op == 18;
  assign W_op_rsv25 = W_iw_op == 25;
  assign W_op_rsv26 = W_iw_op == 26;
  assign W_op_rsv33 = W_iw_op == 33;
  assign W_op_rsv34 = W_iw_op == 34;
  assign W_op_rsv41 = W_iw_op == 41;
  assign W_op_rsv42 = W_iw_op == 42;
  assign W_op_rsv49 = W_iw_op == 49;
  assign W_op_rsv57 = W_iw_op == 57;
  assign W_op_rsv61 = W_iw_op == 61;
  assign W_op_rsv62 = W_iw_op == 62;
  assign W_op_rsv63 = W_iw_op == 63;
  assign W_op_eret = W_op_opx & (W_iw_opx == 1);
  assign W_op_roli = W_op_opx & (W_iw_opx == 2);
  assign W_op_rol = W_op_opx & (W_iw_opx == 3);
  assign W_op_flushp = W_op_opx & (W_iw_opx == 4);
  assign W_op_ret = W_op_opx & (W_iw_opx == 5);
  assign W_op_nor = W_op_opx & (W_iw_opx == 6);
  assign W_op_mulxuu = W_op_opx & (W_iw_opx == 7);
  assign W_op_cmpge = W_op_opx & (W_iw_opx == 8);
  assign W_op_bret = W_op_opx & (W_iw_opx == 9);
  assign W_op_ror = W_op_opx & (W_iw_opx == 11);
  assign W_op_flushi = W_op_opx & (W_iw_opx == 12);
  assign W_op_jmp = W_op_opx & (W_iw_opx == 13);
  assign W_op_and = W_op_opx & (W_iw_opx == 14);
  assign W_op_cmplt = W_op_opx & (W_iw_opx == 16);
  assign W_op_slli = W_op_opx & (W_iw_opx == 18);
  assign W_op_sll = W_op_opx & (W_iw_opx == 19);
  assign W_op_wrprs = W_op_opx & (W_iw_opx == 20);
  assign W_op_or = W_op_opx & (W_iw_opx == 22);
  assign W_op_mulxsu = W_op_opx & (W_iw_opx == 23);
  assign W_op_cmpne = W_op_opx & (W_iw_opx == 24);
  assign W_op_srli = W_op_opx & (W_iw_opx == 26);
  assign W_op_srl = W_op_opx & (W_iw_opx == 27);
  assign W_op_nextpc = W_op_opx & (W_iw_opx == 28);
  assign W_op_callr = W_op_opx & (W_iw_opx == 29);
  assign W_op_xor = W_op_opx & (W_iw_opx == 30);
  assign W_op_mulxss = W_op_opx & (W_iw_opx == 31);
  assign W_op_cmpeq = W_op_opx & (W_iw_opx == 32);
  assign W_op_divu = W_op_opx & (W_iw_opx == 36);
  assign W_op_div = W_op_opx & (W_iw_opx == 37);
  assign W_op_rdctl = W_op_opx & (W_iw_opx == 38);
  assign W_op_mul = W_op_opx & (W_iw_opx == 39);
  assign W_op_cmpgeu = W_op_opx & (W_iw_opx == 40);
  assign W_op_initi = W_op_opx & (W_iw_opx == 41);
  assign W_op_trap = W_op_opx & (W_iw_opx == 45);
  assign W_op_wrctl = W_op_opx & (W_iw_opx == 46);
  assign W_op_cmpltu = W_op_opx & (W_iw_opx == 48);
  assign W_op_add = W_op_opx & (W_iw_opx == 49);
  assign W_op_break = W_op_opx & (W_iw_opx == 52);
  assign W_op_hbreak = W_op_opx & (W_iw_opx == 53);
  assign W_op_sync = W_op_opx & (W_iw_opx == 54);
  assign W_op_sub = W_op_opx & (W_iw_opx == 57);
  assign W_op_srai = W_op_opx & (W_iw_opx == 58);
  assign W_op_sra = W_op_opx & (W_iw_opx == 59);
  assign W_op_intr = W_op_opx & (W_iw_opx == 61);
  assign W_op_crst = W_op_opx & (W_iw_opx == 62);
  assign W_op_rsvx00 = W_op_opx & (W_iw_opx == 0);
  assign W_op_rsvx10 = W_op_opx & (W_iw_opx == 10);
  assign W_op_rsvx15 = W_op_opx & (W_iw_opx == 15);
  assign W_op_rsvx17 = W_op_opx & (W_iw_opx == 17);
  assign W_op_rsvx21 = W_op_opx & (W_iw_opx == 21);
  assign W_op_rsvx25 = W_op_opx & (W_iw_opx == 25);
  assign W_op_rsvx33 = W_op_opx & (W_iw_opx == 33);
  assign W_op_rsvx34 = W_op_opx & (W_iw_opx == 34);
  assign W_op_rsvx35 = W_op_opx & (W_iw_opx == 35);
  assign W_op_rsvx42 = W_op_opx & (W_iw_opx == 42);
  assign W_op_rsvx43 = W_op_opx & (W_iw_opx == 43);
  assign W_op_rsvx44 = W_op_opx & (W_iw_opx == 44);
  assign W_op_rsvx47 = W_op_opx & (W_iw_opx == 47);
  assign W_op_rsvx50 = W_op_opx & (W_iw_opx == 50);
  assign W_op_rsvx51 = W_op_opx & (W_iw_opx == 51);
  assign W_op_rsvx55 = W_op_opx & (W_iw_opx == 55);
  assign W_op_rsvx56 = W_op_opx & (W_iw_opx == 56);
  assign W_op_rsvx60 = W_op_opx & (W_iw_opx == 60);
  assign W_op_rsvx63 = W_op_opx & (W_iw_opx == 63);
  assign W_op_opx = W_iw_op == 58;
  assign W_op_custom = W_iw_op == 50;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          A_target_pcb <= 0;
      else if (A_en)
          A_target_pcb <= M_target_pcb;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          A_mem_baddr <= 0;
      else if (A_en)
          A_mem_baddr <= M_mem_baddr;
    end


  assign E_src1_eq_src2 = E_logic_result == 0;
  //Propagating 'X' data bits
  assign E_add_br_to_taken_history_filtered = E_add_br_to_taken_history_unfiltered;

  //Propagating 'X' data bits
  assign M_bht_wr_en_filtered = M_bht_wr_en_unfiltered;

  //Propagating 'X' data bits
  assign M_bht_wr_data_filtered = M_bht_wr_data_unfiltered;

  //Propagating 'X' data bits
  assign M_bht_ptr_filtered = M_bht_ptr_unfiltered;

  assign test_has_ended = 1'b0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //Clearing 'X' data bits
  assign A_wr_data_unfiltered_0_is_x = ^(A_wr_data_unfiltered[0]) === 1'bx;

  assign A_wr_data_filtered[0] = (A_wr_data_unfiltered_0_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[0];
  assign A_wr_data_unfiltered_1_is_x = ^(A_wr_data_unfiltered[1]) === 1'bx;
  assign A_wr_data_filtered[1] = (A_wr_data_unfiltered_1_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[1];
  assign A_wr_data_unfiltered_2_is_x = ^(A_wr_data_unfiltered[2]) === 1'bx;
  assign A_wr_data_filtered[2] = (A_wr_data_unfiltered_2_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[2];
  assign A_wr_data_unfiltered_3_is_x = ^(A_wr_data_unfiltered[3]) === 1'bx;
  assign A_wr_data_filtered[3] = (A_wr_data_unfiltered_3_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[3];
  assign A_wr_data_unfiltered_4_is_x = ^(A_wr_data_unfiltered[4]) === 1'bx;
  assign A_wr_data_filtered[4] = (A_wr_data_unfiltered_4_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[4];
  assign A_wr_data_unfiltered_5_is_x = ^(A_wr_data_unfiltered[5]) === 1'bx;
  assign A_wr_data_filtered[5] = (A_wr_data_unfiltered_5_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[5];
  assign A_wr_data_unfiltered_6_is_x = ^(A_wr_data_unfiltered[6]) === 1'bx;
  assign A_wr_data_filtered[6] = (A_wr_data_unfiltered_6_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[6];
  assign A_wr_data_unfiltered_7_is_x = ^(A_wr_data_unfiltered[7]) === 1'bx;
  assign A_wr_data_filtered[7] = (A_wr_data_unfiltered_7_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[7];
  assign A_wr_data_unfiltered_8_is_x = ^(A_wr_data_unfiltered[8]) === 1'bx;
  assign A_wr_data_filtered[8] = (A_wr_data_unfiltered_8_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[8];
  assign A_wr_data_unfiltered_9_is_x = ^(A_wr_data_unfiltered[9]) === 1'bx;
  assign A_wr_data_filtered[9] = (A_wr_data_unfiltered_9_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[9];
  assign A_wr_data_unfiltered_10_is_x = ^(A_wr_data_unfiltered[10]) === 1'bx;
  assign A_wr_data_filtered[10] = (A_wr_data_unfiltered_10_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[10];
  assign A_wr_data_unfiltered_11_is_x = ^(A_wr_data_unfiltered[11]) === 1'bx;
  assign A_wr_data_filtered[11] = (A_wr_data_unfiltered_11_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[11];
  assign A_wr_data_unfiltered_12_is_x = ^(A_wr_data_unfiltered[12]) === 1'bx;
  assign A_wr_data_filtered[12] = (A_wr_data_unfiltered_12_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[12];
  assign A_wr_data_unfiltered_13_is_x = ^(A_wr_data_unfiltered[13]) === 1'bx;
  assign A_wr_data_filtered[13] = (A_wr_data_unfiltered_13_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[13];
  assign A_wr_data_unfiltered_14_is_x = ^(A_wr_data_unfiltered[14]) === 1'bx;
  assign A_wr_data_filtered[14] = (A_wr_data_unfiltered_14_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[14];
  assign A_wr_data_unfiltered_15_is_x = ^(A_wr_data_unfiltered[15]) === 1'bx;
  assign A_wr_data_filtered[15] = (A_wr_data_unfiltered_15_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[15];
  assign A_wr_data_unfiltered_16_is_x = ^(A_wr_data_unfiltered[16]) === 1'bx;
  assign A_wr_data_filtered[16] = (A_wr_data_unfiltered_16_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[16];
  assign A_wr_data_unfiltered_17_is_x = ^(A_wr_data_unfiltered[17]) === 1'bx;
  assign A_wr_data_filtered[17] = (A_wr_data_unfiltered_17_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[17];
  assign A_wr_data_unfiltered_18_is_x = ^(A_wr_data_unfiltered[18]) === 1'bx;
  assign A_wr_data_filtered[18] = (A_wr_data_unfiltered_18_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[18];
  assign A_wr_data_unfiltered_19_is_x = ^(A_wr_data_unfiltered[19]) === 1'bx;
  assign A_wr_data_filtered[19] = (A_wr_data_unfiltered_19_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[19];
  assign A_wr_data_unfiltered_20_is_x = ^(A_wr_data_unfiltered[20]) === 1'bx;
  assign A_wr_data_filtered[20] = (A_wr_data_unfiltered_20_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[20];
  assign A_wr_data_unfiltered_21_is_x = ^(A_wr_data_unfiltered[21]) === 1'bx;
  assign A_wr_data_filtered[21] = (A_wr_data_unfiltered_21_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[21];
  assign A_wr_data_unfiltered_22_is_x = ^(A_wr_data_unfiltered[22]) === 1'bx;
  assign A_wr_data_filtered[22] = (A_wr_data_unfiltered_22_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[22];
  assign A_wr_data_unfiltered_23_is_x = ^(A_wr_data_unfiltered[23]) === 1'bx;
  assign A_wr_data_filtered[23] = (A_wr_data_unfiltered_23_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[23];
  assign A_wr_data_unfiltered_24_is_x = ^(A_wr_data_unfiltered[24]) === 1'bx;
  assign A_wr_data_filtered[24] = (A_wr_data_unfiltered_24_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[24];
  assign A_wr_data_unfiltered_25_is_x = ^(A_wr_data_unfiltered[25]) === 1'bx;
  assign A_wr_data_filtered[25] = (A_wr_data_unfiltered_25_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[25];
  assign A_wr_data_unfiltered_26_is_x = ^(A_wr_data_unfiltered[26]) === 1'bx;
  assign A_wr_data_filtered[26] = (A_wr_data_unfiltered_26_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[26];
  assign A_wr_data_unfiltered_27_is_x = ^(A_wr_data_unfiltered[27]) === 1'bx;
  assign A_wr_data_filtered[27] = (A_wr_data_unfiltered_27_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[27];
  assign A_wr_data_unfiltered_28_is_x = ^(A_wr_data_unfiltered[28]) === 1'bx;
  assign A_wr_data_filtered[28] = (A_wr_data_unfiltered_28_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[28];
  assign A_wr_data_unfiltered_29_is_x = ^(A_wr_data_unfiltered[29]) === 1'bx;
  assign A_wr_data_filtered[29] = (A_wr_data_unfiltered_29_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[29];
  assign A_wr_data_unfiltered_30_is_x = ^(A_wr_data_unfiltered[30]) === 1'bx;
  assign A_wr_data_filtered[30] = (A_wr_data_unfiltered_30_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[30];
  assign A_wr_data_unfiltered_31_is_x = ^(A_wr_data_unfiltered[31]) === 1'bx;
  assign A_wr_data_filtered[31] = (A_wr_data_unfiltered_31_is_x & (A_ctrl_ld_non_bypass)) ? 1'b0 : A_wr_data_unfiltered[31];
  always @(posedge clk)
    begin
      if (reset_n)
          if (^(W_wr_dst_reg) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/W_wr_dst_reg is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (W_wr_dst_reg)
          if (^(W_dst_regnum) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/W_dst_regnum is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(W_valid) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/W_valid is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (W_valid)
          if (^(W_pcb) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/W_pcb is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (W_valid)
          if (^(W_iw) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/W_iw is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(A_en) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/A_en is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(E_valid) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/E_valid is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(M_valid) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/M_valid is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(A_valid) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/A_valid is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (A_valid & A_en & A_wr_dst_reg)
          if (^(A_wr_data_unfiltered) === 1'bx)
            begin
              $write("%0d ns: WARNING: cpu_test_bench/A_wr_data_unfiltered is 'x'\n", $time);
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(A_status_reg) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/A_status_reg is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(A_estatus_reg) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/A_estatus_reg is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(A_bstatus_reg) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/A_bstatus_reg is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(i_read) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/i_read is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (i_read)
          if (^(i_address) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/i_address is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(i_readdatavalid) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/i_readdatavalid is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(d_write) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/d_write is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (d_write)
          if (^(d_byteenable) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/d_byteenable is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
        begin
        end
      else if (d_write | d_read)
          if (^(d_address) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/d_address is 'x'\n", $time);
              $stop;
            end
    end


  always @(posedge clk)
    begin
      if (reset_n)
          if (^(d_read) === 1'bx)
            begin
              $write("%0d ns: ERROR: cpu_test_bench/d_read is 'x'\n", $time);
              $stop;
            end
    end


  
  reg [31:0] trace_handle; // for $fopen
  initial  
  begin
    trace_handle = $fopen("cpu.tr");
    $fwrite(trace_handle, "version 3\nnumThreads 1\n");
  end
  always @(posedge clk)
    begin
      if ((~reset_n || (A_valid & A_en)) && ~test_has_ended)
          $fwrite(trace_handle, "%0d ns: %0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h,%0h\n", $time, ~reset_n, A_pcb, 0, A_op_intr, A_op_hbreak, A_iw, ~(A_op_intr | A_op_hbreak), A_wr_dst_reg, A_dst_regnum, 0, A_wr_data_filtered, A_mem_baddr, A_st_data, A_mem_byte_en, A_cmp_result, A_target_pcb, A_status_reg, A_estatus_reg, A_bstatus_reg, A_ienable_reg, A_ipending_reg, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, A_ctrl_exception ? 1 : 0, 0, 0, 0, 0);
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign A_wr_data_filtered = A_wr_data_unfiltered;
//
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20485 "custom_dma.v" 2 */
/* SLline 1 "cpu_mult_cell.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_mult_cell (
                       // inputs:
                        A_en,
                        E_ctrl_mul_shift_src1_signed,
                        E_ctrl_mul_shift_src2_signed,
                        E_src1_mul_cell,
                        E_src2_mul_cell,
                        M_en,
                        clk,
                        reset_n,

                       // outputs:
                        A_mul_cell_result
                     )
;

  output  [ 63: 0] A_mul_cell_result;
  input            A_en;
  input            E_ctrl_mul_shift_src1_signed;
  input            E_ctrl_mul_shift_src2_signed;
  input   [ 31: 0] E_src1_mul_cell;
  input   [ 31: 0] E_src2_mul_cell;
  input            M_en;
  input            clk;
  input            reset_n;

  wire    [ 63: 0] A_mul_cell_result;
  wire             mul_clr;
  assign mul_clr = ~reset_n;
  altmult_add the_altmult_add
    (
      .aclr0 (mul_clr),
      .aclr1 (mul_clr),
      .clock0 (clk),
      .clock1 (clk),
      .dataa (E_src1_mul_cell),
      .datab (E_src2_mul_cell),
      .ena0 (M_en),
      .ena1 (A_en),
      .result (A_mul_cell_result),
      .signa (E_ctrl_mul_shift_src1_signed),
      .signb (E_ctrl_mul_shift_src2_signed)
    );

  defparam the_altmult_add.addnsub_multiplier_aclr1 = "UNUSED",
           the_altmult_add.addnsub_multiplier_pipeline_aclr1 = "UNUSED",
           the_altmult_add.addnsub_multiplier_register1 = "CLOCK0",
           the_altmult_add.dedicated_multiplier_circuitry = "YES",
           the_altmult_add.input_aclr_a0 = "ACLR0",
           the_altmult_add.input_aclr_b0 = "ACLR0",
           the_altmult_add.input_register_a0 = "CLOCK0",
           the_altmult_add.input_register_b0 = "CLOCK0",
           the_altmult_add.input_source_a0 = "DATAA",
           the_altmult_add.input_source_b0 = "DATAB",
           the_altmult_add.intended_device_family = "STRATIXII",
           the_altmult_add.lpm_type = "altmult_add",
           the_altmult_add.multiplier1_direction = "ADD",
           the_altmult_add.multiplier_register0 = "UNREGISTERED",
           the_altmult_add.number_of_multipliers = 1,
           the_altmult_add.output_aclr = "ACLR1",
           the_altmult_add.output_register = "CLOCK1",
           the_altmult_add.signed_aclr_a = "ACLR0",
           the_altmult_add.signed_aclr_b = "ACLR0",
           the_altmult_add.signed_pipeline_register_a = "UNREGISTERED",
           the_altmult_add.signed_pipeline_register_b = "UNREGISTERED",
           the_altmult_add.signed_register_a = "CLOCK0",
           the_altmult_add.signed_register_b = "CLOCK0",
           the_altmult_add.width_a = 32,
           the_altmult_add.width_b = 32,
           the_altmult_add.width_result = 64;


endmodule


/* SLline 20486 "custom_dma.v" 2 */
/* SLline 1 "cpu_oci_test_bench.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_oci_test_bench (
                            // inputs:
                             dct_buffer,
                             dct_count,
                             test_ending,
                             test_has_ended
                          )
;

  input   [ 29: 0] dct_buffer;
  input   [  3: 0] dct_count;
  input            test_ending;
  input            test_has_ended;


endmodule


/* SLline 20487 "custom_dma.v" 2 */
/* SLline 1 "cpu_jtag_debug_module_tck.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_tck (
                                   // inputs:
                                    MonDReg,
                                    break_readreg,
                                    dbrk_hit0_latch,
                                    dbrk_hit1_latch,
                                    dbrk_hit2_latch,
                                    dbrk_hit3_latch,
                                    debugack,
                                    ir_in,
                                    jtag_state_rti,
                                    monitor_error,
                                    monitor_ready,
                                    reset_n,
                                    resetlatch,
                                    tck,
                                    tdi,
                                    tracemem_on,
                                    tracemem_trcdata,
                                    tracemem_tw,
                                    trc_im_addr,
                                    trc_on,
                                    trc_wrap,
                                    trigbrktype,
                                    trigger_state_1,
                                    vs_cdr,
                                    vs_sdr,
                                    vs_uir,

                                   // outputs:
                                    ir_out,
                                    jrst_n,
                                    sr,
                                    st_ready_test_idle,
                                    tdo
                                 )
;

  output  [  1: 0] ir_out;
  output           jrst_n;
  output  [ 37: 0] sr;
  output           st_ready_test_idle;
  output           tdo;
  input   [ 31: 0] MonDReg;
  input   [ 31: 0] break_readreg;
  input            dbrk_hit0_latch;
  input            dbrk_hit1_latch;
  input            dbrk_hit2_latch;
  input            dbrk_hit3_latch;
  input            debugack;
  input   [  1: 0] ir_in;
  input            jtag_state_rti;
  input            monitor_error;
  input            monitor_ready;
  input            reset_n;
  input            resetlatch;
  input            tck;
  input            tdi;
  input            tracemem_on;
  input   [ 35: 0] tracemem_trcdata;
  input            tracemem_tw;
  input   [  6: 0] trc_im_addr;
  input            trc_on;
  input            trc_wrap;
  input            trigbrktype;
  input            trigger_state_1;
  input            vs_cdr;
  input            vs_sdr;
  input            vs_uir;

  reg     [  2: 0] DRsize /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103,R101\""  */;
  wire             debugack_sync;
  reg     [  1: 0] ir_out;
  wire             jrst_n;
  wire             monitor_ready_sync;
  reg     [ 37: 0] sr /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103,R101\""  */;
  wire             st_ready_test_idle;
  wire             tdo;
  wire             unxcomplemented_resetxx0;
  wire             unxcomplemented_resetxx1;
  always @(posedge tck)
    begin
      if (vs_cdr)
          case (ir_in)
          
              2'b00: begin
                  sr[35] <= debugack_sync;
                  sr[34] <= monitor_error;
                  sr[33] <= resetlatch;
                  sr[32 : 1] <= MonDReg;
                  sr[0] <= monitor_ready_sync;
              end // 2'b00 
          
              2'b01: begin
                  sr[35 : 0] <= tracemem_trcdata;
                  sr[37] <= tracemem_tw;
                  sr[36] <= tracemem_on;
              end // 2'b01 
          
              2'b10: begin
                  sr[37] <= trigger_state_1;
                  sr[36] <= dbrk_hit3_latch;
                  sr[35] <= dbrk_hit2_latch;
                  sr[34] <= dbrk_hit1_latch;
                  sr[33] <= dbrk_hit0_latch;
                  sr[32 : 1] <= break_readreg;
                  sr[0] <= trigbrktype;
              end // 2'b10 
          
              2'b11: begin
                  sr[15 : 12] <= 1'b0;
                  sr[11 : 2] <= trc_im_addr;
                  sr[1] <= trc_wrap;
                  sr[0] <= trc_on;
              end // 2'b11 
          
          endcase // ir_in
      if (vs_sdr)
          case (DRsize)
          
              3'b000: begin
                  sr <= {tdi, sr[37 : 2], tdi};
              end // 3'b000 
          
              3'b001: begin
                  sr <= {tdi, sr[37 : 9], tdi, sr[7 : 1]};
              end // 3'b001 
          
              3'b010: begin
                  sr <= {tdi, sr[37 : 17], tdi, sr[15 : 1]};
              end // 3'b010 
          
              3'b011: begin
                  sr <= {tdi, sr[37 : 33], tdi, sr[31 : 1]};
              end // 3'b011 
          
              3'b100: begin
                  sr <= {tdi, sr[37],         tdi, sr[35 : 1]};
              end // 3'b100 
          
              3'b101: begin
                  sr <= {tdi, sr[37 : 1]};
              end // 3'b101 
          
              default: begin
                  sr <= {tdi, sr[37 : 2], tdi};
              end // default
          
          endcase // DRsize
      if (vs_uir)
          case (ir_in)
          
              2'b00: begin
                  DRsize <= 3'b100;
              end // 2'b00 
          
              2'b01: begin
                  DRsize <= 3'b101;
              end // 2'b01 
          
              2'b10: begin
                  DRsize <= 3'b101;
              end // 2'b10 
          
              2'b11: begin
                  DRsize <= 3'b010;
              end // 2'b11 
          
          endcase // ir_in
    end


  assign tdo = sr[0];
  assign st_ready_test_idle = jtag_state_rti;
  assign unxcomplemented_resetxx0 = jrst_n;
  altera_std_synchronizer the_altera_std_synchronizer
    (
      .clk (tck),
      .din (debugack),
      .dout (debugack_sync),
      .reset_n (unxcomplemented_resetxx0)
    );

  defparam the_altera_std_synchronizer.depth = 2;

  assign unxcomplemented_resetxx1 = jrst_n;
  altera_std_synchronizer the_altera_std_synchronizer1
    (
      .clk (tck),
      .din (monitor_ready),
      .dout (monitor_ready_sync),
      .reset_n (unxcomplemented_resetxx1)
    );

  defparam the_altera_std_synchronizer1.depth = 2;

  always @(posedge tck or negedge jrst_n)
    begin
      if (jrst_n == 0)
          ir_out <= 2'b0;
      else 
        ir_out <= {debugack_sync, monitor_ready_sync};
    end



//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign jrst_n = reset_n;

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  assign jrst_n = 1;
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20488 "custom_dma.v" 2 */
/* SLline 1 "cpu_jtag_debug_module_sysclk.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_sysclk (
                                      // inputs:
                                       clk,
                                       ir_in,
                                       sr,
                                       vs_udr,
                                       vs_uir,

                                      // outputs:
                                       jdo,
                                       take_action_break_a,
                                       take_action_break_b,
                                       take_action_break_c,
                                       take_action_ocimem_a,
                                       take_action_ocimem_b,
                                       take_action_tracectrl,
                                       take_action_tracemem_a,
                                       take_action_tracemem_b,
                                       take_no_action_break_a,
                                       take_no_action_break_b,
                                       take_no_action_break_c,
                                       take_no_action_ocimem_a,
                                       take_no_action_tracemem_a
                                    )
;

  output  [ 37: 0] jdo;
  output           take_action_break_a;
  output           take_action_break_b;
  output           take_action_break_c;
  output           take_action_ocimem_a;
  output           take_action_ocimem_b;
  output           take_action_tracectrl;
  output           take_action_tracemem_a;
  output           take_action_tracemem_b;
  output           take_no_action_break_a;
  output           take_no_action_break_b;
  output           take_no_action_break_c;
  output           take_no_action_ocimem_a;
  output           take_no_action_tracemem_a;
  input            clk;
  input   [  1: 0] ir_in;
  input   [ 37: 0] sr;
  input            vs_udr;
  input            vs_uir;

  reg              enable_action_strobe /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103\""  */;
  reg     [  1: 0] ir /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,R101\""  */;
  reg     [ 37: 0] jdo /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,R101\""  */;
  reg              jxuir /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103\""  */;
  reg              sync2_udr /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103\""  */;
  reg              sync2_uir /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103\""  */;
  wire             sync_udr;
  wire             sync_uir;
  wire             take_action_break_a;
  wire             take_action_break_b;
  wire             take_action_break_c;
  wire             take_action_ocimem_a;
  wire             take_action_ocimem_b;
  wire             take_action_tracectrl;
  wire             take_action_tracemem_a;
  wire             take_action_tracemem_b;
  wire             take_no_action_break_a;
  wire             take_no_action_break_b;
  wire             take_no_action_break_c;
  wire             take_no_action_ocimem_a;
  wire             take_no_action_tracemem_a;
  wire             unxunused_resetxx2;
  wire             unxunused_resetxx3;
  reg              update_jdo_strobe /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=\"D101,D103\""  */;
  assign unxunused_resetxx2 = 1'b1;
  altera_std_synchronizer the_altera_std_synchronizer2
    (
      .clk (clk),
      .din (vs_udr),
      .dout (sync_udr),
      .reset_n (unxunused_resetxx2)
    );

  defparam the_altera_std_synchronizer2.depth = 2;

  assign unxunused_resetxx3 = 1'b1;
  altera_std_synchronizer the_altera_std_synchronizer3
    (
      .clk (clk),
      .din (vs_uir),
      .dout (sync_uir),
      .reset_n (unxunused_resetxx3)
    );

  defparam the_altera_std_synchronizer3.depth = 2;

  always @(posedge clk)
    begin
      sync2_udr <= sync_udr;
      update_jdo_strobe <= sync_udr & ~sync2_udr;
      enable_action_strobe <= update_jdo_strobe;
      sync2_uir <= sync_uir;
      jxuir <= sync_uir & ~sync2_uir;
    end


  assign take_action_ocimem_a = enable_action_strobe && (ir == 2'b00) && 
    ~jdo[35] && jdo[34];

  assign take_no_action_ocimem_a = enable_action_strobe && (ir == 2'b00) && 
    ~jdo[35] && ~jdo[34];

  assign take_action_ocimem_b = enable_action_strobe && (ir == 2'b00) && 
    jdo[35];

  assign take_action_tracemem_a = enable_action_strobe && (ir == 2'b01) &&
    ~jdo[37] && 
    jdo[36];

  assign take_no_action_tracemem_a = enable_action_strobe && (ir == 2'b01) &&
    ~jdo[37] && 
    ~jdo[36];

  assign take_action_tracemem_b = enable_action_strobe && (ir == 2'b01) &&
    jdo[37];

  assign take_action_break_a = enable_action_strobe && (ir == 2'b10) && 
    ~jdo[36] && 
    jdo[37];

  assign take_no_action_break_a = enable_action_strobe && (ir == 2'b10) && 
    ~jdo[36] && 
    ~jdo[37];

  assign take_action_break_b = enable_action_strobe && (ir == 2'b10) && 
    jdo[36] && ~jdo[35] &&
    jdo[37];

  assign take_no_action_break_b = enable_action_strobe && (ir == 2'b10) && 
    jdo[36] && ~jdo[35] &&
    ~jdo[37];

  assign take_action_break_c = enable_action_strobe && (ir == 2'b10) && 
    jdo[36] &&  jdo[35] &&
    jdo[37];

  assign take_no_action_break_c = enable_action_strobe && (ir == 2'b10) && 
    jdo[36] &&  jdo[35] &&
    ~jdo[37];

  assign take_action_tracectrl = enable_action_strobe && (ir == 2'b11) &&  
    jdo[15];

  always @(posedge clk)
    begin
      if (jxuir)
          ir <= ir_in;
      if (update_jdo_strobe)
          jdo <= sr;
    end



endmodule


/* SLline 20489 "custom_dma.v" 2 */
/* SLline 1 "cpu_jtag_debug_module_wrapper.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.


// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_jtag_debug_module_wrapper (
                                       // inputs:
                                        MonDReg,
                                        break_readreg,
                                        clk,
                                        dbrk_hit0_latch,
                                        dbrk_hit1_latch,
                                        dbrk_hit2_latch,
                                        dbrk_hit3_latch,
                                        debugack,
                                        monitor_error,
                                        monitor_ready,
                                        reset_n,
                                        resetlatch,
                                        tracemem_on,
                                        tracemem_trcdata,
                                        tracemem_tw,
                                        trc_im_addr,
                                        trc_on,
                                        trc_wrap,
                                        trigbrktype,
                                        trigger_state_1,

                                       // outputs:
                                        jdo,
                                        jrst_n,
                                        st_ready_test_idle,
                                        take_action_break_a,
                                        take_action_break_b,
                                        take_action_break_c,
                                        take_action_ocimem_a,
                                        take_action_ocimem_b,
                                        take_action_tracectrl,
                                        take_action_tracemem_a,
                                        take_action_tracemem_b,
                                        take_no_action_break_a,
                                        take_no_action_break_b,
                                        take_no_action_break_c,
                                        take_no_action_ocimem_a,
                                        take_no_action_tracemem_a
                                     )
;

  output  [ 37: 0] jdo;
  output           jrst_n;
  output           st_ready_test_idle;
  output           take_action_break_a;
  output           take_action_break_b;
  output           take_action_break_c;
  output           take_action_ocimem_a;
  output           take_action_ocimem_b;
  output           take_action_tracectrl;
  output           take_action_tracemem_a;
  output           take_action_tracemem_b;
  output           take_no_action_break_a;
  output           take_no_action_break_b;
  output           take_no_action_break_c;
  output           take_no_action_ocimem_a;
  output           take_no_action_tracemem_a;
  input   [ 31: 0] MonDReg;
  input   [ 31: 0] break_readreg;
  input            clk;
  input            dbrk_hit0_latch;
  input            dbrk_hit1_latch;
  input            dbrk_hit2_latch;
  input            dbrk_hit3_latch;
  input            debugack;
  input            monitor_error;
  input            monitor_ready;
  input            reset_n;
  input            resetlatch;
  input            tracemem_on;
  input   [ 35: 0] tracemem_trcdata;
  input            tracemem_tw;
  input   [  6: 0] trc_im_addr;
  input            trc_on;
  input            trc_wrap;
  input            trigbrktype;
  input            trigger_state_1;

  wire    [ 37: 0] jdo;
  wire             jrst_n;
  wire    [ 37: 0] sr;
  wire             st_ready_test_idle;
  wire             take_action_break_a;
  wire             take_action_break_b;
  wire             take_action_break_c;
  wire             take_action_ocimem_a;
  wire             take_action_ocimem_b;
  wire             take_action_tracectrl;
  wire             take_action_tracemem_a;
  wire             take_action_tracemem_b;
  wire             take_no_action_break_a;
  wire             take_no_action_break_b;
  wire             take_no_action_break_c;
  wire             take_no_action_ocimem_a;
  wire             take_no_action_tracemem_a;
  wire             vji_cdr;
  wire    [  1: 0] vji_ir_in;
  wire    [  1: 0] vji_ir_out;
  wire             vji_rti;
  wire             vji_sdr;
  wire             vji_tck;
  wire             vji_tdi;
  wire             vji_tdo;
  wire             vji_udr;
  wire             vji_uir;
  cpu_jtag_debug_module_tck the_cpu_jtag_debug_module_tck
    (
      .MonDReg            (MonDReg),
      .break_readreg      (break_readreg),
      .dbrk_hit0_latch    (dbrk_hit0_latch),
      .dbrk_hit1_latch    (dbrk_hit1_latch),
      .dbrk_hit2_latch    (dbrk_hit2_latch),
      .dbrk_hit3_latch    (dbrk_hit3_latch),
      .debugack           (debugack),
      .ir_in              (vji_ir_in),
      .ir_out             (vji_ir_out),
      .jrst_n             (jrst_n),
      .jtag_state_rti     (vji_rti),
      .monitor_error      (monitor_error),
      .monitor_ready      (monitor_ready),
      .reset_n            (reset_n),
      .resetlatch         (resetlatch),
      .sr                 (sr),
      .st_ready_test_idle (st_ready_test_idle),
      .tck                (vji_tck),
      .tdi                (vji_tdi),
      .tdo                (vji_tdo),
      .tracemem_on        (tracemem_on),
      .tracemem_trcdata   (tracemem_trcdata),
      .tracemem_tw        (tracemem_tw),
      .trc_im_addr        (trc_im_addr),
      .trc_on             (trc_on),
      .trc_wrap           (trc_wrap),
      .trigbrktype        (trigbrktype),
      .trigger_state_1    (trigger_state_1),
      .vs_cdr             (vji_cdr),
      .vs_sdr             (vji_sdr),
      .vs_uir             (vji_uir)
    );

  cpu_jtag_debug_module_sysclk the_cpu_jtag_debug_module_sysclk
    (
      .clk                       (clk),
      .ir_in                     (vji_ir_in),
      .jdo                       (jdo),
      .sr                        (sr),
      .take_action_break_a       (take_action_break_a),
      .take_action_break_b       (take_action_break_b),
      .take_action_break_c       (take_action_break_c),
      .take_action_ocimem_a      (take_action_ocimem_a),
      .take_action_ocimem_b      (take_action_ocimem_b),
      .take_action_tracectrl     (take_action_tracectrl),
      .take_action_tracemem_a    (take_action_tracemem_a),
      .take_action_tracemem_b    (take_action_tracemem_b),
      .take_no_action_break_a    (take_no_action_break_a),
      .take_no_action_break_b    (take_no_action_break_b),
      .take_no_action_break_c    (take_no_action_break_c),
      .take_no_action_ocimem_a   (take_no_action_ocimem_a),
      .take_no_action_tracemem_a (take_no_action_tracemem_a),
      .vs_udr                    (vji_udr),
      .vs_uir                    (vji_uir)
    );


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign vji_tck = 1'b0;
  assign vji_tdi = 1'b0;
  assign vji_sdr = 1'b0;
  assign vji_cdr = 1'b0;
  assign vji_rti = 1'b0;
  assign vji_uir = 1'b0;
  assign vji_udr = 1'b0;
  assign vji_ir_in = 2'b0;

//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  sld_virtual_jtag_basic cpu_jtag_debug_module_phy
//    (
//      .ir_in (vji_ir_in),
//      .ir_out (vji_ir_out),
//      .jtag_state_rti (vji_rti),
//      .tck (vji_tck),
//      .tdi (vji_tdi),
//      .tdo (vji_tdo),
//      .virtual_state_cdr (vji_cdr),
//      .virtual_state_sdr (vji_sdr),
//      .virtual_state_udr (vji_udr),
//      .virtual_state_uir (vji_uir)
//    );
//
//  defparam cpu_jtag_debug_module_phy.sld_auto_instance_index = "YES",
//           cpu_jtag_debug_module_phy.sld_instance_index = 0,
//           cpu_jtag_debug_module_phy.sld_ir_width = 2,
//           cpu_jtag_debug_module_phy.sld_mfg_id = 70,
//           cpu_jtag_debug_module_phy.sld_sim_action = "",
//           cpu_jtag_debug_module_phy.sld_sim_n_scan = 0,
//           cpu_jtag_debug_module_phy.sld_sim_total_length = 0,
//           cpu_jtag_debug_module_phy.sld_type_id = 34,
//           cpu_jtag_debug_module_phy.sld_version = 3;
//
//synthesis read_comments_as_HDL off

endmodule


/* SLline 20490 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_clock_0.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_edge_to_pulse (
                                          // inputs:
                                           clock,
                                           data_in,
                                           reset_n,

                                          // outputs:
                                           data_out
                                        )
;

  output           data_out;
  input            clock;
  input            data_in;
  input            reset_n;

  reg              data_in_d1;
  wire             data_out;
  always @(posedge clock or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  assign data_out = data_in ^ data_in_d1;

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_slave_FSM (
                                      // inputs:
                                       master_read_done_token,
                                       master_write_done_token,
                                       slave_clk,
                                       slave_read,
                                       slave_reset_n,
                                       slave_write,

                                      // outputs:
                                       slave_read_request,
                                       slave_waitrequest,
                                       slave_write_request
                                    )
;

  output           slave_read_request;
  output           slave_waitrequest;
  output           slave_write_request;
  input            master_read_done_token;
  input            master_write_done_token;
  input            slave_clk;
  input            slave_read;
  input            slave_reset_n;
  input            slave_write;

  reg              next_slave_read_request;
  reg     [  2: 0] next_slave_state;
  reg              next_slave_write_request;
  reg              slave_read_request;
  reg     [  2: 0] slave_state;
  reg              slave_waitrequest;
  reg              slave_write_request;
  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_read_request <= 0;
      else if (1)
          slave_read_request <= next_slave_read_request;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_write_request <= 0;
      else if (1)
          slave_write_request <= next_slave_write_request;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_state <= 3'b001;
      else if (1)
          slave_state <= next_slave_state;
    end


  always @(master_read_done_token or master_write_done_token or slave_read or slave_read_request or slave_state or slave_write or slave_write_request)
    begin
      case (slave_state) // synthesis parallel_case
      
          3'b001: begin
              //read request: go from IDLE state to READ_WAIT state
              if (slave_read)
                begin
                  next_slave_state = 3'b010;
                  slave_waitrequest = 1;
                  next_slave_read_request = !slave_read_request;
                  next_slave_write_request = slave_write_request;
                end
              else if (slave_write)
                begin
                  next_slave_state = 3'b100;
                  slave_waitrequest = 1;
                  next_slave_read_request = slave_read_request;
                  next_slave_write_request = !slave_write_request;
                end
              else 
                begin
                  next_slave_state = slave_state;
                  slave_waitrequest = 0;
                  next_slave_read_request = slave_read_request;
                  next_slave_write_request = slave_write_request;
                end
          end // 3'b001 
      
          3'b010: begin
              //stay in READ_WAIT state until master passes read done token
              if (master_read_done_token)
                begin
                  next_slave_state = 3'b001;
                  slave_waitrequest = 0;
                end
              else 
                begin
                  next_slave_state = 3'b010;
                  slave_waitrequest = 1;
                end
              next_slave_read_request = slave_read_request;
              next_slave_write_request = slave_write_request;
          end // 3'b010 
      
          3'b100: begin
              //stay in WRITE_WAIT state until master passes write done token
              if (master_write_done_token)
                begin
                  next_slave_state = 3'b001;
                  slave_waitrequest = 0;
                end
              else 
                begin
                  next_slave_state = 3'b100;
                  slave_waitrequest = 1;
                end
              next_slave_read_request = slave_read_request;
              next_slave_write_request = slave_write_request;
          end // 3'b100 
      
          default: begin
              next_slave_state = 3'b001;
              slave_waitrequest = 0;
              next_slave_read_request = slave_read_request;
              next_slave_write_request = slave_write_request;
          end // default
      
      endcase // slave_state
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_master_FSM (
                                       // inputs:
                                        master_clk,
                                        master_reset_n,
                                        master_waitrequest,
                                        slave_read_request_token,
                                        slave_write_request_token,

                                       // outputs:
                                        master_read,
                                        master_read_done,
                                        master_write,
                                        master_write_done
                                     )
;

  output           master_read;
  output           master_read_done;
  output           master_write;
  output           master_write_done;
  input            master_clk;
  input            master_reset_n;
  input            master_waitrequest;
  input            slave_read_request_token;
  input            slave_write_request_token;

  reg              master_read;
  reg              master_read_done;
  reg     [  2: 0] master_state;
  reg              master_write;
  reg              master_write_done;
  reg              next_master_read;
  reg              next_master_read_done;
  reg     [  2: 0] next_master_state;
  reg              next_master_write;
  reg              next_master_write_done;
  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_read_done <= 0;
      else if (1)
          master_read_done <= next_master_read_done;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_write_done <= 0;
      else if (1)
          master_write_done <= next_master_write_done;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_read <= 0;
      else if (1)
          master_read <= next_master_read;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_write <= 0;
      else if (1)
          master_write <= next_master_write;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_state <= 3'b001;
      else if (1)
          master_state <= next_master_state;
    end


  always @(master_read or master_read_done or master_state or master_waitrequest or master_write or master_write_done or slave_read_request_token or slave_write_request_token)
    begin
      case (master_state) // synthesis parallel_case
      
          3'b001: begin
              //if read request token from slave then goto READ_WAIT state
              if (slave_read_request_token)
                begin
                  next_master_state = 3'b010;
                  next_master_read = 1;
                  next_master_write = 0;
                end
              else if (slave_write_request_token)
                begin
                  next_master_state = 3'b100;
                  next_master_read = 0;
                  next_master_write = 1;
                end
              else 
                begin
                  next_master_state = master_state;
                  next_master_read = 0;
                  next_master_write = 0;
                end
              next_master_read_done = master_read_done;
              next_master_write_done = master_write_done;
          end // 3'b001 
      
          3'b010: begin
              //stay in READ_WAIT state until master wait is deasserted
              if (!master_waitrequest)
                begin
                  next_master_state = 3'b001;
                  next_master_read_done = !master_read_done;
                  next_master_read = 0;
                end
              else 
                begin
                  next_master_state = 3'b010;
                  next_master_read_done = master_read_done;
                  next_master_read = master_read;
                end
              next_master_write_done = master_write_done;
              next_master_write = 0;
          end // 3'b010 
      
          3'b100: begin
              //stay in WRITE_WAIT state until slave wait is deasserted
              if (!master_waitrequest)
                begin
                  next_master_state = 3'b001;
                  next_master_write = 0;
                  next_master_write_done = !master_write_done;
                end
              else 
                begin
                  next_master_state = 3'b100;
                  next_master_write = master_write;
                  next_master_write_done = master_write_done;
                end
              next_master_read_done = master_read_done;
              next_master_read = 0;
          end // 3'b100 
      
          default: begin
              next_master_state = 3'b001;
              next_master_write = 0;
              next_master_write_done = master_write_done;
              next_master_read = 0;
              next_master_read_done = master_read_done;
          end // default
      
      endcase // master_state
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module custom_dma_clock_0_bit_pipe (
                                     // inputs:
                                      clk1,
                                      clk2,
                                      data_in,
                                      reset_clk1_n,
                                      reset_clk2_n,

                                     // outputs:
                                      data_out
                                   )
;

  output           data_out;
  input            clk1;
  input            clk2;
  input            data_in;
  input            reset_clk1_n;
  input            reset_clk2_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-to \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  always @(posedge clk1 or negedge reset_clk1_n)
    begin
      if (reset_clk1_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk2 or negedge reset_clk2_n)
    begin
      if (reset_clk2_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//Clock Domain Crossing Adaptercustom_dma_clock_0


module custom_dma_clock_0 (
                            // inputs:
                             master_clk,
                             master_endofpacket,
                             master_readdata,
                             master_reset_n,
                             master_waitrequest,
                             slave_address,
                             slave_byteenable,
                             slave_clk,
                             slave_nativeaddress,
                             slave_read,
                             slave_reset_n,
                             slave_write,
                             slave_writedata,

                            // outputs:
                             master_address,
                             master_byteenable,
                             master_nativeaddress,
                             master_read,
                             master_write,
                             master_writedata,
                             slave_endofpacket,
                             slave_readdata,
                             slave_waitrequest
                          )
;

  output  [  3: 0] master_address;
  output  [  1: 0] master_byteenable;
  output  [  2: 0] master_nativeaddress;
  output           master_read;
  output           master_write;
  output  [ 15: 0] master_writedata;
  output           slave_endofpacket;
  output  [ 15: 0] slave_readdata;
  output           slave_waitrequest;
  input            master_clk;
  input            master_endofpacket;
  input   [ 15: 0] master_readdata;
  input            master_reset_n;
  input            master_waitrequest;
  input   [  3: 0] slave_address;
  input   [  1: 0] slave_byteenable;
  input            slave_clk;
  input   [  2: 0] slave_nativeaddress;
  input            slave_read;
  input            slave_reset_n;
  input            slave_write;
  input   [ 15: 0] slave_writedata;

  reg     [  3: 0] master_address /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  reg     [  1: 0] master_byteenable /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  reg     [  2: 0] master_nativeaddress /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  wire             master_read;
  wire             master_read_done;
  wire             master_read_done_sync;
  wire             master_read_done_token;
  wire             master_write;
  wire             master_write_done;
  wire             master_write_done_sync;
  wire             master_write_done_token;
  reg     [ 15: 0] master_writedata /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON"  */;
  reg     [  3: 0] slave_address_d1 /* synthesis ALTERA_ATTRIBUTE = "{-to \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  reg     [  1: 0] slave_byteenable_d1 /* synthesis ALTERA_ATTRIBUTE = "{-to \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  wire             slave_endofpacket;
  reg     [  2: 0] slave_nativeaddress_d1 /* synthesis ALTERA_ATTRIBUTE = "{-to \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  wire             slave_read_request;
  wire             slave_read_request_sync;
  wire             slave_read_request_token;
  reg     [ 15: 0] slave_readdata /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON"  */;
  reg     [ 15: 0] slave_readdata_p1;
  wire             slave_waitrequest;
  wire             slave_write_request;
  wire             slave_write_request_sync;
  wire             slave_write_request_token;
  reg     [ 15: 0] slave_writedata_d1 /* synthesis ALTERA_ATTRIBUTE = "{-to \"*\"} CUT=ON ; PRESERVE_REGISTER=ON"  */;
  //in, which is an e_avalon_slave
  //out, which is an e_avalon_master
  altera_std_synchronizer the_altera_std_synchronizer
    (
      .clk (slave_clk),
      .din (master_read_done),
      .dout (master_read_done_sync),
      .reset_n (slave_reset_n)
    );

  defparam the_altera_std_synchronizer.depth = 2;

  altera_std_synchronizer the_altera_std_synchronizer1
    (
      .clk (slave_clk),
      .din (master_write_done),
      .dout (master_write_done_sync),
      .reset_n (slave_reset_n)
    );

  defparam the_altera_std_synchronizer1.depth = 2;

  //read_done_edge_to_pulse, which is an e_instance
  custom_dma_clock_0_edge_to_pulse read_done_edge_to_pulse
    (
      .clock    (slave_clk),
      .data_in  (master_read_done_sync),
      .data_out (master_read_done_token),
      .reset_n  (slave_reset_n)
    );

  //write_done_edge_to_pulse, which is an e_instance
  custom_dma_clock_0_edge_to_pulse write_done_edge_to_pulse
    (
      .clock    (slave_clk),
      .data_in  (master_write_done_sync),
      .data_out (master_write_done_token),
      .reset_n  (slave_reset_n)
    );

  //slave_FSM, which is an e_instance
  custom_dma_clock_0_slave_FSM slave_FSM
    (
      .master_read_done_token  (master_read_done_token),
      .master_write_done_token (master_write_done_token),
      .slave_clk               (slave_clk),
      .slave_read              (slave_read),
      .slave_read_request      (slave_read_request),
      .slave_reset_n           (slave_reset_n),
      .slave_waitrequest       (slave_waitrequest),
      .slave_write             (slave_write),
      .slave_write_request     (slave_write_request)
    );

  altera_std_synchronizer the_altera_std_synchronizer2
    (
      .clk (master_clk),
      .din (slave_read_request),
      .dout (slave_read_request_sync),
      .reset_n (master_reset_n)
    );

  defparam the_altera_std_synchronizer2.depth = 2;

  altera_std_synchronizer the_altera_std_synchronizer3
    (
      .clk (master_clk),
      .din (slave_write_request),
      .dout (slave_write_request_sync),
      .reset_n (master_reset_n)
    );

  defparam the_altera_std_synchronizer3.depth = 2;

  //read_request_edge_to_pulse, which is an e_instance
  custom_dma_clock_0_edge_to_pulse read_request_edge_to_pulse
    (
      .clock    (master_clk),
      .data_in  (slave_read_request_sync),
      .data_out (slave_read_request_token),
      .reset_n  (master_reset_n)
    );

  //write_request_edge_to_pulse, which is an e_instance
  custom_dma_clock_0_edge_to_pulse write_request_edge_to_pulse
    (
      .clock    (master_clk),
      .data_in  (slave_write_request_sync),
      .data_out (slave_write_request_token),
      .reset_n  (master_reset_n)
    );

  //master_FSM, which is an e_instance
  custom_dma_clock_0_master_FSM master_FSM
    (
      .master_clk                (master_clk),
      .master_read               (master_read),
      .master_read_done          (master_read_done),
      .master_reset_n            (master_reset_n),
      .master_waitrequest        (master_waitrequest),
      .master_write              (master_write),
      .master_write_done         (master_write_done),
      .slave_read_request_token  (slave_read_request_token),
      .slave_write_request_token (slave_write_request_token)
    );

  //endofpacket_bit_pipe, which is an e_instance
  custom_dma_clock_0_bit_pipe endofpacket_bit_pipe
    (
      .clk1         (slave_clk),
      .clk2         (master_clk),
      .data_in      (master_endofpacket),
      .data_out     (slave_endofpacket),
      .reset_clk1_n (slave_reset_n),
      .reset_clk2_n (master_reset_n)
    );

  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          slave_readdata_p1 <= 0;
      else if (master_read & ~master_waitrequest)
          slave_readdata_p1 <= master_readdata;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_readdata <= 0;
      else 
        slave_readdata <= slave_readdata_p1;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_writedata_d1 <= 0;
      else 
        slave_writedata_d1 <= slave_writedata;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_writedata <= 0;
      else 
        master_writedata <= slave_writedata_d1;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_address_d1 <= 0;
      else 
        slave_address_d1 <= slave_address;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_address <= 0;
      else 
        master_address <= slave_address_d1;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_nativeaddress_d1 <= 0;
      else 
        slave_nativeaddress_d1 <= slave_nativeaddress;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_nativeaddress <= 0;
      else 
        master_nativeaddress <= slave_nativeaddress_d1;
    end


  always @(posedge slave_clk or negedge slave_reset_n)
    begin
      if (slave_reset_n == 0)
          slave_byteenable_d1 <= 0;
      else 
        slave_byteenable_d1 <= slave_byteenable;
    end


  always @(posedge master_clk or negedge master_reset_n)
    begin
      if (master_reset_n == 0)
          master_byteenable <= 0;
      else 
        master_byteenable <= slave_byteenable_d1;
    end



endmodule


/* SLline 20492 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_1.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: cpu/instruction_master
//adapter masters: pipeline_bridge/s1
//asp_debug: 0
//byteaddr_width: 14
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 4
//downstream_addr_shift: 2
//downstream_burstcount_width: 1
//downstream_max_burstcount: 1
//downstream_pipeline: 1
//dynamic_slave: 1
//master_always_burst_max_burst: 1
//master_burst_on_burst_boundaries_only: 0
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 1
//nativeaddr_width: 12
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 0
//upstream_burstcount: 4'h8
//upstream_burstcount_width: 4
//upstream_max_burstcount: 8
//zero_address_width: 0


module custom_dma_burst_1 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             reg_downstream_address,
                             reg_downstream_arbitrationshare,
                             reg_downstream_burstcount,
                             reg_downstream_byteenable,
                             reg_downstream_debugaccess,
                             reg_downstream_nativeaddress,
                             reg_downstream_read,
                             reg_downstream_write,
                             reg_downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 11: 0] reg_downstream_address;
  output  [  3: 0] reg_downstream_arbitrationshare;
  output           reg_downstream_burstcount;
  output  [  3: 0] reg_downstream_byteenable;
  output           reg_downstream_debugaccess;
  output  [ 11: 0] reg_downstream_nativeaddress;
  output           reg_downstream_read;
  output           reg_downstream_write;
  output  [ 31: 0] reg_downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 13: 0] upstream_address;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 11: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  2: 0] address_offset;
  reg              atomic_counter;
  wire    [  2: 0] burst_offset;
  wire    [ 13: 0] current_upstream_address;
  wire    [  3: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  3: 0] data_counter;
  wire    [  3: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 11: 0] downstream_address;
  wire    [ 13: 0] downstream_address_base;
  wire    [  3: 0] downstream_arbitrationshare;
  wire             downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 11: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire             max_burst_size;
  wire             p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  2: 0] read_address_offset;
  wire             read_update_count;
  wire    [  3: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 11: 0] reg_downstream_address;
  reg     [  3: 0] reg_downstream_arbitrationshare;
  reg              reg_downstream_burstcount;
  reg     [  3: 0] reg_downstream_byteenable;
  reg              reg_downstream_debugaccess;
  reg     [ 11: 0] reg_downstream_nativeaddress;
  reg              reg_downstream_read;
  reg              reg_downstream_write;
  reg     [ 31: 0] reg_downstream_writedata;
  reg     [  3: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 13: 0] registered_upstream_address;
  reg     [  3: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 11: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  3: 0] transactions_remaining;
  reg     [  3: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  2: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = 4'h8;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= 4'h8;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? 4'h8 : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 1;
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign downstream_arbitrationshare = current_upstream_read ? (dbs_adjusted_upstream_burstcount) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign burst_offset = downstream_address_base[4 : 2] + address_offset;
  assign downstream_address = {downstream_address_base[13 : 5],
    burst_offset,
    2'b00};

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_address <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_address <= downstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_arbitrationshare <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_arbitrationshare <= downstream_arbitrationshare;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_burstcount <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_burstcount <= downstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_byteenable <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_byteenable <= downstream_byteenable;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_debugaccess <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_debugaccess <= downstream_debugaccess;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_nativeaddress <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_nativeaddress <= downstream_nativeaddress;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_read <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_read <= downstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_write <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_write <= downstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_writedata <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_writedata <= downstream_writedata;
    end



endmodule


/* SLline 20493 "custom_dma.v" 2 */
/* SLline 1 "timestamp_timer.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module timestamp_timer (
                         // inputs:
                          address,
                          chipselect,
                          clk,
                          reset_n,
                          write_n,
                          writedata,

                         // outputs:
                          irq,
                          readdata
                       )
;

  output           irq;
  output  [ 15: 0] readdata;
  input   [  2: 0] address;
  input            chipselect;
  input            clk;
  input            reset_n;
  input            write_n;
  input   [ 15: 0] writedata;

  wire             clk_en;
  wire             control_continuous;
  wire             control_interrupt_enable;
  reg     [  3: 0] control_register;
  wire             control_wr_strobe;
  reg              counter_is_running;
  wire             counter_is_zero;
  wire    [ 31: 0] counter_load_value;
  reg     [ 31: 0] counter_snapshot;
  reg              delayed_unxcounter_is_zeroxx0;
  wire             do_start_counter;
  wire             do_stop_counter;
  reg              force_reload;
  reg     [ 31: 0] internal_counter;
  wire             irq;
  reg     [ 15: 0] period_h_register;
  wire             period_h_wr_strobe;
  reg     [ 15: 0] period_l_register;
  wire             period_l_wr_strobe;
  wire    [ 15: 0] read_mux_out;
  reg     [ 15: 0] readdata;
  wire             snap_h_wr_strobe;
  wire             snap_l_wr_strobe;
  wire    [ 31: 0] snap_read_value;
  wire             snap_strobe;
  wire             start_strobe;
  wire             status_wr_strobe;
  wire             stop_strobe;
  wire             timeout_event;
  reg              timeout_occurred;
  assign clk_en = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          internal_counter <= 32'h3E7;
      else if (counter_is_running || force_reload)
          if (counter_is_zero    || force_reload)
              internal_counter <= counter_load_value;
          else 
            internal_counter <= internal_counter - 1;
    end


  assign counter_is_zero = internal_counter == 0;
  assign counter_load_value = {period_h_register,
    period_l_register};

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          force_reload <= 0;
      else if (clk_en)
          force_reload <= period_h_wr_strobe || period_l_wr_strobe;
    end


  assign do_start_counter = start_strobe;
  assign do_stop_counter = (stop_strobe                            ) ||
    (force_reload                           ) ||
    (counter_is_zero && ~control_continuous );

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          counter_is_running <= 1'b0;
      else if (clk_en)
          if (do_start_counter)
              counter_is_running <= -1;
          else if (do_stop_counter)
              counter_is_running <= 0;
    end


  //delayed_unxcounter_is_zeroxx0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          delayed_unxcounter_is_zeroxx0 <= 0;
      else if (clk_en)
          delayed_unxcounter_is_zeroxx0 <= counter_is_zero;
    end


  assign timeout_event = (counter_is_zero) & ~(delayed_unxcounter_is_zeroxx0);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          timeout_occurred <= 0;
      else if (clk_en)
          if (status_wr_strobe)
              timeout_occurred <= 0;
          else if (timeout_event)
              timeout_occurred <= -1;
    end


  assign irq = timeout_occurred && control_interrupt_enable;
  //s1, which is an e_avalon_slave
  assign read_mux_out = ({16 {(address == 2)}} & period_l_register) |
    ({16 {(address == 3)}} & period_h_register) |
    ({16 {(address == 4)}} & snap_read_value[15 : 0]) |
    ({16 {(address == 5)}} & snap_read_value[31 : 16]) |
    ({16 {(address == 1)}} & control_register) |
    ({16 {(address == 0)}} & {counter_is_running,
    timeout_occurred});

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          readdata <= 0;
      else if (clk_en)
          readdata <= read_mux_out;
    end


  assign period_l_wr_strobe = chipselect && ~write_n && (address == 2);
  assign period_h_wr_strobe = chipselect && ~write_n && (address == 3);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          period_l_register <= 999;
      else if (period_l_wr_strobe)
          period_l_register <= writedata;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          period_h_register <= 0;
      else if (period_h_wr_strobe)
          period_h_register <= writedata;
    end


  assign snap_l_wr_strobe = chipselect && ~write_n && (address == 4);
  assign snap_h_wr_strobe = chipselect && ~write_n && (address == 5);
  assign snap_strobe = snap_l_wr_strobe || snap_h_wr_strobe;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          counter_snapshot <= 0;
      else if (snap_strobe)
          counter_snapshot <= internal_counter;
    end


  assign snap_read_value = counter_snapshot;
  assign control_wr_strobe = chipselect && ~write_n && (address == 1);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          control_register <= 0;
      else if (control_wr_strobe)
          control_register <= writedata[3 : 0];
    end


  assign stop_strobe = writedata[3] && control_wr_strobe;
  assign start_strobe = writedata[2] && control_wr_strobe;
  assign control_continuous = control_register[1];
  assign control_interrupt_enable = control_register;
  assign status_wr_strobe = chipselect && ~write_n && (address == 0);

endmodule


/* SLline 20494 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_3.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: cpu/instruction_master
//adapter masters: ddr_sdram/s1
//asp_debug: 0
//byteaddr_width: 27
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 4
//downstream_addr_shift: 2
//downstream_burstcount_width: 3
//downstream_max_burstcount: 4
//downstream_pipeline: 1
//dynamic_slave: 1
//master_always_burst_max_burst: 1
//master_burst_on_burst_boundaries_only: 0
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 1
//nativeaddr_width: 25
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 1
//upstream_burstcount: 4'h8
//upstream_burstcount_width: 4
//upstream_max_burstcount: 8
//zero_address_width: 0


module custom_dma_burst_3 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             reg_downstream_address,
                             reg_downstream_arbitrationshare,
                             reg_downstream_burstcount,
                             reg_downstream_byteenable,
                             reg_downstream_debugaccess,
                             reg_downstream_nativeaddress,
                             reg_downstream_read,
                             reg_downstream_write,
                             reg_downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 24: 0] reg_downstream_address;
  output  [  3: 0] reg_downstream_arbitrationshare;
  output  [  2: 0] reg_downstream_burstcount;
  output  [  3: 0] reg_downstream_byteenable;
  output           reg_downstream_debugaccess;
  output  [ 24: 0] reg_downstream_nativeaddress;
  output           reg_downstream_read;
  output           reg_downstream_write;
  output  [ 31: 0] reg_downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 26: 0] upstream_address;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 24: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  2: 0] address_offset;
  reg     [  2: 0] atomic_counter;
  wire    [  2: 0] burst_offset;
  wire    [ 26: 0] current_upstream_address;
  wire    [  3: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  3: 0] data_counter;
  wire    [  3: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 24: 0] downstream_address;
  wire    [ 26: 0] downstream_address_base;
  wire    [  3: 0] downstream_arbitrationshare;
  wire    [  2: 0] downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 24: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire    [  3: 0] interleave_end;
  wire    [  2: 0] max_burst_size;
  wire    [  2: 0] p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  2: 0] read_address_offset;
  wire             read_update_count;
  wire    [  3: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 24: 0] reg_downstream_address;
  reg     [  3: 0] reg_downstream_arbitrationshare;
  reg     [  2: 0] reg_downstream_burstcount;
  reg     [  3: 0] reg_downstream_byteenable;
  reg              reg_downstream_debugaccess;
  reg     [ 24: 0] reg_downstream_nativeaddress;
  reg              reg_downstream_read;
  reg              reg_downstream_write;
  reg     [ 31: 0] reg_downstream_writedata;
  reg     [  3: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 26: 0] registered_upstream_address;
  reg     [  3: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 24: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  3: 0] transactions_remaining;
  reg     [  3: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  2: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = 4'h8;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= 4'h8;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? 4'h8 : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 4 - burst_offset[1 : 0];
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign interleave_end = (dbs_adjusted_upstream_burstcount > 0) ? (dbs_adjusted_upstream_burstcount - 0) : 0;
  assign downstream_arbitrationshare = current_upstream_read ? (|burst_offset[1 : 0] + (interleave_end >> 2) + |(interleave_end[1 : 0])) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign burst_offset = downstream_address_base[4 : 2] + address_offset;
  assign downstream_address = {downstream_address_base[26 : 5],
    burst_offset,
    2'b00};

  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_address <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_address <= downstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_arbitrationshare <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_arbitrationshare <= downstream_arbitrationshare;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_burstcount <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_burstcount <= downstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_byteenable <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_byteenable <= downstream_byteenable;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_debugaccess <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_debugaccess <= downstream_debugaccess;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_nativeaddress <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_nativeaddress <= downstream_nativeaddress;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_read <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_read <= downstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_write <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_write <= downstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_writedata <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_writedata <= downstream_writedata;
    end



endmodule


/* SLline 20495 "custom_dma.v" 2 */
/* SLline 1 "custom_dma_burst_4.v" 1 */
//Legal Notice: (C)2010 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

//
//Burst adapter parameters:
//adapter is mastered by: cpu/data_master
//adapter masters: ddr_sdram/s1
//asp_debug: 0
//byteaddr_width: 27
//ceil_data_width: 32
//data_width: 32
//dbs_shift: 0
//dbs_upstream_burstcount_width: 4
//downstream_addr_shift: 2
//downstream_burstcount_width: 3
//downstream_max_burstcount: 4
//downstream_pipeline: 1
//dynamic_slave: 1
//master_always_burst_max_burst: 0
//master_burst_on_burst_boundaries_only: 1
//master_data_width: 32
//master_interleave: 0
//master_linewrap_bursts: 0
//nativeaddr_width: 25
//slave_always_burst_max_burst: 0
//slave_burst_on_burst_boundaries_only: 0
//slave_interleave: 0
//slave_linewrap_bursts: 1
//upstream_burstcount: upstream_burstcount
//upstream_burstcount_width: 4
//upstream_max_burstcount: 8
//zero_address_width: 0


module custom_dma_burst_4 (
                            // inputs:
                             clk,
                             downstream_readdata,
                             downstream_readdatavalid,
                             downstream_waitrequest,
                             reset_n,
                             upstream_address,
                             upstream_burstcount,
                             upstream_byteenable,
                             upstream_debugaccess,
                             upstream_nativeaddress,
                             upstream_read,
                             upstream_write,
                             upstream_writedata,

                            // outputs:
                             reg_downstream_address,
                             reg_downstream_arbitrationshare,
                             reg_downstream_burstcount,
                             reg_downstream_byteenable,
                             reg_downstream_debugaccess,
                             reg_downstream_nativeaddress,
                             reg_downstream_read,
                             reg_downstream_write,
                             reg_downstream_writedata,
                             upstream_readdata,
                             upstream_readdatavalid,
                             upstream_waitrequest
                          )
;

  output  [ 24: 0] reg_downstream_address;
  output  [  3: 0] reg_downstream_arbitrationshare;
  output  [  2: 0] reg_downstream_burstcount;
  output  [  3: 0] reg_downstream_byteenable;
  output           reg_downstream_debugaccess;
  output  [ 24: 0] reg_downstream_nativeaddress;
  output           reg_downstream_read;
  output           reg_downstream_write;
  output  [ 31: 0] reg_downstream_writedata;
  output  [ 31: 0] upstream_readdata;
  output           upstream_readdatavalid;
  output           upstream_waitrequest;
  input            clk;
  input   [ 31: 0] downstream_readdata;
  input            downstream_readdatavalid;
  input            downstream_waitrequest;
  input            reset_n;
  input   [ 26: 0] upstream_address;
  input   [  3: 0] upstream_burstcount;
  input   [  3: 0] upstream_byteenable;
  input            upstream_debugaccess;
  input   [ 24: 0] upstream_nativeaddress;
  input            upstream_read;
  input            upstream_write;
  input   [ 31: 0] upstream_writedata;

  wire    [  2: 0] address_offset;
  reg     [  2: 0] atomic_counter;
  wire    [ 26: 0] current_upstream_address;
  wire    [  3: 0] current_upstream_burstcount;
  wire             current_upstream_read;
  wire             current_upstream_write;
  reg     [  3: 0] data_counter;
  wire    [  3: 0] dbs_adjusted_upstream_burstcount;
  wire    [ 24: 0] downstream_address;
  wire    [ 26: 0] downstream_address_base;
  wire    [  3: 0] downstream_arbitrationshare;
  wire    [  2: 0] downstream_burstcount;
  wire             downstream_burstdone;
  wire    [  3: 0] downstream_byteenable;
  wire             downstream_debugaccess;
  wire    [ 24: 0] downstream_nativeaddress;
  reg              downstream_read;
  wire             downstream_write;
  reg              downstream_write_reg;
  wire    [ 31: 0] downstream_writedata;
  wire             enable_state_change;
  wire             fifo_empty;
  wire    [  3: 0] interleave_end;
  wire    [  2: 0] max_burst_size;
  wire    [  2: 0] p1_atomic_counter;
  wire             p1_fifo_empty;
  wire             p1_state_busy;
  wire             p1_state_idle;
  wire             pending_register_enable;
  wire             pending_upstream_read;
  reg              pending_upstream_read_reg;
  wire             pending_upstream_write;
  reg              pending_upstream_write_reg;
  reg     [  2: 0] read_address_offset;
  wire             read_update_count;
  wire    [  3: 0] read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 24: 0] reg_downstream_address;
  reg     [  3: 0] reg_downstream_arbitrationshare;
  reg     [  2: 0] reg_downstream_burstcount;
  reg     [  3: 0] reg_downstream_byteenable;
  reg              reg_downstream_debugaccess;
  reg     [ 24: 0] reg_downstream_nativeaddress;
  reg              reg_downstream_read;
  reg              reg_downstream_write;
  reg     [ 31: 0] reg_downstream_writedata;
  reg     [  3: 0] registered_read_write_dbs_adjusted_upstream_burstcount;
  reg     [ 26: 0] registered_upstream_address;
  reg     [  3: 0] registered_upstream_burstcount;
  reg     [  3: 0] registered_upstream_byteenable;
  reg     [ 24: 0] registered_upstream_nativeaddress;
  reg              registered_upstream_read;
  reg              registered_upstream_write;
  reg              state_busy;
  reg              state_idle;
  wire             sync_nativeaddress;
  wire    [  3: 0] transactions_remaining;
  reg     [  3: 0] transactions_remaining_reg;
  wire             update_count;
  wire             upstream_burstdone;
  wire             upstream_read_run;
  wire    [ 31: 0] upstream_readdata;
  wire             upstream_readdatavalid;
  wire             upstream_waitrequest;
  wire             upstream_write_run;
  reg     [  2: 0] write_address_offset;
  wire             write_update_count;
  assign sync_nativeaddress = |upstream_nativeaddress;
  //downstream, which is an e_avalon_master
  //upstream, which is an e_avalon_slave
  assign upstream_burstdone = current_upstream_read ? (transactions_remaining == downstream_burstcount) & downstream_read & ~downstream_waitrequest : (transactions_remaining == (atomic_counter + 1)) & downstream_write & ~downstream_waitrequest;
  assign p1_atomic_counter = atomic_counter + (downstream_read ? downstream_burstcount : 1);
  assign downstream_burstdone = (downstream_read | downstream_write) & ~downstream_waitrequest & (p1_atomic_counter == downstream_burstcount);
  assign dbs_adjusted_upstream_burstcount = pending_register_enable ? read_write_dbs_adjusted_upstream_burstcount : registered_read_write_dbs_adjusted_upstream_burstcount;
  assign read_write_dbs_adjusted_upstream_burstcount = upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_read_write_dbs_adjusted_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_read_write_dbs_adjusted_upstream_burstcount <= read_write_dbs_adjusted_upstream_burstcount;
    end


  assign p1_state_idle = state_idle & ~upstream_read & ~upstream_write | state_busy & (data_counter == 0) & p1_fifo_empty & ~pending_upstream_read & ~pending_upstream_write;
  assign p1_state_busy = state_idle & (upstream_read | upstream_write) | state_busy & (~(data_counter == 0) | ~p1_fifo_empty | pending_upstream_read | pending_upstream_write);
  assign enable_state_change = ~(downstream_read | downstream_write) | ~downstream_waitrequest;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_read_reg <= 0;
      else if (upstream_read & state_idle)
          pending_upstream_read_reg <= -1;
      else if (upstream_burstdone)
          pending_upstream_read_reg <= 0;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          pending_upstream_write_reg <= 0;
      else if (upstream_burstdone)
          pending_upstream_write_reg <= 0;
      else if (upstream_write & (state_idle | ~upstream_waitrequest))
          pending_upstream_write_reg <= -1;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_idle <= 1;
      else if (enable_state_change)
          state_idle <= p1_state_idle;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          state_busy <= 0;
      else if (enable_state_change)
          state_busy <= p1_state_busy;
    end


  assign pending_upstream_read = pending_upstream_read_reg;
  assign pending_upstream_write = pending_upstream_write_reg & ~upstream_burstdone;
  assign pending_register_enable = state_idle | ((upstream_read | upstream_write) & ~upstream_waitrequest);
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_read <= 0;
      else if (pending_register_enable)
          registered_upstream_read <= upstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_write <= 0;
      else if (pending_register_enable)
          registered_upstream_write <= upstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_burstcount <= 0;
      else if (pending_register_enable)
          registered_upstream_burstcount <= upstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_address <= 0;
      else if (pending_register_enable)
          registered_upstream_address <= upstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_nativeaddress <= 0;
      else if (pending_register_enable)
          registered_upstream_nativeaddress <= upstream_nativeaddress;
    end


  assign current_upstream_read = registered_upstream_read & !downstream_write;
  assign current_upstream_write = registered_upstream_write;
  assign current_upstream_address = registered_upstream_address;
  assign current_upstream_burstcount = pending_register_enable ? upstream_burstcount : registered_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          atomic_counter <= 0;
      else if ((downstream_read | downstream_write) & ~downstream_waitrequest)
          atomic_counter <= downstream_burstdone ? 0 : p1_atomic_counter;
    end


  assign read_update_count = current_upstream_read & ~downstream_waitrequest;
  assign write_update_count = current_upstream_write & downstream_write & downstream_burstdone;
  assign update_count = read_update_count | write_update_count;
  assign transactions_remaining = (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : transactions_remaining_reg;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          transactions_remaining_reg <= 0;
      else 
        transactions_remaining_reg <= (state_idle & (upstream_read | upstream_write)) ? dbs_adjusted_upstream_burstcount : update_count ? transactions_remaining_reg - downstream_burstcount : transactions_remaining_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_counter <= 0;
      else 
        data_counter <= state_idle & upstream_read & ~upstream_waitrequest ?  dbs_adjusted_upstream_burstcount : downstream_readdatavalid ? data_counter - 1 : data_counter;
    end


  assign max_burst_size = 4;
  assign downstream_burstcount = (transactions_remaining > max_burst_size) ? max_burst_size : transactions_remaining;
  assign interleave_end = (dbs_adjusted_upstream_burstcount > 0) ? (dbs_adjusted_upstream_burstcount - 0) : 0;
  assign downstream_arbitrationshare = current_upstream_read ? (0 + (interleave_end >> 2) + |(interleave_end[1 : 0])) : dbs_adjusted_upstream_burstcount;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_address_offset <= 0;
      else 
        write_address_offset <= state_idle & upstream_write ? 0 : ((downstream_write & ~downstream_waitrequest & downstream_burstdone)) ? write_address_offset + downstream_burstcount : write_address_offset;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_address_offset <= 0;
      else 
        read_address_offset <= state_idle & upstream_read ? 0 : (downstream_read & ~downstream_waitrequest) ? read_address_offset + downstream_burstcount : read_address_offset;
    end


  assign downstream_nativeaddress = registered_upstream_nativeaddress >> 2;
  assign address_offset = current_upstream_read ? read_address_offset : write_address_offset;
  assign downstream_address_base = current_upstream_address;
  assign downstream_address = downstream_address_base + {address_offset, 2'b00};
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_read <= 0;
      else if (~downstream_read | ~downstream_waitrequest)
          downstream_read <= state_idle & upstream_read ? 1 : (transactions_remaining == downstream_burstcount) ? 0 : downstream_read;
    end


  assign upstream_readdatavalid = downstream_readdatavalid;
  assign upstream_readdata = downstream_readdata;
  assign fifo_empty = 1;
  assign p1_fifo_empty = 1;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          downstream_write_reg <= 0;
      else if (~downstream_write_reg | ~downstream_waitrequest)
          downstream_write_reg <= state_idle & upstream_write ? 1 : ((transactions_remaining == downstream_burstcount) & downstream_burstdone) ? 0 : downstream_write_reg;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          registered_upstream_byteenable <= 4'b1111;
      else if (pending_register_enable)
          registered_upstream_byteenable <= upstream_byteenable;
    end


  assign downstream_write = downstream_write_reg & upstream_write & !downstream_read;
  assign downstream_byteenable = downstream_write_reg ? upstream_byteenable : registered_upstream_byteenable;
  assign downstream_writedata = upstream_writedata;
  assign upstream_read_run = state_idle & upstream_read;
  assign upstream_write_run = state_busy & upstream_write & ~downstream_waitrequest & !downstream_read;
  assign upstream_waitrequest = (upstream_read | current_upstream_read) ? ~upstream_read_run : current_upstream_write ? ~upstream_write_run : 1;
  assign downstream_debugaccess = upstream_debugaccess;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_address <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_address <= downstream_address;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_arbitrationshare <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_arbitrationshare <= downstream_arbitrationshare;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_burstcount <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_burstcount <= downstream_burstcount;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_byteenable <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_byteenable <= downstream_byteenable;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_debugaccess <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_debugaccess <= downstream_debugaccess;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_nativeaddress <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_nativeaddress <= downstream_nativeaddress;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_read <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_read <= downstream_read;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_write <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_write <= downstream_write;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          reg_downstream_writedata <= 0;
      else if (~downstream_waitrequest)
          reg_downstream_writedata <= downstream_writedata;
    end



endmodule


/* SLline 20496 "custom_dma.v" 2 */

`timescale 1ns / 1ps

module test_bench 
;


  wire             adsc_n_to_the_ext_ssram;
  wire    [  3: 0] bw_n_to_the_ext_ssram;
  wire             bwe_n_to_the_ext_ssram;
  wire             chipenable1_n_to_the_ext_ssram;
  wire             clk;
  wire             clk_to_sdram_from_the_ddr_sdram;
  wire             clk_to_sdram_n_from_the_ddr_sdram;
  wire             custom_dma_burst_0_downstream_debugaccess;
  wire    [ 20: 0] custom_dma_burst_0_downstream_nativeaddress;
  wire    [ 31: 0] custom_dma_burst_1_upstream_writedata;
  wire             custom_dma_burst_3_downstream_debugaccess;
  wire    [ 24: 0] custom_dma_burst_3_downstream_nativeaddress;
  wire    [ 31: 0] custom_dma_burst_3_upstream_writedata;
  wire             custom_dma_burst_4_downstream_debugaccess;
  wire    [ 24: 0] custom_dma_burst_4_downstream_nativeaddress;
  wire             custom_dma_burst_5_downstream_debugaccess;
  wire    [ 24: 0] custom_dma_burst_5_downstream_nativeaddress;
  wire    [ 31: 0] custom_dma_burst_5_upstream_readdata_from_sa;
  wire             custom_dma_burst_5_upstream_readdatavalid_from_sa;
  wire             custom_dma_clock_0_out_endofpacket;
  wire    [ 12: 0] ddr_a_from_the_ddr_sdram;
  wire    [  1: 0] ddr_ba_from_the_ddr_sdram;
  wire             ddr_cas_n_from_the_ddr_sdram;
  wire             ddr_cke_from_the_ddr_sdram;
  wire             ddr_cs_n_from_the_ddr_sdram;
  wire    [  1: 0] ddr_dm_from_the_ddr_sdram;
  wire    [ 15: 0] ddr_dq_to_and_from_the_ddr_sdram;
  wire    [  1: 0] ddr_dqs_to_and_from_the_ddr_sdram;
  wire             ddr_ras_n_from_the_ddr_sdram;
  wire             ddr_we_n_from_the_ddr_sdram;
  wire    [  5: 0] dqs_delay_ctrl_to_the_ddr_sdram;
  wire             dqsupdate_to_the_ddr_sdram;
  wire    [ 20: 0] ext_ssram_bus_address;
  wire    [ 31: 0] ext_ssram_bus_data;
  reg              external_clk;
  wire             jtag_uart_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_avalon_jtag_slave_readyfordata_from_sa;
  wire             outputenable_n_to_the_ext_ssram;
  wire             pipeline_bridge_s1_endofpacket_from_sa;
  reg              reset_n;
  wire             sdram_write_clk;
  wire             ssram_clk;
  wire             stratix_dll_control_from_the_ddr_sdram;
  wire             system_clk;
  wire             write_clk_to_the_ddr_sdram;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  custom_dma DUT
    (
      .adsc_n_to_the_ext_ssram                (adsc_n_to_the_ext_ssram),
      .bw_n_to_the_ext_ssram                  (bw_n_to_the_ext_ssram),
      .bwe_n_to_the_ext_ssram                 (bwe_n_to_the_ext_ssram),
      .chipenable1_n_to_the_ext_ssram         (chipenable1_n_to_the_ext_ssram),
      .clk_to_sdram_from_the_ddr_sdram        (clk_to_sdram_from_the_ddr_sdram),
      .clk_to_sdram_n_from_the_ddr_sdram      (clk_to_sdram_n_from_the_ddr_sdram),
      .ddr_a_from_the_ddr_sdram               (ddr_a_from_the_ddr_sdram),
      .ddr_ba_from_the_ddr_sdram              (ddr_ba_from_the_ddr_sdram),
      .ddr_cas_n_from_the_ddr_sdram           (ddr_cas_n_from_the_ddr_sdram),
      .ddr_cke_from_the_ddr_sdram             (ddr_cke_from_the_ddr_sdram),
      .ddr_cs_n_from_the_ddr_sdram            (ddr_cs_n_from_the_ddr_sdram),
      .ddr_dm_from_the_ddr_sdram              (ddr_dm_from_the_ddr_sdram),
      .ddr_dq_to_and_from_the_ddr_sdram       (ddr_dq_to_and_from_the_ddr_sdram),
      .ddr_dqs_to_and_from_the_ddr_sdram      (ddr_dqs_to_and_from_the_ddr_sdram),
      .ddr_ras_n_from_the_ddr_sdram           (ddr_ras_n_from_the_ddr_sdram),
      .ddr_we_n_from_the_ddr_sdram            (ddr_we_n_from_the_ddr_sdram),
      .dqs_delay_ctrl_to_the_ddr_sdram        (dqs_delay_ctrl_to_the_ddr_sdram),
      .dqsupdate_to_the_ddr_sdram             (dqsupdate_to_the_ddr_sdram),
      .ext_ssram_bus_address                  (ext_ssram_bus_address),
      .ext_ssram_bus_data                     (ext_ssram_bus_data),
      .external_clk                           (external_clk),
      .outputenable_n_to_the_ext_ssram        (outputenable_n_to_the_ext_ssram),
      .reset_n                                (reset_n),
      .sdram_write_clk                        (sdram_write_clk),
      .ssram_clk                              (ssram_clk),
      .stratix_dll_control_from_the_ddr_sdram (stratix_dll_control_from_the_ddr_sdram),
      .system_clk                             (system_clk),
      .write_clk_to_the_ddr_sdram             (write_clk_to_the_ddr_sdram)
    );

  ext_ssram the_ext_ssram
    (
      .address        (ext_ssram_bus_address[20 : 2]),
      .adsc_n         (adsc_n_to_the_ext_ssram),
      .bw_n           (bw_n_to_the_ext_ssram),
      .bwe_n          (bwe_n_to_the_ext_ssram),
      .chipenable1_n  (chipenable1_n_to_the_ext_ssram),
      .clk            (system_clk),
      .data           (ext_ssram_bus_data),
      .outputenable_n (outputenable_n_to_the_ext_ssram),
      .reset_n        (reset_n)
    );

  ddr_sdram_test_component the_ddr_sdram_test_component
    (
      .clk       (system_clk),
      .ddr_a     (ddr_a_from_the_ddr_sdram),
      .ddr_ba    (ddr_ba_from_the_ddr_sdram),
      .ddr_cas_n (ddr_cas_n_from_the_ddr_sdram),
      .ddr_cke   (ddr_cke_from_the_ddr_sdram),
      .ddr_cs_n  (ddr_cs_n_from_the_ddr_sdram),
      .ddr_dm    (ddr_dm_from_the_ddr_sdram),
      .ddr_dq    (ddr_dq_to_and_from_the_ddr_sdram),
      .ddr_dqs   (ddr_dqs_to_and_from_the_ddr_sdram),
      .ddr_ras_n (ddr_ras_n_from_the_ddr_sdram),
      .ddr_we_n  (ddr_we_n_from_the_ddr_sdram)
    );

  initial
    external_clk = 1'b0;
  always
    #10 external_clk <= ~external_clk;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end

endmodule


//synthesis translate_on