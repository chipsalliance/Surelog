/*
:name: desc_test_12
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`ifdef DEBUGGER
`MACRO(stuff, morestuff)
`SCHMACRO()
`endif
