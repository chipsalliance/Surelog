/*
:name: class_member_test_20
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subr(ducktype #(3) x);
endclass