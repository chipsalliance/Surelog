/*
:name: class_test_61
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
`ifndef DEBUGGER
`endif
endclass