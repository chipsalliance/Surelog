// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: behavior_of_randomization_methods_0
:description: static random variables test
:tags: 18.6.3
*/

class a;
    static rand int b;
    constraint c { b > 5; b < 12; }
endclass
