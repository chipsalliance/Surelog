/*
:name: system-functions
:description: Calling system functions
:tags: 5.6.3
*/
module systemfn();
  /* Note:
   * This does not test all the individual system calls.
   * It just verifies if the concept exists using one of the
   * calls.
   */

  initial $display("hello world");
endmodule
