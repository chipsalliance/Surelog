/*
:name: string-basic
:description: Basic string example
:should_fail: 0
:tags: 5.9 5.3
*/
module top();

  initial begin;
    $display("one line");
  end

endmodule
