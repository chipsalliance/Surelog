`pragma pragma_number_other a = 123, b = 4


module top();
   wire context;

 enmodule
   
