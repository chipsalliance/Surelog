// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: string_atoreal
:description: string.atoreal()  tests
:tags: 6.16.10
*/
module top();
	string a = "4.76";
	real b = a.atoreal();
endmodule
