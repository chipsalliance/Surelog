module t;
    event e;
endmodule

