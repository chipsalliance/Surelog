/*
:name: class_member_test_49
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
virtual splinterface grinterface, winterface;
virtual interface foo_if bar_if, baz_if;
endclass