module SIM();
   initial begin
      #1 ;
      
   end
endmodule // OR
