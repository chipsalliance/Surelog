/*
:name: string_atohex
:description: string.atohex()  tests
:tags: 6.16.9
*/
module top();
	string a = "0xff";
	int b = a.atohex();
endmodule
