module MODULE_NAME_DOES_NOT_MATCH_FILE_NAME();
endmodule
