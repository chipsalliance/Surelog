/*
:name: 22.7--timescale-basic-4
:description: Test
:should_fail_because: only integers 1, 10 and 100 are allowed in this type of expression
:tags: 22.7
:type: simulation
*/
`timescale 1 ns / 1000 ps
