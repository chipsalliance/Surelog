/*
:name: 22.10--celldefine-invalid
:description: Test
:should_fail: 1
:tags: 22.10
:type: preprocessing
*/
`celldefine foo
