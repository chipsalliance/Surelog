module top;
  task simutil_memload;
    input string file;
    input int files  [1:0] ;
    input [1:0]  implic;
  endtask
endmodule // top
