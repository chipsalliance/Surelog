module test(output var a, input b);
    always_comb a = b;
endmodule
