module InoutConnect(
                    .X1(internal), 
                    .X2(internal)
                    );
   inout internal;
endmodule 
