/*
:name: string_toupper
:description: string.toupper()  tests
:should_fail: 0
:tags: 6.16.4
*/
module top();
	string a = "Test";
	string b = a.toupper();
endmodule
