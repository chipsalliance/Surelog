module mylib();
endmodule
