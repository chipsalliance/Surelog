module dut (b);                                                                                          
        wire a = 0;      
        output reg b = 0;                                                                        
        
   assign c = a;
                                                                                           
endmodule
