module top();

function automatic logic
bsg_mul_booth(
  [2:0] sdn);
  return 1;
endfunction

endmodule
