/*
:name: macromodule_definition
:description: macromodule definition test
:should_fail: 0
:tags: 23.2
*/
macromodule top();

endmodule
