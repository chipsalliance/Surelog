/*
:name: iface_class_test_2
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic #(int N = 8, type T = string);
endclass