/*
:name: net_decl_assignment
:description: net declaration assignment test
:tags: 10.3.1
*/
module top(input a, input b);

wire w = a & b;

endmodule
