/*
:name: parameter_real
:description: parameter with real value test
:should_fail: 0
:tags: 6.20.2
*/
module top();
	parameter p = 4.76;
endmodule
