/*
:name: class_test_11
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo #(int N, int P);
endclass