/*
:name: localparam
:description: localparam tests
:should_fail: 0
:tags: 6.20.4
*/
module top();
	localparam p = 123;
endmodule
