/*
:name: associative-arrays-integral
:description: Test associative arrays support
:should_fail: 0
:tags: 7.8.4 7.8
*/
module top ();

int arr [ integer ];

endmodule
