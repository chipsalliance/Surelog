// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: logic_vector
:description: logic vector tests
:tags: 6.9.1
*/
module top();
	logic [15:0] a;
endmodule
