/*
:name: class_test_23
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo implements Bar; endclass