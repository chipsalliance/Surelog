/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s001
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 15762
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_pi_4g_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_pi_4g_wphy_pi_4g_outdrv, View -
//schematic
// LAST TIME SAVED: Sep 18 06:30:05 2020
// NETLIST TIME: Oct 28 22:02:33 2020
`timescale 1ps / 1ps 




 

module wphy_pi_4g_wphy_pi_4g_outdrv (outn, outp, vdda, vss, inn, inp, tiehi, 
    tielo);

output  outn, outp;

inout  vdda, vss;

input  inn, inp, tiehi, tielo;


wphy_pi_4g_INV_D2_GL16_RVT INV0_1 ( .in(n1), .vss(vss), .out(net014), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV0_0 ( .in(n1), .vss(vss), .out(net014), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV2_1 ( .in(p1), .vss(vss), .out(net013), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV2_0 ( .in(p1), .vss(vss), .out(net013), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_3 ( .in(net013), .vss(vss), .out(outp), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_2 ( .in(net013), .vss(vss), .out(outp), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_1 ( .in(net013), .vss(vss), .out(outp), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_0 ( .in(net013), .vss(vss), .out(outp), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV3_1 ( .in(inn), .vss(vss), .out(p1), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV3_0 ( .in(inn), .vss(vss), .out(p1), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV1_1 ( .in(inp), .vss(vss), .out(n1), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV1_0 ( .in(inp), .vss(vss), .out(n1), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_3 ( .in(net014), .vss(vss), .out(outn), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_2 ( .in(net014), .vss(vss), .out(outn), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_1 ( .in(net014), .vss(vss), .out(outn), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_0 ( .in(net014), .vss(vss), .out(outn), 
    .vdd(vdda));

wphy_pi_4g_INV_D1_GL16_RVT_Mmod_nomodel INV5 ( .tiehi(tiehi), .tielo(tielo), 
    .in(net014), .vss(vss), .out(net013), .vdd(vdda));

wphy_pi_4g_INV_D1_GL16_RVT_Mmod_nomodel INV4 ( .tiehi(tiehi), .tielo(tielo), 
    .in(net013), .vss(vss), .out(net014), .vdd(vdda));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_pi_4g_wphy_pi_logic, View -
//schematic
// LAST TIME SAVED: Sep 18 06:51:38 2020
// NETLIST TIME: Oct 28 22:02:33 2020
`timescale 1ps / 1ps 




 

module wphy_pi_4g_wphy_pi_logic (en_int, enb_int, gear_out, gear_outb, sel0, 
    sel0b, sel90, sel90b, sel180, sel180b, sel270, sel270b, xcpl, 
    xcplb, vdda, vss, code, en, gear, quad, tiehi, tielo, xcpl_in);

output  en_int, enb_int;

inout  vdda, vss;

input  en, tiehi, tielo;

output [15:0]  sel270;
output [15:0]  sel270b;
output [3:0]  xcpl;
output [3:0]  gear_out;
output [3:0]  xcplb;
output [3:0]  gear_outb;
output [15:0]  sel180b;
output [15:0]  sel0b;
output [15:0]  sel180;
output [15:0]  sel90;
output [15:0]  sel90b;
output [15:0]  sel0;

input [3:0]  gear;
input [1:0]  quad;
input [15:0]  code;
input [3:0]  xcpl_in;

// Buses in the design

wire  [1:0]  quadb;

wire  [1:0]  quada;


wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_15 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[15]), 
    .vss(vss), .vdd(vdda), .b(code[15]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_14 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[14]), 
    .vss(vss), .vdd(vdda), .b(code[14]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_13 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[13]), 
    .vss(vss), .vdd(vdda), .b(code[13]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_12 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[12]), 
    .vss(vss), .vdd(vdda), .b(code[12]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_11 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[11]), 
    .vss(vss), .vdd(vdda), .b(code[11]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_10 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[10]), 
    .vss(vss), .vdd(vdda), .b(code[10]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_9 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[9]), 
    .vss(vss), .vdd(vdda), .b(code[9]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_8 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[8]), 
    .vss(vss), .vdd(vdda), .b(code[8]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_7 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[7]), 
    .vss(vss), .vdd(vdda), .b(code[7]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_6 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[6]), 
    .vss(vss), .vdd(vdda), .b(code[6]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_5 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[5]), 
    .vss(vss), .vdd(vdda), .b(code[5]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_4 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[4]), 
    .vss(vss), .vdd(vdda), .b(code[4]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_3 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[3]), 
    .vss(vss), .vdd(vdda), .b(code[3]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_2 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[2]), 
    .vss(vss), .vdd(vdda), .b(code[2]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_1 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[1]), 
    .vss(vss), .vdd(vdda), .b(code[1]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR0_0 ( .tielo(tielo), .tiehi(tiehi), .y(sel90[0]), 
    .vss(vss), .vdd(vdda), .b(code[0]), .a(quada[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_15 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[15]), .vss(vss), .vdd(vdda), .b(code[15]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_14 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[14]), .vss(vss), .vdd(vdda), .b(code[14]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_13 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[13]), .vss(vss), .vdd(vdda), .b(code[13]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_12 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[12]), .vss(vss), .vdd(vdda), .b(code[12]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_11 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[11]), .vss(vss), .vdd(vdda), .b(code[11]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_10 ( .tielo(tielo), .tiehi(tiehi), 
    .y(sel270[10]), .vss(vss), .vdd(vdda), .b(code[10]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_9 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[9]), 
    .vss(vss), .vdd(vdda), .b(code[9]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_8 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[8]), 
    .vss(vss), .vdd(vdda), .b(code[8]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_7 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[7]), 
    .vss(vss), .vdd(vdda), .b(code[7]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_6 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[6]), 
    .vss(vss), .vdd(vdda), .b(code[6]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_5 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[5]), 
    .vss(vss), .vdd(vdda), .b(code[5]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_4 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[4]), 
    .vss(vss), .vdd(vdda), .b(code[4]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_3 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[3]), 
    .vss(vss), .vdd(vdda), .b(code[3]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_2 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[2]), 
    .vss(vss), .vdd(vdda), .b(code[2]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_1 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[1]), 
    .vss(vss), .vdd(vdda), .b(code[1]), .a(quadb[0]));

wphy_pi_4g_NOR2_D1_GL16_RVT NOR1_0 ( .tielo(tielo), .tiehi(tiehi), .y(sel270[0]), 
    .vss(vss), .vdd(vdda), .b(code[0]), .a(quadb[0]));

wphy_pi_4g_INV_D2_GL16_RVT INV3 ( .in(enb_int), .vss(vss), .out(en_int), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV1_1 ( .in(quadb[1]), .vss(vss), .out(quada[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV1_0 ( .in(quadb[0]), .vss(vss), .out(quada[0]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV10_3 ( .in(gear_outb[3]), .vss(vss), 
    .out(gear_out[3]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV10_2 ( .in(gear_outb[2]), .vss(vss), 
    .out(gear_out[2]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV10_1 ( .in(gear_outb[1]), .vss(vss), 
    .out(gear_out[1]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV10_0 ( .in(gear_outb[0]), .vss(vss), 
    .out(gear_out[0]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV2 ( .in(en), .vss(vss), .out(enb_int), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_15 ( .in(sel0b[15]), .vss(vss), .out(sel0[15]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_14 ( .in(sel0b[14]), .vss(vss), .out(sel0[14]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_13 ( .in(sel0b[13]), .vss(vss), .out(sel0[13]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_12 ( .in(sel0b[12]), .vss(vss), .out(sel0[12]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_11 ( .in(sel0b[11]), .vss(vss), .out(sel0[11]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_10 ( .in(sel0b[10]), .vss(vss), .out(sel0[10]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_9 ( .in(sel0b[9]), .vss(vss), .out(sel0[9]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_8 ( .in(sel0b[8]), .vss(vss), .out(sel0[8]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_7 ( .in(sel0b[7]), .vss(vss), .out(sel0[7]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_6 ( .in(sel0b[6]), .vss(vss), .out(sel0[6]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_5 ( .in(sel0b[5]), .vss(vss), .out(sel0[5]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_4 ( .in(sel0b[4]), .vss(vss), .out(sel0[4]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_3 ( .in(sel0b[3]), .vss(vss), .out(sel0[3]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_2 ( .in(sel0b[2]), .vss(vss), .out(sel0[2]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_1 ( .in(sel0b[1]), .vss(vss), .out(sel0[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV4_0 ( .in(sel0b[0]), .vss(vss), .out(sel0[0]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_15 ( .in(sel90[15]), .vss(vss), .out(sel90b[15]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_14 ( .in(sel90[14]), .vss(vss), .out(sel90b[14]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_13 ( .in(sel90[13]), .vss(vss), .out(sel90b[13]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_12 ( .in(sel90[12]), .vss(vss), .out(sel90b[12]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_11 ( .in(sel90[11]), .vss(vss), .out(sel90b[11]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_10 ( .in(sel90[10]), .vss(vss), .out(sel90b[10]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_9 ( .in(sel90[9]), .vss(vss), .out(sel90b[9]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_8 ( .in(sel90[8]), .vss(vss), .out(sel90b[8]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_7 ( .in(sel90[7]), .vss(vss), .out(sel90b[7]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_6 ( .in(sel90[6]), .vss(vss), .out(sel90b[6]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_5 ( .in(sel90[5]), .vss(vss), .out(sel90b[5]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_4 ( .in(sel90[4]), .vss(vss), .out(sel90b[4]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_3 ( .in(sel90[3]), .vss(vss), .out(sel90b[3]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_2 ( .in(sel90[2]), .vss(vss), .out(sel90b[2]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_1 ( .in(sel90[1]), .vss(vss), .out(sel90b[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV5_0 ( .in(sel90[0]), .vss(vss), .out(sel90b[0]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV8_3 ( .in(xcplb[3]), .vss(vss), .out(xcpl[3]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV8_2 ( .in(xcplb[2]), .vss(vss), .out(xcpl[2]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV8_1 ( .in(xcplb[1]), .vss(vss), .out(xcpl[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV8_0 ( .in(xcplb[0]), .vss(vss), .out(xcpl[0]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_15 ( .in(sel180b[15]), .vss(vss), 
    .out(sel180[15]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_14 ( .in(sel180b[14]), .vss(vss), 
    .out(sel180[14]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_13 ( .in(sel180b[13]), .vss(vss), 
    .out(sel180[13]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_12 ( .in(sel180b[12]), .vss(vss), 
    .out(sel180[12]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_11 ( .in(sel180b[11]), .vss(vss), 
    .out(sel180[11]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_10 ( .in(sel180b[10]), .vss(vss), 
    .out(sel180[10]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_9 ( .in(sel180b[9]), .vss(vss), .out(sel180[9]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_8 ( .in(sel180b[8]), .vss(vss), .out(sel180[8]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_7 ( .in(sel180b[7]), .vss(vss), .out(sel180[7]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_6 ( .in(sel180b[6]), .vss(vss), .out(sel180[6]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_5 ( .in(sel180b[5]), .vss(vss), .out(sel180[5]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_4 ( .in(sel180b[4]), .vss(vss), .out(sel180[4]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_3 ( .in(sel180b[3]), .vss(vss), .out(sel180[3]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_2 ( .in(sel180b[2]), .vss(vss), .out(sel180[2]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_1 ( .in(sel180b[1]), .vss(vss), .out(sel180[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV6_0 ( .in(sel180b[0]), .vss(vss), .out(sel180[0]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_15 ( .in(sel270[15]), .vss(vss), 
    .out(sel270b[15]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_14 ( .in(sel270[14]), .vss(vss), 
    .out(sel270b[14]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_13 ( .in(sel270[13]), .vss(vss), 
    .out(sel270b[13]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_12 ( .in(sel270[12]), .vss(vss), 
    .out(sel270b[12]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_11 ( .in(sel270[11]), .vss(vss), 
    .out(sel270b[11]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_10 ( .in(sel270[10]), .vss(vss), 
    .out(sel270b[10]), .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_9 ( .in(sel270[9]), .vss(vss), .out(sel270b[9]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_8 ( .in(sel270[8]), .vss(vss), .out(sel270b[8]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_7 ( .in(sel270[7]), .vss(vss), .out(sel270b[7]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_6 ( .in(sel270[6]), .vss(vss), .out(sel270b[6]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_5 ( .in(sel270[5]), .vss(vss), .out(sel270b[5]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_4 ( .in(sel270[4]), .vss(vss), .out(sel270b[4]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_3 ( .in(sel270[3]), .vss(vss), .out(sel270b[3]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_2 ( .in(sel270[2]), .vss(vss), .out(sel270b[2]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_1 ( .in(sel270[1]), .vss(vss), .out(sel270b[1]), 
    .vdd(vdda));

wphy_pi_4g_INV_D2_GL16_RVT INV7_0 ( .in(sel270[0]), .vss(vss), .out(sel270b[0]), 
    .vdd(vdda));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND7_3 ( .tielo(tielo), .vdd(vdda), .y(xcplb[3]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(xcpl_in[3]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND7_2 ( .tielo(tielo), .vdd(vdda), .y(xcplb[2]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(xcpl_in[2]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND7_1 ( .tielo(tielo), .vdd(vdda), .y(xcplb[1]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(xcpl_in[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND7_0 ( .tielo(tielo), .vdd(vdda), .y(xcplb[0]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(xcpl_in[0]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_15 ( .tielo(tielo), .vdd(vdda), .y(sel0b[15]), 
    .vss(vss), .tiehi(tiehi), .b(code[15]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_14 ( .tielo(tielo), .vdd(vdda), .y(sel0b[14]), 
    .vss(vss), .tiehi(tiehi), .b(code[14]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_13 ( .tielo(tielo), .vdd(vdda), .y(sel0b[13]), 
    .vss(vss), .tiehi(tiehi), .b(code[13]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_12 ( .tielo(tielo), .vdd(vdda), .y(sel0b[12]), 
    .vss(vss), .tiehi(tiehi), .b(code[12]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_11 ( .tielo(tielo), .vdd(vdda), .y(sel0b[11]), 
    .vss(vss), .tiehi(tiehi), .b(code[11]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_10 ( .tielo(tielo), .vdd(vdda), .y(sel0b[10]), 
    .vss(vss), .tiehi(tiehi), .b(code[10]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_9 ( .tielo(tielo), .vdd(vdda), .y(sel0b[9]), 
    .vss(vss), .tiehi(tiehi), .b(code[9]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_8 ( .tielo(tielo), .vdd(vdda), .y(sel0b[8]), 
    .vss(vss), .tiehi(tiehi), .b(code[8]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_7 ( .tielo(tielo), .vdd(vdda), .y(sel0b[7]), 
    .vss(vss), .tiehi(tiehi), .b(code[7]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_6 ( .tielo(tielo), .vdd(vdda), .y(sel0b[6]), 
    .vss(vss), .tiehi(tiehi), .b(code[6]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_5 ( .tielo(tielo), .vdd(vdda), .y(sel0b[5]), 
    .vss(vss), .tiehi(tiehi), .b(code[5]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_4 ( .tielo(tielo), .vdd(vdda), .y(sel0b[4]), 
    .vss(vss), .tiehi(tiehi), .b(code[4]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_3 ( .tielo(tielo), .vdd(vdda), .y(sel0b[3]), 
    .vss(vss), .tiehi(tiehi), .b(code[3]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_2 ( .tielo(tielo), .vdd(vdda), .y(sel0b[2]), 
    .vss(vss), .tiehi(tiehi), .b(code[2]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_1 ( .tielo(tielo), .vdd(vdda), .y(sel0b[1]), 
    .vss(vss), .tiehi(tiehi), .b(code[1]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND0_0 ( .tielo(tielo), .vdd(vdda), .y(sel0b[0]), 
    .vss(vss), .tiehi(tiehi), .b(code[0]), .a(quadb[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND2_1 ( .tielo(tielo), .vdd(vdda), .y(quadb[1]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(quad[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND2_0 ( .tielo(tielo), .vdd(vdda), .y(quadb[0]), 
    .vss(vss), .tiehi(tiehi), .b(en), .a(quad[0]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_15 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[15]), .vss(vss), .tiehi(tiehi), .b(code[15]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_14 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[14]), .vss(vss), .tiehi(tiehi), .b(code[14]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_13 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[13]), .vss(vss), .tiehi(tiehi), .b(code[13]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_12 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[12]), .vss(vss), .tiehi(tiehi), .b(code[12]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_11 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[11]), .vss(vss), .tiehi(tiehi), .b(code[11]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_10 ( .tielo(tielo), .vdd(vdda), 
    .y(sel180b[10]), .vss(vss), .tiehi(tiehi), .b(code[10]), 
    .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_9 ( .tielo(tielo), .vdd(vdda), .y(sel180b[9]), 
    .vss(vss), .tiehi(tiehi), .b(code[9]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_8 ( .tielo(tielo), .vdd(vdda), .y(sel180b[8]), 
    .vss(vss), .tiehi(tiehi), .b(code[8]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_7 ( .tielo(tielo), .vdd(vdda), .y(sel180b[7]), 
    .vss(vss), .tiehi(tiehi), .b(code[7]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_6 ( .tielo(tielo), .vdd(vdda), .y(sel180b[6]), 
    .vss(vss), .tiehi(tiehi), .b(code[6]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_5 ( .tielo(tielo), .vdd(vdda), .y(sel180b[5]), 
    .vss(vss), .tiehi(tiehi), .b(code[5]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_4 ( .tielo(tielo), .vdd(vdda), .y(sel180b[4]), 
    .vss(vss), .tiehi(tiehi), .b(code[4]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_3 ( .tielo(tielo), .vdd(vdda), .y(sel180b[3]), 
    .vss(vss), .tiehi(tiehi), .b(code[3]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_2 ( .tielo(tielo), .vdd(vdda), .y(sel180b[2]), 
    .vss(vss), .tiehi(tiehi), .b(code[2]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_1 ( .tielo(tielo), .vdd(vdda), .y(sel180b[1]), 
    .vss(vss), .tiehi(tiehi), .b(code[1]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND5_0 ( .tielo(tielo), .vdd(vdda), .y(sel180b[0]), 
    .vss(vss), .tiehi(tiehi), .b(code[0]), .a(quada[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND1_3 ( .tielo(tielo), .vdd(vdda), 
    .y(gear_outb[3]), .vss(vss), .tiehi(tiehi), .b(en), .a(gear[3]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND1_2 ( .tielo(tielo), .vdd(vdda), 
    .y(gear_outb[2]), .vss(vss), .tiehi(tiehi), .b(en), .a(gear[2]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND1_1 ( .tielo(tielo), .vdd(vdda), 
    .y(gear_outb[1]), .vss(vss), .tiehi(tiehi), .b(en), .a(gear[1]));

wphy_pi_4g_NAND2_D1_GL16_RVT NAND1_0 ( .tielo(tielo), .vdd(vdda), 
    .y(gear_outb[0]), .vss(vss), .tiehi(tiehi), .b(en), .a(gear[0]));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_pi_4g_wphy_pi_4g_predrv, View -
//schematic
// LAST TIME SAVED: Sep 18 06:30:31 2020
// NETLIST TIME: Oct 28 22:02:33 2020
`timescale 1ps / 1ps 




 

module wphy_pi_4g_wphy_pi_4g_predrv (outn, outp, vdda, vss, en, enb, gear, gearb, 
    inn, inp);

output  outn, outp;

inout  vdda, vss;

input  en, enb, inn, inp;

input [3:0]  gear;
input [3:0]  gearb;


wphy_pi_4g_PU_D1_GL16_RVT PUDUM1 ( .vdd(vdda), .en(vdda), .y(outp));

wphy_pi_4g_PU_D1_GL16_RVT PU0 ( .vdd(vdda), .en(en), .y(outn));

wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p5 INV7 ( .en(gear[0]), .enb(gearb[0]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p5 INV0 ( .en(gear[0]), .enb(gearb[0]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p25 I3 ( .en(en), .enb(enb), .in(inp), .vss(vss), 
    .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p25 I2 ( .en(en), .enb(enb), .in(inn), .vss(vss), 
    .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV6_1 ( .en(gear[2]), .enb(gearb[2]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV6_0 ( .en(gear[2]), .enb(gearb[2]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve I1 ( .en(gear[1]), .enb(gearb[1]), .in(inn), .vss(vss), 
    .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve I0 ( .en(gear[1]), .enb(gearb[1]), .in(inp), .vss(vss), 
    .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV1_1 ( .en(gear[2]), .enb(gearb[2]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV1_0 ( .en(gear[2]), .enb(gearb[2]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV2_3 ( .en(gear[3]), .enb(gearb[3]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV2_2 ( .en(gear[3]), .enb(gearb[3]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV2_1 ( .en(gear[3]), .enb(gearb[3]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV2_0 ( .en(gear[3]), .enb(gearb[3]), .in(inn), 
    .vss(vss), .out(outp), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV4_3 ( .en(gear[3]), .enb(gearb[3]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV4_2 ( .en(gear[3]), .enb(gearb[3]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV4_1 ( .en(gear[3]), .enb(gearb[3]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_wphy_pi_4g_inve INV4_0 ( .en(gear[3]), .enb(gearb[3]), .in(inp), 
    .vss(vss), .out(outn), .vdda(vdda));

wphy_pi_4g_PD_D1_GL16_RVT PDDUM1 ( .vss(vss), .enb(vss), .y(outn));

wphy_pi_4g_PD_D1_GL16_RVT PD0 ( .vss(vss), .enb(enb), .y(outp));

endmodule
// Library - wphy_gf12lp_ips_lib, Cell - wphy_pi_4g, View - schematic
// LAST TIME SAVED: Oct 23 12:01:12 2020
// NETLIST TIME: Oct 28 22:02:33 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_pi_4g (out, outb,   clk0, clk90, clk180, clk270, 
    code, ena, gear, quad, xcpl
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  out, outb;



input  clk0, clk90, clk180, clk270, ena;

input [15:0]  code;
input [3:0]  gear;
input [3:0]  xcpl;
input [1:0]  quad;

// Buses in the design 
`ifdef SYNTHESIS 
`else

wire  [15:0]  sel90;

wire  [15:0]  sel0;

wire  [15:0]  sel90b;

wire  [15:0]  sel0b;

wire  [3:0]  gear_intb;

wire  [15:0]  sel270;

wire  [15:0]  sel180b;

wire  [15:0]  sel270b;

wire  [3:0]  gear_int;

wire  [3:0]  xcpl_int;

wire  [15:0]  sel180;

wire  [3:0]  xcplb_int;


wphy_pi_4g_TIELO_D2_GL16_RVT TIELO0 ( .tielo(tielo), .vss(vss), .vdd(vdda));

wphy_pi_4g_TIEHI_D2_GL16_RVT TIEHI0 ( .tiehi(tiehi), .vss(vss), .vdd(vdda));

wphy_pi_4g_wphy_pi_4g_outdrv Ioutdrv ( .vss(vss), .tielo(tielo), .outp(out), 
    .outn(outb), .inp(mix_outp), .inn(mix_outn), .vdda(vdda), 
    .tiehi(tiehi));

wphy_pi_4g_wphy_pi_4g_core core ( .vdda(vdda), .vss(vss), .outn(mix_outn), 
    .outp(mix_outp), .clk0(preclk0), .clk90(preclk90), 
    .clk180(preclk180), .clk270(preclk270), .sel0(sel0), .sel0b(sel0b), 
    .sel90(sel90), .sel90b(sel90b), .sel180(sel180), .sel180b(sel180b), 
    .sel270(sel270), .sel270b(sel270b), .xcpl(xcpl_int), 
    .xcplb(xcplb_int));

wphy_pi_4g_wphy_pi_logic Ipi_logic ( .gear_out(gear_int[3:0]), 
    .gear_outb(gear_intb[3:0]), .enb_int(enb_int), .en_int(en_int), 
    .en(ena), .xcpl_in(xcpl[3:0]), .gear(gear[3:0]), .vss(vss), 
    .tielo(tielo), .xcplb(xcplb_int[3:0]), .xcpl(xcpl_int[3:0]), 
    .sel270b(sel270b[15:0]), .sel270(sel270[15:0]), 
    .sel180b(sel180b[15:0]), .sel180(sel180[15:0]), 
    .sel90b(sel90b[15:0]), .sel90(sel90[15:0]), .sel0b(sel0b[15:0]), 
    .sel0(sel0[15:0]), .tiehi(tiehi), .vdda(vdda), .quad(quad[1:0]), 
    .code(code[15:0]));

wphy_pi_4g_wphy_pi_4g_predrv predrvQ ( .vdda(vdda), .en(en_int), .enb(enb_int), 
    .gearb(gear_intb[3:0]), .vss(vss), .inp(clk90), .inn(clk270), 
    .outp(preclk90), .outn(preclk270), .gear(gear_int[3:0]));

wphy_pi_4g_wphy_pi_4g_predrv predrvI ( .vdda(vdda), .en(en_int), .enb(enb_int), 
    .gearb(gear_intb[3:0]), .vss(vss), .inp(clk0), .inn(clk180), 
    .outp(preclk0), .outn(preclk180), .gear(gear_int[3:0]));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// HDL file - wphy_gf12lp_ips_sim_lib, wphy_pi_4g_stim, systemVerilog.

// Library - wphy_gf12lp_ips_sim_lib, Cell - wphy_pi_4g_tb, View -
//schematic
// LAST TIME SAVED: Oct 28 21:48:07 2020
// NETLIST TIME: Oct 28 22:02:33 2020

module wphy_pi_4g_PD_D1_GL16_RVT( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//Verilog HDL for "wmx_d2d_serdes_lib", "wmx_d2d_pi_cmos_inv1_en" "functional"


module wphy_pi_4g_wphy_pi_4g_inve ( in, vdda, vss, out, en, enb );

  input in;
  inout vdda;
  output out;
  input en;
  input enb;
  inout vss;
  wire pwr_ok;

  assign pwr_ok = vdda & ~vss;
  assign out= pwr_ok ? ( en ? ~in:1'bz) : 1'bx ;

endmodule
//Verilog HDL for "wphy_ln08lpu_ips_lib", "wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p25" "functional"


module wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p25 ( in, vdda, vss, out, en, enb );

  input in;
  inout vdda;
  output out;
  input en;
  input enb;
  inout vss;

  wire polarity_ok = en ^ enb;
  wire pwr_ok;

  assign pwr_ok = vdda & ~vss;
  assign out= (pwr_ok&polarity_ok) ? ( en ? ~in:1'bz) : 1'bx ;


endmodule
//Verilog HDL for "wmx_d2d_serdes_lib", "wmx_d2d_pi_cmos_inv1_en" "functional"


module wphy_pi_4g_wphy_pi_4g_wphy_pi_4g_inve_0p5 ( in, vdda, vss, out, en, enb );

  input in;
  inout vdda;
  output out;
  input en;
  input enb;
  inout vss;
  wire pwr_ok;

  assign pwr_ok = vdda & ~vss;
  assign out= pwr_ok ? ( en ? ~in:1'bz) : 1'bx ;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_pi_4g_PU_D1_GL16_RVT" "systemVerilog"


module wphy_pi_4g_PU_D1_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule



module wphy_pi_4g_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_pi_4g_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_pi_4g_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//systemVerilog HDL for "wphy_ln08lpu_ips_lib", "wphy_pi_4g_wphy_pi_4g_core" "systemVerilog"

`timescale 1ps/1fs
module wphy_pi_4g_wphy_pi_4g_core ( outn, outp, vdda, vss, clk0, clk90, clk180, clk270,
sel0, sel0b, sel90, sel90b, sel180, sel180b, sel270, sel270b, xcpl, xcplb );

  input  [3:0] xcplb;
  input  [3:0] xcpl;
  input  [15:0] sel270;
  input  [15:0] sel270b;
  input clk270;
  input  [15:0] sel90b;
  input clk90;
  input  [15:0] sel90;

  input  [15:0] sel180;
  input  [15:0] sel180b;
  input clk180;
  input clk0;

  input  [15:0] sel0b;
  input  [15:0] sel0;

  inout vdda;
  inout vss;
  output reg outp = 1'b0;
  output wire outn;

//reg outp = 1'b0;

reg outp_int = 1'b0;
//reg       outp_int;


wire [63:0]       therm_code;
real        current_edge0, previous_edge0, current_period0;
real        current_edge90, previous_edge90, current_period90;
real        current_edge180, previous_edge180, current_period180;
real        current_edge270, previous_edge270, current_period270;
real        phase_step0, phase_step90, phase_step180, phase_step270;
real        phase_delay0, phase_delay90, phase_delay180, phase_delay270;
integer        delay_count, delay_count_mod;
reg         out_int;
wire [15:0]    tsel0, tsel90, tsel180, tsel270;
wire        power_ok;
reg         del_270_0, del_0_90, del_90_180, del_180_270;

reg         genclk0, genclk90, genclk180, genclk270;

assign power_ok = (vdda & ~vss);

assign tsel0      =  sel0     & ~sel0b;
assign tsel90     =  sel90    & ~sel90b;
assign tsel180 =  sel180   & ~sel180b;
assign tsel270 =  sel270   & ~sel270b;


assign therm_code = {tsel0, tsel90, tsel180, tsel270};

integer ones0;
integer ones90;
integer ones180;
integer ones270;
integer ones [3:0];
real tmin_delay=0.0;
reg assert_en=1'b0;
integer clk0_edges=0;

initial begin
  ones0=$countones(tsel0);
  ones90=$countones(tsel90);
  ones180=$countones(tsel180);
  ones270=$countones(tsel270);

  ones[0]=ones0;
  ones[1]=ones90;
  ones[2]=ones180;
  ones[3]=ones270;
end

initial begin
   if ($value$plusargs("WPHY_ANA_ASSERT_EN=%f", assert_en)) begin
      assert_en=assert_en;
   end
end


always @(tsel0) begin
  ones0=$countones(tsel0);
end
always @(tsel90) begin
  ones90=$countones(tsel90);
end
always @(tsel180) begin
  ones180=$countones(tsel180);
end
always @(tsel270) begin
  ones270=$countones(tsel270);
end

always @(*) begin
  ones[0]=ones0;
  ones[1]=ones90;
  ones[2]=ones180;
  ones[3]=ones270;
end


// BIG TABLE, will change if I have some time
always @(*) begin

   //therm_code_ones = $countones
   case({ones[0],ones[1],ones[2],ones[3]})
    {32'd00,32'd0,32'd0,32'd16}:delay_count = 0;
    {32'd01,32'd0,32'd0,32'd15}:delay_count = 1;
    {32'd02,32'd0,32'd0,32'd14}:delay_count = 2;
    {32'd03,32'd0,32'd0,32'd13}:delay_count = 3;
    {32'd04,32'd0,32'd0,32'd12}:delay_count = 4;
    {32'd05,32'd0,32'd0,32'd11}:delay_count = 5;
    {32'd06,32'd0,32'd0,32'd10}:delay_count = 6;
    {32'd07,32'd0,32'd0,32'd09}:delay_count = 7;
    {32'd08,32'd0,32'd0,32'd08}:delay_count = 8;
    {32'd09,32'd0,32'd0,32'd07}:delay_count = 9;
    {32'd10,32'd0,32'd0,32'd06}:delay_count = 10;
    {32'd11,32'd0,32'd0,32'd05}:delay_count = 11;
    {32'd12,32'd0,32'd0,32'd04}:delay_count = 12;
    {32'd13,32'd0,32'd0,32'd03}:delay_count = 13;
    {32'd14,32'd0,32'd0,32'd02}:delay_count = 14;
    {32'd15,32'd0,32'd0,32'd01}:delay_count = 15;

    {32'd16,32'd00,32'd0,32'd0}:delay_count = 16;
    {32'd15,32'd01,32'd0,32'd0}:delay_count = 17;
    {32'd14,32'd02,32'd0,32'd0}:delay_count = 18;
    {32'd13,32'd03,32'd0,32'd0}:delay_count = 19;
    {32'd12,32'd04,32'd0,32'd0}:delay_count = 20;
    {32'd11,32'd05,32'd0,32'd0}:delay_count = 21;
    {32'd10,32'd06,32'd0,32'd0}:delay_count = 22;
    {32'd09,32'd07,32'd0,32'd0}:delay_count = 23;
    {32'd08,32'd08,32'd0,32'd0}:delay_count = 24;
    {32'd07,32'd09,32'd0,32'd0}:delay_count = 25;
    {32'd06,32'd10,32'd0,32'd0}:delay_count = 26;
    {32'd05,32'd11,32'd0,32'd0}:delay_count = 27;
    {32'd04,32'd12,32'd0,32'd0}:delay_count = 28;
    {32'd03,32'd13,32'd0,32'd0}:delay_count = 29;
    {32'd02,32'd14,32'd0,32'd0}:delay_count = 30;
    {32'd01,32'd15,32'd0,32'd0}:delay_count = 31;

    {32'd00,32'd16,32'd00,32'd0}:delay_count = 32;
    {32'd00,32'd15,32'd01,32'd0}:delay_count = 33;
    {32'd00,32'd14,32'd02,32'd0}:delay_count = 34;
    {32'd00,32'd13,32'd03,32'd0}:delay_count = 35;
    {32'd00,32'd12,32'd04,32'd0}:delay_count = 36;
    {32'd00,32'd11,32'd05,32'd0}:delay_count = 37;
    {32'd00,32'd10,32'd06,32'd0}:delay_count = 38;
    {32'd00,32'd09,32'd07,32'd0}:delay_count = 39;
    {32'd00,32'd08,32'd08,32'd0}:delay_count = 40;
    {32'd00,32'd07,32'd09,32'd0}:delay_count = 41;
    {32'd00,32'd06,32'd10,32'd0}:delay_count = 42;
    {32'd00,32'd05,32'd11,32'd0}:delay_count = 43;
    {32'd00,32'd04,32'd12,32'd0}:delay_count = 44;
    {32'd00,32'd03,32'd13,32'd0}:delay_count = 45;
    {32'd00,32'd02,32'd14,32'd0}:delay_count = 46;
    {32'd00,32'd01,32'd15,32'd0}:delay_count = 47;

    {32'd00,32'd00,32'd16,32'd00}:delay_count = 48;
    {32'd00,32'd00,32'd15,32'd01}:delay_count = 49;
    {32'd00,32'd00,32'd14,32'd02}:delay_count = 50;
    {32'd00,32'd00,32'd13,32'd03}:delay_count = 51;
    {32'd00,32'd00,32'd12,32'd04}:delay_count = 52;
    {32'd00,32'd00,32'd11,32'd05}:delay_count = 53;
    {32'd00,32'd00,32'd10,32'd06}:delay_count = 54;
    {32'd00,32'd00,32'd09,32'd07}:delay_count = 55;
    {32'd00,32'd00,32'd08,32'd08}:delay_count = 56;
    {32'd00,32'd00,32'd07,32'd09}:delay_count = 57;
    {32'd00,32'd00,32'd06,32'd10}:delay_count = 58;
    {32'd00,32'd00,32'd05,32'd11}:delay_count = 59;
    {32'd00,32'd00,32'd04,32'd12}:delay_count = 60;
    {32'd00,32'd00,32'd03,32'd13}:delay_count = 61;
    {32'd00,32'd00,32'd02,32'd14}:delay_count = 62;
    {32'd00,32'd00,32'd01,32'd15}:delay_count = 63;

    default : delay_count = delay_count;
   endcase
  delay_count_mod = delay_count % 16;
end


                  


//period
always @(posedge clk0) begin 
  current_edge0            = $realtime;
  current_period0          = current_edge0 - previous_edge0;
  if(current_period0 > 5000) begin
    current_period0     = 5000;
  end
  previous_edge0           = current_edge0;
  phase_step0              = current_period0 / 64;
  //phase_delay0             = del_270_0 ? ((delay_count_mod+1) * phase_step0) : (del_0_90 ? ((15 - delay_count_mod) * phase_step0) : 0);
  phase_delay0             = del_0_90 ? ((delay_count_mod) * phase_step0) : 0;


  
  if(Ipi_logic.en & assert_en) begin
    if(clk0_edges<5)
     clk0_edges = clk0_edges+1;
    else
      if(current_period0 > 5000)
        $display("WPHY_ANA_ERROR: input PI frequency too low (needs to be >500MHz),  %m at %t",$realtime);

  end
  else
    clk0_edges=0;

end

always @(posedge clk90) begin 
  current_edge90           = $realtime;
  current_period90         = current_edge90 - previous_edge90;
  if(current_period90 > 5000) begin
    current_period90     = 5000;
  end
  previous_edge90          = current_edge90;
  phase_step90                = current_period90 / 64;
  //phase_delay90            = del_0_90 ? ((delay_count_mod+1) * phase_step90) : (del_90_180 ? ((15 - delay_count_mod) * phase_step90) : 0);
  phase_delay90            = del_90_180 ? ((delay_count_mod) * phase_step90) : 0;
end

always @(posedge clk180) begin 
  current_edge180             = $realtime;
  current_period180        = current_edge180 - previous_edge180;
  if(current_period180 > 5000) begin
    current_period180     = 5000;
  end
  previous_edge180            = current_edge180;
  phase_step180               = current_period180 / 64;
  //phase_delay180              = del_90_180 ? ((delay_count_mod+1) * phase_step180) : (del_180_270 ? ((15 - delay_count_mod) * phase_step180) : 0);
  phase_delay180              = del_180_270 ? ((delay_count_mod) * phase_step180) : 0;
end

always @(posedge clk270) begin 
  current_edge270             = $realtime;
  current_period270        = current_edge270 - previous_edge270;
  if(current_period270 > 5000) begin
    current_period270     = 5000;
  end
  previous_edge270            = current_edge270;
  phase_step270               = (current_period270 / 64) + 0.001;
  //phase_delay270              = del_180_270 ? ((delay_count_mod+1) * phase_step270) : (del_270_0 ? ((15 - delay_count_mod) * phase_step270) : 0);
  phase_delay270              = del_270_0 ? ((delay_count_mod) * phase_step270) : 0;
end



always @(clk0) begin
   if(clk0) genclk0 = #(phase_delay0) 1'b1;
  else         genclk0 = #(phase_delay0) 1'b0;
end        
          
always @(clk90) begin
 if(clk90) genclk90 = #(phase_delay90) 1'b1;
 else      genclk90 = #(phase_delay90) 1'b0;
end  

always @(clk180) begin
   if(clk180) genclk180 = #(phase_delay180) 1'b1;
 else        genclk180 = #(phase_delay180) 1'b0;
end  

always @(clk270) begin
   if(clk270) genclk270 = #(phase_delay270) 1'b1;
 else        genclk270 = #(phase_delay270) 1'b0;
end  


//always @(*) begin
always@(genclk0 or genclk90 or genclk180 or genclk270) begin
    #0;
   //case({del_270_0, del_0_90, del_90_180, del_180_270})
   case({del_0_90, del_90_180, del_180_270,del_270_0})
    4'b1000 : outp_int = genclk0;
    4'b0100 : outp_int = genclk90;
    4'b0010 : outp_int = genclk180;
    4'b0001 : outp_int = genclk270;
    default : outp_int = outp;
  endcase
end

initial begin
   case(Ipi_logic.gear)
      0: tmin_delay = 454.0;
      1: tmin_delay = 335.0;
      2: tmin_delay = 250.0;
      3: tmin_delay = 245.0;
      4: tmin_delay = 160.0;
      5: tmin_delay = 157.0;
      6: tmin_delay = 154.0;
      7: tmin_delay = 153.0;
      8: tmin_delay = 140.0;
      9: tmin_delay = 134.0;
      10: tmin_delay = 126.0;
      11: tmin_delay = 125.0;
      12: tmin_delay = 109.0;
      13: tmin_delay = 108.0;
      14: tmin_delay = 107.0;
      15: tmin_delay = 106.0;
      default: tmin_delay = 50.0;
   endcase
end
always @(Ipi_logic.gear) begin
   case(Ipi_logic.gear)
      0: tmin_delay = 454.0;
      1: tmin_delay = 335.0;
      2: tmin_delay = 250.0;
      3: tmin_delay = 245.0;
      4: tmin_delay = 160.0;
      5: tmin_delay = 157.0;
      6: tmin_delay = 154.0;
      7: tmin_delay = 153.0;
      8: tmin_delay = 140.0;
      9: tmin_delay = 134.0;
      10: tmin_delay = 126.0;
      11: tmin_delay = 125.0;
      12: tmin_delay = 109.0;
      13: tmin_delay = 108.0;
      14: tmin_delay = 107.0;
      15: tmin_delay = 106.0;
      default: tmin_delay = 50.0;
   endcase
end

always @(outp_int) begin
  outp <= #(tmin_delay) outp_int;
end

always @(delay_count) begin
  del_270_0    = (delay_count>=0)   && (delay_count<=15);
  del_0_90     = (delay_count>=16)  && (delay_count<=31);
  del_90_180   = (delay_count>=32)  && (delay_count<=47);
  del_180_270  = (delay_count>=48)  && (delay_count<=63);
end


assign outn = ~outp;              

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_pi_4g_INV_D1_GL16_RVT_Mmod_nomodel"
//"systemVerilog"


module wphy_pi_4g_INV_D1_GL16_RVT_Mmod_nomodel ( in, out, tiehi, tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
  input tiehi;
  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_pi_4g_INV_D2_GL16_RVT" "systemVerilog"


module wphy_pi_4g_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_pi_4g_TIEHI_D2_GL16_RVT" "systemVerilog"


module wphy_pi_4g_TIEHI_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);


  output tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tiehi = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tiehi =  1'b1 ;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_pi_4g_TIELO_D2_GL16_RVT" "systemVerilog"


module wphy_pi_4g_TIELO_D2_GL16_RVT ( tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd
`endif //WLOGIC_MODEL_NO_PG
);

  output tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;

  assign tielo = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign tielo =  1'b0 ;


endmodule
`endif //SYNTHESIS
