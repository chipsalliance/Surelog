// CRC32 based on https://msdn.microsoft.com/en-us/library/dd905031.aspx
//
// 
//
//
//

module crc32 (input [7:0] din, input clk, input rst_n, output [31:0] dout);

  reg [31:0] crctbl [255:0];
  reg [31:0] crc;

  initial
    begin
        crctbl[0] <= 32'h00000000;
        crctbl[1] <= 32'h77073096;
        crctbl[2] <= 32'hEE0E612C;
        crctbl[3] <= 32'h990951BA;
        crctbl[4] <= 32'h076DC419;
        crctbl[5] <= 32'h706AF48F;
        crctbl[6] <= 32'hE963A535;
        crctbl[7] <= 32'h9E6495A3;
        crctbl[8] <= 32'h0EDB8832;
        crctbl[9] <= 32'h79DCB8A4;
        crctbl[10] <= 32'hE0D5E91E;
        crctbl[11] <= 32'h97D2D988;
        crctbl[12] <= 32'h09B64C2B;
        crctbl[13] <= 32'h7EB17CBD;
        crctbl[14] <= 32'hE7B82D07;
        crctbl[15] <= 32'h90BF1D91;
        crctbl[16] <= 32'h1DB71064;
        crctbl[17] <= 32'h6AB020F2;
        crctbl[18] <= 32'hF3B97148;
        crctbl[19] <= 32'h84BE41DE;
        crctbl[20] <= 32'h1ADAD47D;
        crctbl[21] <= 32'h6DDDE4EB;
        crctbl[22] <= 32'hF4D4B551;
        crctbl[23] <= 32'h83D385C7;
        crctbl[24] <= 32'h136C9856;
        crctbl[25] <= 32'h646BA8C0;
        crctbl[26] <= 32'hFD62F97A;
        crctbl[27] <= 32'h8A65C9EC;
        crctbl[28] <= 32'h14015C4F;
        crctbl[29] <= 32'h63066CD9;
        crctbl[30] <= 32'hFA0F3D63;
        crctbl[31] <= 32'h8D080DF5;
        crctbl[32] <= 32'h3B6E20C8;
        crctbl[33] <= 32'h4C69105E;
        crctbl[34] <= 32'hD56041E4;
        crctbl[35] <= 32'hA2677172;
        crctbl[36] <= 32'h3C03E4D1;
        crctbl[37] <= 32'h4B04D447;
        crctbl[38] <= 32'hD20D85FD;
        crctbl[39] <= 32'hA50AB56B;
        crctbl[40] <= 32'h35B5A8FA;
        crctbl[41] <= 32'h42B2986C;
        crctbl[42] <= 32'hDBBBC9D6;
        crctbl[43] <= 32'hACBCF940;
        crctbl[44] <= 32'h32D86CE3;
        crctbl[45] <= 32'h45DF5C75;
        crctbl[46] <= 32'hDCD60DCF;
        crctbl[47] <= 32'hABD13D59;
        crctbl[48] <= 32'h26D930AC;
        crctbl[49] <= 32'h51DE003A;
        crctbl[50] <= 32'hC8D75180;
        crctbl[51] <= 32'hBFD06116;
        crctbl[52] <= 32'h21B4F4B5;
        crctbl[53] <= 32'h56B3C423;
        crctbl[54] <= 32'hCFBA9599;
        crctbl[55] <= 32'hB8BDA50F;
        crctbl[56] <= 32'h2802B89E;
        crctbl[57] <= 32'h5F058808;
        crctbl[58] <= 32'hC60CD9B2;
        crctbl[59] <= 32'hB10BE924;
        crctbl[60] <= 32'h2F6F7C87;
        crctbl[61] <= 32'h58684C11;
        crctbl[62] <= 32'hC1611DAB;
        crctbl[63] <= 32'hB6662D3D;
        crctbl[64] <= 32'h76DC4190;
        crctbl[65] <= 32'h01DB7106;
        crctbl[66] <= 32'h98D220BC;
        crctbl[67] <= 32'hEFD5102A;
        crctbl[68] <= 32'h71B18589;
        crctbl[69] <= 32'h06B6B51F;
        crctbl[70] <= 32'h9FBFE4A5;
        crctbl[71] <= 32'hE8B8D433;
        crctbl[72] <= 32'h7807C9A2;
        crctbl[73] <= 32'h0F00F934;
        crctbl[74] <= 32'h9609A88E;
        crctbl[75] <= 32'hE10E9818;
        crctbl[76] <= 32'h7F6A0DBB;
        crctbl[77] <= 32'h086D3D2D;
        crctbl[78] <= 32'h91646C97;
        crctbl[79] <= 32'hE6635C01;
        crctbl[80] <= 32'h6B6B51F4;
        crctbl[81] <= 32'h1C6C6162;
        crctbl[82] <= 32'h856530D8;
        crctbl[83] <= 32'hF262004E;
        crctbl[84] <= 32'h6C0695ED;
        crctbl[85] <= 32'h1B01A57B;
        crctbl[86] <= 32'h8208F4C1;
        crctbl[87] <= 32'hF50FC457;
        crctbl[88] <= 32'h65B0D9C6;
        crctbl[89] <= 32'h12B7E950;
        crctbl[90] <= 32'h8BBEB8EA;
        crctbl[91] <= 32'hFCB9887C;
        crctbl[92] <= 32'h62DD1DDF;
        crctbl[93] <= 32'h15DA2D49;
        crctbl[94] <= 32'h8CD37CF3;
        crctbl[95] <= 32'hFBD44C65;
        crctbl[96] <= 32'h4DB26158;
        crctbl[97] <= 32'h3AB551CE;
        crctbl[98] <= 32'hA3BC0074;
        crctbl[99] <= 32'hD4BB30E2;
        crctbl[100] <= 32'h4ADFA541;
        crctbl[101] <= 32'h3DD895D7;
        crctbl[102] <= 32'hA4D1C46D;
        crctbl[103] <= 32'hD3D6F4FB;
        crctbl[104] <= 32'h4369E96A;
        crctbl[105] <= 32'h346ED9FC;
        crctbl[106] <= 32'hAD678846;
        crctbl[107] <= 32'hDA60B8D0;
        crctbl[108] <= 32'h44042D73;
        crctbl[109] <= 32'h33031DE5;
        crctbl[110] <= 32'hAA0A4C5F;
        crctbl[111] <= 32'hDD0D7CC9;
        crctbl[112] <= 32'h5005713C;
        crctbl[113] <= 32'h270241AA;
        crctbl[114] <= 32'hBE0B1010;
        crctbl[115] <= 32'hC90C2086;
        crctbl[116] <= 32'h5768B525;
        crctbl[117] <= 32'h206F85B3;
        crctbl[118] <= 32'hB966D409;
        crctbl[119] <= 32'hCE61E49F;
        crctbl[120] <= 32'h5EDEF90E;
        crctbl[121] <= 32'h29D9C998;
        crctbl[122] <= 32'hB0D09822;
        crctbl[123] <= 32'hC7D7A8B4;
        crctbl[124] <= 32'h59B33D17;
        crctbl[125] <= 32'h2EB40D81;
        crctbl[126] <= 32'hB7BD5C3B;
        crctbl[127] <= 32'hC0BA6CAD;
        crctbl[128] <= 32'hEDB88320;
        crctbl[129] <= 32'h9ABFB3B6;
        crctbl[130] <= 32'h03B6E20C;
        crctbl[131] <= 32'h74B1D29A;
        crctbl[132] <= 32'hEAD54739;
        crctbl[133] <= 32'h9DD277AF;
        crctbl[134] <= 32'h04DB2615;
        crctbl[135] <= 32'h73DC1683;
        crctbl[136] <= 32'hE3630B12;
        crctbl[137] <= 32'h94643B84;
        crctbl[138] <= 32'h0D6D6A3E;
        crctbl[139] <= 32'h7A6A5AA8;
        crctbl[140] <= 32'hE40ECF0B;
        crctbl[141] <= 32'h9309FF9D;
        crctbl[142] <= 32'h0A00AE27;
        crctbl[143] <= 32'h7D079EB1;
        crctbl[144] <= 32'hF00F9344;
        crctbl[145] <= 32'h8708A3D2;
        crctbl[146] <= 32'h1E01F268;
        crctbl[147] <= 32'h6906C2FE;
        crctbl[148] <= 32'hF762575D;
        crctbl[149] <= 32'h806567CB;
        crctbl[150] <= 32'h196C3671;
        crctbl[151] <= 32'h6E6B06E7;
        crctbl[152] <= 32'hFED41B76;
        crctbl[153] <= 32'h89D32BE0;
        crctbl[154] <= 32'h10DA7A5A;
        crctbl[155] <= 32'h67DD4ACC;
        crctbl[156] <= 32'hF9B9DF6F;
        crctbl[157] <= 32'h8EBEEFF9;
        crctbl[158] <= 32'h17B7BE43;
        crctbl[159] <= 32'h60B08ED5;
        crctbl[160] <= 32'hD6D6A3E8;
        crctbl[161] <= 32'hA1D1937E;
        crctbl[162] <= 32'h38D8C2C4;
        crctbl[163] <= 32'h4FDFF252;
        crctbl[164] <= 32'hD1BB67F1;
        crctbl[165] <= 32'hA6BC5767;
        crctbl[166] <= 32'h3FB506DD;
        crctbl[167] <= 32'h48B2364B;
        crctbl[168] <= 32'hD80D2BDA;
        crctbl[169] <= 32'hAF0A1B4C;
        crctbl[170] <= 32'h36034AF6;
        crctbl[171] <= 32'h41047A60;
        crctbl[172] <= 32'hDF60EFC3;
        crctbl[173] <= 32'hA867DF55;
        crctbl[174] <= 32'h316E8EEF;
        crctbl[175] <= 32'h4669BE79;
        crctbl[176] <= 32'hCB61B38C;
        crctbl[177] <= 32'hBC66831A;
        crctbl[178] <= 32'h256FD2A0;
        crctbl[179] <= 32'h5268E236;
        crctbl[180] <= 32'hCC0C7795;
        crctbl[181] <= 32'hBB0B4703;
        crctbl[182] <= 32'h220216B9;
        crctbl[183] <= 32'h5505262F;
        crctbl[184] <= 32'hC5BA3BBE;
        crctbl[185] <= 32'hB2BD0B28;
        crctbl[186] <= 32'h2BB45A92;
        crctbl[187] <= 32'h5CB36A04;
        crctbl[188] <= 32'hC2D7FFA7;
        crctbl[189] <= 32'hB5D0CF31;
        crctbl[190] <= 32'h2CD99E8B;
        crctbl[191] <= 32'h5BDEAE1D;
        crctbl[192] <= 32'h9B64C2B0;
        crctbl[193] <= 32'hEC63F226;
        crctbl[194] <= 32'h756AA39C;
        crctbl[195] <= 32'h026D930A;
        crctbl[196] <= 32'h9C0906A9;
        crctbl[197] <= 32'hEB0E363F;
        crctbl[198] <= 32'h72076785;
        crctbl[199] <= 32'h05005713;
        crctbl[200] <= 32'h95BF4A82;
        crctbl[201] <= 32'hE2B87A14;
        crctbl[202] <= 32'h7BB12BAE;
        crctbl[203] <= 32'h0CB61B38;
        crctbl[204] <= 32'h92D28E9B;
        crctbl[205] <= 32'hE5D5BE0D;
        crctbl[206] <= 32'h7CDCEFB7;
        crctbl[207] <= 32'h0BDBDF21;
        crctbl[208] <= 32'h86D3D2D4;
        crctbl[209] <= 32'hF1D4E242;
        crctbl[210] <= 32'h68DDB3F8;
        crctbl[211] <= 32'h1FDA836E;
        crctbl[212] <= 32'h81BE16CD;
        crctbl[213] <= 32'hF6B9265B;
        crctbl[214] <= 32'h6FB077E1;
        crctbl[215] <= 32'h18B74777;
        crctbl[216] <= 32'h88085AE6;
        crctbl[217] <= 32'hFF0F6A70;
        crctbl[218] <= 32'h66063BCA;
        crctbl[219] <= 32'h11010B5C;
        crctbl[220] <= 32'h8F659EFF;
        crctbl[221] <= 32'hF862AE69;
        crctbl[222] <= 32'h616BFFD3;
        crctbl[223] <= 32'h166CCF45;
        crctbl[224] <= 32'hA00AE278;
        crctbl[225] <= 32'hD70DD2EE;
        crctbl[226] <= 32'h4E048354;
        crctbl[227] <= 32'h3903B3C2;
        crctbl[228] <= 32'hA7672661;
        crctbl[229] <= 32'hD06016F7;
        crctbl[230] <= 32'h4969474D;
        crctbl[231] <= 32'h3E6E77DB;
        crctbl[232] <= 32'hAED16A4A;
        crctbl[233] <= 32'hD9D65ADC;
        crctbl[234] <= 32'h40DF0B66;
        crctbl[235] <= 32'h37D83BF0;
        crctbl[236] <= 32'hA9BCAE53;
        crctbl[237] <= 32'hDEBB9EC5;
        crctbl[238] <= 32'h47B2CF7F;
        crctbl[239] <= 32'h30B5FFE9;
        crctbl[240] <= 32'hBDBDF21C;
        crctbl[241] <= 32'hCABAC28A;
        crctbl[242] <= 32'h53B39330;
        crctbl[243] <= 32'h24B4A3A6;
        crctbl[244] <= 32'hBAD03605;
        crctbl[245] <= 32'hCDD70693;
        crctbl[246] <= 32'h54DE5729;
        crctbl[247] <= 32'h23D967BF;
        crctbl[248] <= 32'hB3667A2E;
        crctbl[249] <= 32'hC4614AB8;
        crctbl[250] <= 32'h5D681B02;
        crctbl[251] <= 32'h2A6F2B94;
        crctbl[252] <= 32'hB40BBE37;
        crctbl[253] <= 32'hC30C8EA1;
        crctbl[254] <= 32'h5A05DF1B;
        crctbl[255] <= 32'h2D02EF8D;
    end

  always @(posedge clk)
  begin
    if (rst_n == 1'b0)
      crc <= 32'hFFFFFFFF;
    else
      crc <= (crc >> 8) ^ crctbl[(crc[7:0] ^ din)];    
  end

  assign dout = crc;

endmodule