/*
:name: class_test_37
:description: Test
:tags: 6.15 8.3
*/
virtual class foo extends bar;
  import fedex_pkg::box;
  import fedex_pkg::*;
endclass