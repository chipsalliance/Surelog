/*
:name: class_member_test_1
:description: Test
:should_fail: 0
:tags: 8.3
*/
class c;
  task intf.task1();
  endtask
endclass