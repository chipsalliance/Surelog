/*
:name: 22.12--line-basic
:description: Test
:should_fail: 0
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 2
