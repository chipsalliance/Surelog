/*
:name: 22.10--celldefine-basic-2
:description: Test
:tags: 22.10
:type: preprocessing
*/
`celldefine
