
`include "inc-1.h"


module a_module(
    input [`BUS_WIDTH] bus
);

endmodule
