/*
:name: class_test_58
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class fields_with_modifiers;
  const static data_type_or_module_type foo1 = 4'hf;
  static const data_type_or_module_type foo3, foo4;
endclass