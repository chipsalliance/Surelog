module test;
    typedef logic [1:0] t_two_bits;
    typedef t_two_bits t_two_bits_copy;
    t_two_bits kkkk;
    t_two_bits_copy zzzz;
endmodule // test
