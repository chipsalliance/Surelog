/*
:name: class_member_test_21
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function sometype #(N+1) subr(ducktype #(3) x);
endclass