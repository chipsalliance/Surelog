module top(output int o);
   localparam unsigned P = 15;
   localparam signed [63:0] n = 32'h8000_0000;
endmodule
