/*
:name: preproc_test_10
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`define LONG_MACRO(\
    a,\
    b, c) text goes here
