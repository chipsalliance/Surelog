module t();
logic [3:0][3:0][7:0] state_d;
assign state_d[2][3][7:0] = 8'b10101010;
endmodule
