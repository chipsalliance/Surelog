module top(output int o);
   function automatic int theta();
      for (int x = 0 ; x < 5 ; x++) begin
         int a, b;
        
         return 0;
      end
      return 0;
   endfunction : theta

endmodule : top
