/*
:name: initial
:description: initial check
:should_fail: 0
:tags: 9.2.1
*/
module initial_tb ();
	reg a = 0;
	initial
		a = 1;
endmodule
