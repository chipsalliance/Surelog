// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: unconnected-drive
:description: Unconnected drive keywords
:tags: 5.6.4
:type: preprocessing
*/


`unconnected_drive pull1

module ts();
endmodule

`nounconnected_drive
