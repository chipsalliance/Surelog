

module mod_3 ();

NO_DEF5 nodef_5();

endmodule
