/*
:name: string_tolower
:description: string.tolower()  tests
:tags: 6.16.5
*/
module top();
	string a = "Test";
	string b = a.tolower();
endmodule
