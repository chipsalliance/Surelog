/*
:name: random_function
:description: $random test
:tags: 20.15
:type: simulation parsing
*/

module top();

initial begin
	$display("%d", $random);
end

endmodule
