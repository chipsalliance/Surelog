module out ();
endmodule
