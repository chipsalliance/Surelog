/*
:name: class_test_36
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class foo;
  import fedex_pkg::box;
  import fedex_pkg::*;
endclass