/*
:name: macromodule_definition
:description: macromodule definition test
:tags: 23.2
*/
macromodule top();

endmodule
