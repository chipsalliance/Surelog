/* wire.h */
reg wire_h;

