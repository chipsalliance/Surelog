/*
:name: resetall-directive
:description: Check for the resetall directive
:tags: 5.6.4
*/

`resetall

module ts();
endmodule
