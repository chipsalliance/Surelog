package pkg;
   typedef struct packed {
      logic 	  x;
   } a;
   typedef a b[5:0];
endpackage // pkg
   
