/*
:name: desc_test_2
:description: Test
:type: preprocessing
:should_fail: 0
:tags: 5.6.4
*/
`ifndef DEBUGGER
`endif
