/*
:name: class_test_3
:description: Test
:tags: 6.15 8.3
*/
class automatic Foo; endclass