/*
:name: union_test_0
:description: Test
:should_fail: 0
:tags: 7.3
*/
typedef union myunion_fwd;