`ifndef BP_COMMON_DEFINES_VH
`define BP_COMMON_DEFINES_VH


`endif

