`define DDR_ANA_CKE_DRVR_LPBK_OVRD_SEL_FIELD      2:0
`define DDR_ANA_CKE_DRVR_LPBK_OVRD_VAL_FIELD      3
`define DDR_ANA_CKE_DRVR_LPBK_RSVD_FIELD          4
`define DDR_ANA_CKE_DRVR_LPBK_SW_OVR_FIELD        5
