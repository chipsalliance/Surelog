// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: comments
:description: A module testing system verilog comments
:tags: 5.4
*/
module empty (
);
  /* multi
     line
     comment
   */

  // single line comment
endmodule
