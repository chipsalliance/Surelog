module top(output string o);
   initial begin
      o = "\\/ _| __| | '_ \\ / _` / ";
   end
endmodule // top
module top(output string o);
   initial begin
      o = "\\/ _| __| | '_ \\ / _` / ";
   end
endmodule // top


