/*
:name: class_test_25
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo implements Package::Bar; endclass