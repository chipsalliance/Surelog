module wtop ();
wsub sub1();
wsub sub2();
wsub sub3();
endmodule

