module top
  (.op({\op[79] ,\op[78] }));

   output \op[79] ;
   output \op[78] ; 
endmodule
