/*
:name: exit_task
:description: $exit test
:should_fail: 0
:tags: 20.2
*/
module top();

initial
	$exit;

endmodule
