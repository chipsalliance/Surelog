/*
:name: class_test_19
:description: Test
:tags: 6.15 8.3
*/
class Foo extends Package::Bar #(x,y,z); endclass