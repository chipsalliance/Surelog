

module Foo ();
 parameter P1 = P2;
 parameter P2 = P1;
 
endmodule

