
module top();

   for (i = 0; i < 3 ; i = i + 1) begin
      assign tmp[i] = 1'b1;
   end

endmodule