/*
:name: class_test_32
:description: Test
:tags: 6.15 8.3
*/
class zzxx;
extern function void set_port(analysis_port #(1) ap);
endclass