module top;
    byte b[] = {1, 1, 1};
    byte o = b.and;
    byte o = b.or;
    byte o = b.xor;
    byte o = b.unique;
endmodule

