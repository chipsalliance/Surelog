module dut();
  unkown_module u0 (a, b, c);
  unkown_module u1 (~a, b, c);
endmodule
