module top(b);integer
inout b;reg c;assign&0=0;assign 0=0;always
i=0;always
if(8)b=_;always
if(8)b=M&0;endmodule
