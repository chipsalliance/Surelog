module top #(
)(
  output bit [6:0]  dmi_req_ram [23:24],
  output bit [6:0]  dmi_req_addr
);
endmodule
