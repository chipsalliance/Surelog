/*
:name: chandle
:description: chandle type tests
:tags: 6.14
*/
module top();
	chandle a;
endmodule
