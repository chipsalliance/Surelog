/*
:name: parameter
:description: parameter tests
:should_fail: 0
:tags: 6.20.2
*/
module top();
	parameter p = 123;
endmodule
