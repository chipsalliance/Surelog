/*
:name: var_local
:description: class with local variable
:tags: 8.18
*/
module class_tb ();
	class a_cls;
		local int a_loc = 2;
	endclass
endmodule
