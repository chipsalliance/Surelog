/*
:name: 22.11--pragma-number
:description: Test
:should_fail: 0
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_number 123
