parameter X = 2;

module top(b,c);
input b;
output c;

parameter Y = 3;

assign c = b;
endmodule

