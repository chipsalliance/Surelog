// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: string_toupper
:description: string.toupper()  tests
:tags: 6.16.4
*/
module top();
	string a = "Test";
	string b = a.toupper();
endmodule
