// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: resetall-directive
:description: Check for the resetall directive
:tags: 5.6.4
*/

`resetall

module ts();
endmodule
