/*
:name: typedef_test_16
:description: Test
:tags: 6.18
*/
typedef struct packed {
  logic [4:0] some_member;
} mystruct_t;