/*
:name: 22.10--celldefine-invalid
:description: Test
:should_fail_because: module must be defined for celldefine to make sense
:tags: 22.10
:type: preprocessing
*/
`celldefine foo
