package pack;

import "DPI-C" context function int uvm_hdl_check_path(string path);

string uvm_aa_string_key;

endpackage

