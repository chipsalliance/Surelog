// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.12--line-complex
:description: Test
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 2
`line 123 "someother" 1
`line 8273 "somefile" 0
`resetall
`line 5 "foo" 2
