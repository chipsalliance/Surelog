/*
:name: 22.7--timescale-basic-1
:description: Test
:tags: 22.7
:type: preprocessing
*/
`timescale 1 ns / 1 ps
