

`define wxyz(I,R = DEFAULT) \
assign abc[I].clk = R.du``I``_clk_x;

