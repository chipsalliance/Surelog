// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.5.2--undef-nonexisting
:description: Test
:tags: 22.5.2
:type: preprocessing
*/
`undef FOO
`undef BAR
