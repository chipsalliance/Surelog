/*
:name: 22.9--unconnected_drive-invalid-2
:description: Test
:should_fail: 1
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull2
`nounconnected_drive
