/*
:name: specparam
:description: specparam tests
:tags: 6.20.5
*/
module top();
	specparam delay = 50;
endmodule
