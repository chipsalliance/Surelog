/*
:name: associative-arrays-wildcard
:description: Test associative arrays support
:tags: 7.8.1 7.8
*/
module top ();

int arr [*];

endmodule
