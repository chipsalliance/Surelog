/*
:name: interface
:description: interface test
:should_fail: 0
:tags: 25.3
*/

interface test_bus;
  logic test_pad;
endinterface: test_bus

module top(test_bus t);

endmodule
