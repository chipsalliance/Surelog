/*
:name: realtime
:description: realtime type tests
:tags: 6.12
*/
module top();
	realtime a = 0.5;
endmodule
