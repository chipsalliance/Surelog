/*
:name: 22.4--include_from_other_directory
:description: Test
:tags: 22.4
:type: preprocessing parsing
*/
`include "include_directory/defs.sv"
module top ();
endmodule
