/*
:name: 22.9--unconnected_drive-basic-2
:description: Test
:should_fail: 0
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull1
