module top(b);
input b;
initial $display("%m");
endmodule

