module test();

reg legal [];

reg [] illegal;

endmodule
