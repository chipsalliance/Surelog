/*
:name: class_member_test_42
:description: Test
:tags: 8.3
*/
class constructible;
function new (string name, virtual time_if vif);
  this.name = name;
endfunction
endclass