/*
:name: real-token
:description: Testing the real variable type
:tags: 5.7.2
*/
module top();
  real a;
endmodule
