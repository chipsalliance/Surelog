module top();
	logic [11:0] first  = 12'h1; 
	logic [11:0] second  = 12'd1; 
	logic [11:0] third  = 12'b1;
	logic [11:0] forth  = 12'o1;
	logic [11:0] fifth  = 1; 
endmodule

