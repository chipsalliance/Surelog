module top ();

   CELL1 cell1();

   CELL2 cell2();

endmodule

