`define DDR_ANA_DQ_DRVR_LPBK_NCAL_FIELD         4:0
`define DDR_ANA_DQ_DRVR_LPBK_PCAL_FIELD         10:5
`define DDR_ANA_DQ_DRVR_LPBK_BS_EN_FIELD        11
`define DDR_ANA_DQ_DRVR_LPBK_LPBK_EN_FIELD      12
