module mytop();
endmodule // mytop
