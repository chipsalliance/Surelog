module top;
   int dynamic1 [];
   int dynamic2 [][1:0];
   int dynamic3 [1:0][];
   int dynamic4 [1:0][][2:0];
   int assoc [int];
   int assoc_string [string];
   int queue [$];
endmodule // top

