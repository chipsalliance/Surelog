/*
:name: class_member_test_24
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subr(mypkg::foo #(4) x[N]);
endclass