module top1 (
input [3:0] S,
input [15:0] D,
output M2,M4,M8,M16
);

endmodule
