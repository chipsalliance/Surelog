/*
:name: typedef_test_0
:description: Test
:tags: 6.18
*/
typedef i_am_a_type_really;