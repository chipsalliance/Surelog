/*
:name: class_member_test_45
:description: Test
:should_fail: 0
:tags: 8.3
*/
class constructible;
extern function new();
endclass