/*
:name: empty_test_1
:description: Test
:type: preprocessing
:tags: 5.3 5.4
*/
    