interface Interface;
    parameter type P;
    P x;
endinterface
module top;
    Interface #(1) intf();
endmodule
