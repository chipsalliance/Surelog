
`unconnected_drive pull0

module test();

endmodule

`nounconnected_drive

`unconnected_drive pull1

`nounconnected_drive
