/*
:name: desc_test_9
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`ifdef FPGA
`ifdef DEBUGGER
module mymod;
endmodule
`endif
`endif
