package pack;

class uvm_port_base;
parameter p1 = 10;
localparam p2 = 5 * p1;
endclass   

endpackage
