/*
:name: class_test_51
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class how_wide;
  localparam Max_int = {$bits(int) - 1{1'b1}};
endclass