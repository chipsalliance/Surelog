`define DDR_ANA_PI_SMALL_CODE_RANGE              4:0
`define DDR_ANA_PI_SMALL_GEAR_RANGE              9:6
`define DDR_ANA_PI_SMALL_EN_RANGE                14

`define DDR_ANA_PI_SMALL_THERM_RANGE             23:16
`define DDR_ANA_PI_SMALL_QUAD_RANGE              33:32

`define DDR_ANA_PI_SMALL_ENC_RANGE               14:0
`define DDR_ANA_PI_SMALL_DEC_RANGE               33:16
