/*
:name: class_test_16
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo #(IFType=virtual x_if);
endclass