module top(b);inout b=0==c;assign c=^K;assign c=9^k;integer c#0;endmodule
