/*
:name: desc_test_7
:description: Test
:type: preprocessing
:should_fail: 0
:tags: 5.6.4
*/
`ifdef DEBUGGER
module mymod;
endmodule
module mymod_different;
endmodule
`endif
