module wsub ();
endmodule

