module adder();
// rtl
m f1();
m f2();
endmodule

module m();
// rtl
endmodule

