module net_vars (input var logic i1 /* var */, input i2 /* net */, input logic i3 /* net */, output var logic o1 /* var */ , output o2 /* net */);

wire a; // net
wire logic b; // net
logic c; // var logic
var d; // var logic
   
endmodule
