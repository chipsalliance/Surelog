/*
:name: class_test_20
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo extends Package::Bar #(.v1(x),.v2(y)); endclass