/*
:name: class_test_26
:description: Test
:tags: 6.15 8.3
*/
class Foo implements Bar#(N); endclass