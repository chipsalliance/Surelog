/*
:name: preproc_test_2
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`include "foo.svh"
`ifndef SANITY
`define SANITY
`endif
