/*
:name: desc_test_4
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
`elsif BORED
`else
`endif
