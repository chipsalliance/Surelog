/*
:name: enum_test_0
:description: Test
:should_fail: 0
:tags: 6.19
*/
typedef enum myenum_fwd;