module top(input clk, output [32:0] o);
assign o = 'bx;
endmodule
