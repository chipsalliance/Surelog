// toto

import wddr_pkg::*;

