/*
:name: 22.5.3--undefineall-basic
:description: Test
:tags: 22.5.3
:type: preprocessing
*/
`undefineall
