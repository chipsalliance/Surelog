/*
:name: 22.9--unconnected_drive-basic-2
:description: Test
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull1
