module OR();
endmodule // OR
