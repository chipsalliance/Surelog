module test;
    typedef logic [1:0] log_two_bits;
    log_two_bits logn;

    typedef reg [1:0] reg_two_bits;
    reg_two_bits regn;

    typedef bit [1:0] bit_two_bits;
    bit_two_bits bitn;

endmodule


