/*
:name: parameter_port_list
:description: parameter port list tests
:tags: 6.20.2
*/
module top #(p = 12);
endmodule
