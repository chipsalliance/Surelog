@0000000  98 00 00 00 78 1c 00 00 3b 9c ff fc b8 00 d8 00
@0000010  78 01 00 00 38 21 80 00 78 02 00 00 38 42 80 08
@0000020  4c 22 00 04 58 20 00 00 34 21 00 04 e3 ff ff fd
@0000030  f8 00 00 46 78 01 de ad 38 02 be ef 58 22 00 00
@0000040  37 9c ff f4 5b 9b 00 08 5b 9d 00 04 34 1b 00 0c
@0000050  b7 7c d8 00 5b 61 00 00 2b 61 00 00 00 21 00 05
@0000060  b8 20 20 00 b8 20 10 00 78 01 00 00 38 21 80 00
@0000070  3c 42 00 02 b4 22 08 00 28 23 00 00 2b 61 00 00
@0000080  20 22 00 1f 34 01 00 01 bc 22 08 00 b8 61 18 00
@0000090  78 01 00 00 38 21 80 00 3c 82 00 02 b4 22 08 00
@00000a0  58 23 00 00 2b 9b 00 08 2b 9d 00 04 37 9c 00 0c
@00000b0  c3 a0 00 00 37 9c ff f4 5b 9b 00 08 5b 9d 00 04
@00000c0  34 1b 00 0c b7 7c d8 00 5b 61 00 00 2b 61 00 00
@00000d0  00 22 00 05 78 01 00 00 38 21 80 00 3c 42 00 02
@00000e0  b4 22 08 00 28 23 00 00 2b 61 00 00 20 22 00 1f
@00000f0  34 01 00 01 bc 22 08 00 a0 61 08 00 7c 21 00 00
@0000100  2b 9b 00 08 2b 9d 00 04 37 9c 00 0c c3 a0 00 00
@0000110  37 9c ff f4 5b 9b 00 08 5b 9d 00 04 34 1b 00 0c
@0000120  b7 7c d8 00 5b 61 00 00 78 01 ff 00 38 21 00 04
@0000130  2b 62 00 00 58 22 00 00 2b 9b 00 08 2b 9d 00 04
@0000140  37 9c 00 0c c3 a0 00 00 37 9c ff ec 5b 9b 00 08
@0000150  5b 9d 00 04 34 1b 00 14 b7 7c d8 00 34 01 00 02
@0000160  fb ff ff ec 34 01 00 00 5b 61 ff f8 e0 00 00 26
@0000170  2b 61 ff f8 fb ff ff d0 b8 20 10 00 34 01 00 00
@0000180  5c 41 00 1e 2b 61 ff f8 b4 21 08 00 34 21 00 03
@0000190  fb ff ff e0 2b 61 ff f8 3c 21 00 02 34 21 00 06
@00001a0  5b 61 ff fc 2b 61 ff fc 20 22 00 01 34 01 00 00
@00001b0  44 41 00 0a 2b 61 ff fc 34 21 ff fd 00 21 00 01
@00001c0  5b 61 00 00 2b 62 00 00 34 01 00 3f 54 41 00 0b
@00001d0  2b 61 00 00 fb ff ff 9b 2b 61 ff f8 b4 21 08 00
@00001e0  b8 20 10 00 2b 61 ff fc b4 41 08 00 34 21 00 03
@00001f0  5b 61 ff fc e3 ff ff ec 2b 61 ff f8 34 21 00 01
@0000200  5b 61 ff f8 2b 62 ff f8 34 01 00 3f 50 22 ff d9
@0000210  34 01 00 00 2b 9b 00 08 2b 9d 00 04 37 9c 00 14
@0000220  c3 a0 00 00                                    
