/*
:name: vector_vectored
:description: vectored vector tests
:should_fail: 0
:tags: 6.9.2
*/
module top();
	tri1 vectored [15:0] a;

endmodule
