/*
:name: class_member_test_10
:description: Test
:should_fail: 0
:tags: 8.3
*/
class outerclass;
  class innerclass;
    class reallyinnerclass;
      task subtask;
      endtask
    endclass
  endclass
endclass