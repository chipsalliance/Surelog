/*
:name: 22.9--unconnected_drive-invalid-2
:description: Test
:should_fail_because: the directive `unconnected_drive takes one of two arguments: pull1 or pull0
:tags: 22.9
:type: preprocessing
*/
`unconnected_drive pull2
`nounconnected_drive
