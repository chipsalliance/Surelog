/*
:name: unconnected-drive
:description: Unconnected drive keywords
:should_fail: 0
:tags: 5.6.4
*/


`unconnected_drive pull1

module ts();
endmodule

`nounconnected_drive
