
`default_nettype wire


module dumb();

endmodule
