/*
:name: iface_class_test_5
:description: Test
:should_fail: 0
:tags: 8.3 8.26
*/
interface class base_ic #(int N = 8) extends pkg1::base1, base2#(N);
endclass