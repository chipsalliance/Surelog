module top();

logic [10:0] product_exponent;

assign p = product_exponent[7:0] == '1;

endmodule // top

