/*
:name: 22.7--timescale-basic-3
:description: Test
:should_fail: 1
:tags: 22.7
:type: simulation
*/
`timescale 9 ns / 1 ps
