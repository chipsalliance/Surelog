/*
:name: typedef_test_19
:description: Test
:tags: 6.18
*/
typedef enum logic {
  Global = 4'h2,
  Local = 4'h3
} myenum_fwd;