// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: defs 
:description: Utility for testing `include directive
:type: preprocessing
:tags: 22.4
*/

`define define_var "define_var"
`define TWO_PLUS_TWO 5
