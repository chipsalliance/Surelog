/*
:name: include-directive
:description: Include empty file
:tags: 5.6.4
*/

`include "/dev/null"

module empty();
endmodule
