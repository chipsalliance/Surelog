/*
:name: desc_test_11
:description: Test
:type: preprocessing
:should_fail: 0
:tags: 5.6.4
*/
`ifdef DEBUGGER
`MACRO(stuff, morestuff)
`endif
