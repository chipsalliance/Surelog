/*
:name: default-nettype
:description: Default nettype check
:should_fail: 0
:tags: 5.6.4
*/

`default_nettype wire
`default_nettype none
module dn();
endmodule
