/*
:name: 22.5.1--define
:description: Test
:tags: 22.5.1
:type: preprocessing
*/
`define FOUR 5
`define SOMESTRING "somestring"
