/*
:name: desc_test_3
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
`else
`endif
