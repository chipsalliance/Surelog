/*
:name: class_member_test_7
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern virtual protected task subtask(arg_type arg);
endclass