module top(b,c);
input b;
output c;

assign c = b;
endmodule
