/*
:name: debug-line
:description: Debugging compiler directives
:should_fail: 0
:tags: 5.6.4
*/

module directives();
  `line 1 "5.6.4--compiler-directives-debug-line.sv" 1
endmodule
