/*
:name: localparam
:description: localparam tests
:tags: 6.20.4
*/
module top();
	localparam p = 123;
endmodule
