// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: variable_assignment
:description: Variable assignment tests
:tags: 6.5
*/
module top();
	int v;

	assign v = 12;
endmodule
