/*
:name: class_test_47
:description: Test
:tags: 6.15 8.3
*/
class macros_id_as_call;
 `uvm_new_func
 `uvm_new_func2  // comment
 `uvm_new_func3  /* comment */
endclass