/*
:name: comments
:description: A module testing system verilog comments
:tags: 5.4
*/
module empty (
);
  /* multi
     line
     comment
   */

  // single line comment
endmodule
