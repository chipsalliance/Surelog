/*
:name: nettype
:description: user-defined nettype tests
:should_fail: 0
:tags: 6.6.7
*/
module top();
	nettype real real_net;
endmodule
