
/*
 * Copyright (c) 2000 Peter monta (pmonta@pacbell.net)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */
// Reworked slightly to be self checking.
module main;

  wire y;
  reg  a,b;
  reg  error;

  assign y = a && (b ? 0 : 1);

  initial 
    begin
       error = 0;
       #1 ; // get passed the time 0 race problems ;-)
       b = 1;
       a = 1;
       #1 ;
       if(y !== 0)
         begin
           $display("FAILED");
           error = 1;
         end   
       #1 ;
       b = 0;
       #1 ;
       if(y !== 1)
         begin
           $display("FAILED");
           error = 1;
         end   
       if(error === 0)
         $display("PASSED");
    end

endmodule
