/*
:name: 22.11--pragma-nested
:description: Test
:should_fail: 0
:tags: 22.11
:type: preprocessing
*/
`pragma foo something, somethingelse = 7, "abcdef", ( hello, ( "world", pr = 4, "gm" ) ), a
