/*
:name: typedef_test_11
:description: Test
:tags: 6.18
*/
typedef bit data_t;

typedef data_t my_array_t [bit];
