// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: debug-line
:description: Debugging compiler directives
:tags: 5.6.4
*/

module directives();
  `line 1 "5.6.4--compiler-directives-debug-line.sv" 1
endmodule
