`define DDR_ANA_DQS_DRVR_LPBK_NCAL_FIELD          4:0
`define DDR_ANA_DQS_DRVR_LPBK_PCAL_FIELD          10:5
`define DDR_ANA_DQS_DRVR_LPBK_BS_EN_FIELD         11
`define DDR_ANA_DQS_DRVR_LPBK_LPBK_EN_FIELD       12
`define DDR_ANA_DQS_DRVR_LPBK_SE_MODE_FIELD       13
