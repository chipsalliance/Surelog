/*
:name: dummy_include
:description: Utility for testing `include directive
:type: preprocessing
:should_fail: 0
:tags: 22.4
*/
