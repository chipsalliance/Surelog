/*
:name: class_test_8
:description: Test
:tags: 6.15 8.3
*/
class Foo extends Bar #(x,y,z); endclass