/*
:name: class_test_12
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo #(int N=1, int P=2) extends Bar #(x,y,z);
endclass