
// Benchmark source:
// https://github.com/jamesbowman/swapforth/tree/master/j1a

// ===================================================================

`timescale 1 ns / 1 ps

`default_nettype none
`define WIDTH 16

module SB_RAM2048x2(
	output [1:0] RDATA,
	input        RCLK, RCLKE, RE,
	input  [10:0] RADDR,
	input         WCLK, WCLKE, WE,
	input  [10:0] WADDR,
	input  [1:0] MASK, WDATA
);
	parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  wire [15:0] rd;

  SB_RAM40_4K #(
    .WRITE_MODE(3),
    .READ_MODE(3),
    .INIT_0(INIT_0),
    .INIT_1(INIT_1),
    .INIT_2(INIT_2),
    .INIT_3(INIT_3),
    .INIT_4(INIT_4),
    .INIT_5(INIT_5),
    .INIT_6(INIT_6),
    .INIT_7(INIT_7),
    .INIT_8(INIT_8),
    .INIT_9(INIT_9),
    .INIT_A(INIT_A),
    .INIT_B(INIT_B),
    .INIT_C(INIT_C),
    .INIT_D(INIT_D),
    .INIT_E(INIT_E),
    .INIT_F(INIT_F)
  ) _ram (
    .RDATA(rd),
    .RADDR(RADDR),
    .RCLK(RCLK), .RCLKE(RCLKE), .RE(RE),
    .WCLK(WCLK), .WCLKE(WCLKE), .WE(WE),
    .WADDR(WADDR),
    .MASK(16'h0000), .WDATA({4'b0, WDATA[1], 7'b0, WDATA[0], 3'b0}));

  assign RDATA[0] = rd[3];
  assign RDATA[1] = rd[11];

endmodule

module ioport(
  input clk,
  inout [7:0] pins,
  input we,
  input [7:0] wd,
  output [7:0] rd,
  input [7:0] dir);

  genvar i;
  generate 
    for (i = 0; i < 8; i = i + 1) begin : io
      // 1001   PIN_OUTPUT_REGISTERED_ENABLE 
      //     01 PIN_INPUT 
      SB_IO #(.PIN_TYPE(6'b1001_01)) _io (
        .PACKAGE_PIN(pins[i]),
        .CLOCK_ENABLE(we),
        .OUTPUT_CLK(clk),
        .D_OUT_0(wd[i]),
        .D_IN_0(rd[i]),
        .OUTPUT_ENABLE(dir[i]));
    end
  endgenerate

endmodule

module outpin(
  input clk,
  output pin,
  input we,
  input wd,
  output rd);

  SB_IO #(.PIN_TYPE(6'b0101_01)) _io (
        .PACKAGE_PIN(pin),
        .CLOCK_ENABLE(we),
        .OUTPUT_CLK(clk),
        .D_OUT_0(wd),
        .D_IN_0(rd));
endmodule

module inpin(
  input clk,
  input pin,
  output rd);

  SB_IO #(.PIN_TYPE(6'b0000_00)) _io (
        .PACKAGE_PIN(pin),
        .INPUT_CLK(clk),
        .D_IN_0(rd));
endmodule

module top(input pclk, output D1, output D2, output D3, output D4, output D5,

           output TXD,        // UART TX
           input RXD,         // UART RX

           output PIOS_00,    // flash SCK
           input PIOS_01,     // flash MISO
           output PIOS_02,    // flash MOSI
           output PIOS_03,    // flash CS

           inout PIO1_02,    // PMOD 1
           inout PIO1_03,    // PMOD 2
           inout PIO1_04,    // PMOD 3
           inout PIO1_05,    // PMOD 4
           inout PIO1_06,    // PMOD 5
           inout PIO1_07,    // PMOD 6
           inout PIO1_08,    // PMOD 7
           inout PIO1_09,    // PMOD 8

           inout PIO0_02,    // HDR1 1
           inout PIO0_03,    // HDR1 2
           inout PIO0_04,    // HDR1 3
           inout PIO0_05,    // HDR1 4
           inout PIO0_06,    // HDR1 5
           inout PIO0_07,    // HDR1 6
           inout PIO0_08,    // HDR1 7
           inout PIO0_09,    // HDR1 8

           inout PIO2_10,    // HDR2 1
           inout PIO2_11,    // HDR2 2
           inout PIO2_12,    // HDR2 3
           inout PIO2_13,    // HDR2 4
           inout PIO2_14,    // HDR2 5
           inout PIO2_15,    // HDR2 6
           inout PIO2_16,    // HDR2 7
           inout PIO2_17,    // HDR2 8

           output PIO1_18,    // IR TXD
           input  PIO1_19,    // IR RXD
           output PIO1_20,    // IR SD

           input resetq
);
  localparam MHZ = 12;

  wire clk;
  SB_PLL40_CORE #(.FEEDBACK_PATH("SIMPLE"),
                  .PLLOUT_SELECT("GENCLK"),
                  .DIVR(4'b0000),
                  .DIVF(7'd3),
                  .DIVQ(3'b000),
                  .FILTER_RANGE(3'b001)
                 ) uut (
                         .REFERENCECLK(pclk),
                         .PLLOUTCORE(clk),
                         //.PLLOUTGLOBAL(clk),
                         // .LOCK(D5),
                         .RESETB(1'b1),
                         .BYPASS(1'b0)
                        );

  wire io_rd, io_wr;
  wire [15:0] mem_addr;
  wire mem_wr;
  wire [15:0] dout;
  wire [15:0] io_din;
  wire [12:0] code_addr;
  reg unlocked = 0;

    wire [15:0] insn0, insn1;
    wire [15:0] insn;

  SB_RAM2048x2 #(
    .INIT_0(256'h5356015230330c46360b2c394049315a400a23690e673f1b3576526a65064505),
    .INIT_1(256'h712a2c5c5339654e2c5806594615236c4549245e0c1b4f465c340d35727f260d),
    .INIT_2(256'h2060281a774c362c0b3f061e0861017c48510c00045c2d716c60045433615f76),
    .INIT_3(256'h0d1613131b730265441e11214e264b4237166b6a4366447c2d5c2f1e163a413b),
    .INIT_4(256'h6c584c642b1f3a55327a0e357b2d29040104003d140202786b13015f0d313157),
    .INIT_5(256'h5c6645571931347c0030653c7c0b1846307f4b7d215a335c3557483e64692e08),
    .INIT_6(256'h24190f13193841541153505e124a545c192c612b48410444706675554a252877),
    .INIT_7(256'h345d292c797c5830602d280c0c7d684806757c0a2d202e72041a3a00083c413f),
    .INIT_8(256'h401004186404393c6040085d244d0c6975742534216c7c342c7d5008352d0460),
    .INIT_9(256'h0019200c3818010d651048254d51452d1c04641d401c405d38241c1914442829),
    .INIT_A(256'h08100515243c11140820002015382d3c21343034200435153130081911252925),
    .INIT_B(256'h04300511203d0031382c1018303d110c252d0010001511102024251d003c0109),
    .INIT_C(256'h3000331410083c3f303c3d0b011b0913231e2414061e0c173d0032262b043614),
    .INIT_D(256'h330b3e24241d04362c1b30180905340d260e0232241b022c331f120c1a02111c),
    .INIT_E(256'h0a271c192e3210201a16043e38040a0f10373429362e020a3c261a2c33252f37),
    .INIT_F(256'h080b213e1d21130a302f191d160712261825161e3325351811241031151e3c16)
  ) _bn00 (
    .RDATA(insn0[1:0]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[1:0]));

  SB_RAM2048x2 #(
    .INIT_0(256'h30300105082d462c203d2c28366752136a5b7327081e154e387e0e02156f7870),
    .INIT_1(256'h005c100c653b1c08092914216c1f72335555101045291804296b073f4a4a0129),
    .INIT_2(256'h486a515100502020332b423240681071486830280919243c195d71313a382109),
    .INIT_3(256'h223b7571442c0c6e217511311602051d424252101b223a2e6b7d001221104535),
    .INIT_4(256'h1246046c7850024a161f65760858520b214119695c180a7a5b53245613250636),
    .INIT_5(256'h30266064055300741c5c5450407a564d614a0a1c60510b1f09477b5134724848),
    .INIT_6(256'h08072c3424356c7d0a48521c0000287a2070475528735033595a5b390f041a10),
    .INIT_7(256'h6001697008281c147d7c4160303416156b193611550a0f3b3c322a3c241c6635),
    .INIT_8(256'h6d7d147c054554544918150c5554054109484c4c3838150d4130707020782c30),
    .INIT_9(256'h143410302c2c28381d182020243c0125217029087c5924605c51657441101c5c),
    .INIT_A(256'h3d2c0c0d1414280c041401202408002530142425293c3c0c3435292808340015),
    .INIT_B(256'h1c1c0804301c0c29252c01212131241c283c2c343014151439390039003d1414),
    .INIT_C(256'h00092931292b0913221a000d29091030383a19333a3a242f0c3e2a2b2203012f),
    .INIT_D(256'h212310010a09112705132012012a22330811233b3d30042818393c362e370a18),
    .INIT_E(256'h390b321e00020607101904053b03111517360404082c1c1b3c0d030221091838),
    .INIT_F(256'h273e0d181c110d1c1c1c14142021040e01113a3c143c06211b123c14381e0c0f)
  ) _bn01 (
    .RDATA(insn0[3:2]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[3:2]));

  SB_RAM2048x2 #(
    .INIT_0(256'h143028722022020051540904633a505e1052161c46404f504a004e0030310203),
    .INIT_1(256'h14447d775226242a296005486618414c2c64307a0b05201004672c3848444526),
    .INIT_2(256'h224863355008424b0820223b2848001c59081c4c09613454410d787016447109),
    .INIT_3(256'h090b70087919421e351e1020122705051a0223021b3614283d210646043d003c),
    .INIT_4(256'h701648090a1b7a395f0549286d65342665471d0d10490a0832382c1415063e6a),
    .INIT_5(256'h1e314670596d7648103d233c1827135f315811571866682c06183a3e64317033),
    .INIT_6(256'h033a08743802797452065a0048051800586c3f5303023a1251146202003d5a17),
    .INIT_7(256'h784051686044201c010d210454781337695a52765a572a54003d3c523d01676a),
    .INIT_8(256'h4834251051501c0c480c1d750149082048000105184c191979595d6011601175),
    .INIT_9(256'h311c11152904203c5c5000751830645830314819047c0435741d6c6958684865),
    .INIT_A(256'h3111041c2439082030013511200c04102010000519013c0438290d3114001919),
    .INIT_B(256'h1c300511211824003d042c3c240d110504080c182810180d342c21200939010c),
    .INIT_C(256'h1838180c08331801300b2d3e291e0c1e221e2a180a1029001b1138140b3f0e2e),
    .INIT_D(256'h05040b223a2a3708362104011b0c31293a3a2a392d331e153904340529090929),
    .INIT_E(256'h2e350205212d0b362204240400260c011502040329090f0c3002072132161a3a),
    .INIT_F(256'h19133c2a3d0a040c110e010718300324192b0e093828012f0c392d2c1c000a01)
  ) _bn02 (
    .RDATA(insn0[5:4]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[5:4]));

  SB_RAM2048x2 #(
    .INIT_0(256'h3014082800200402104124050203005000102316004c1054304a044e24317b0a),
    .INIT_1(256'h1010045433100020002300011000300011200020000208082408032802480004),
    .INIT_2(256'h0000507000100021231012220020101100302018002800201000094830100020),
    .INIT_3(256'h280101741c70024004252118421600280a1a1021221200120010000000313500),
    .INIT_4(256'h06380c082047285a005f0449324910200861005064544042097a10214413003c),
    .INIT_5(256'h101a0002094102400034620710422033003f0c5720106546194a006b00001a60),
    .INIT_6(256'h303b1c600f0b60680258005a004932025008326c401358120950134040094a48),
    .INIT_7(256'h0070213d08411c387041602100481411106942340157190e002d0a5620350245),
    .INIT_8(256'h116804046451401c4808101534014c080008400920104d010059000870211819),
    .INIT_9(256'h2900301021201828440060000024084011604041784c402401544c3958082048),
    .INIT_A(256'h24090c00240105040120142d0c20000121002100200114282008040d14001410),
    .INIT_B(256'h001c20250029082400311d2c0434150c0034380428080c152d34200828051001),
    .INIT_C(256'h3e2e23081912000a0820143802230c08092a290208222c05263b160c022b030c),
    .INIT_D(256'h30312a2120122112211200241a213021321811082128203a2018221426091607),
    .INIT_E(256'h153e10022c2d1a193a2a25253b38190c01050004183130252c280106112a282a),
    .INIT_F(256'h251025350c1c25051011302108180109181c3000283c0706131d1c240018250b)
  ) _bn03 (
    .RDATA(insn0[7:6]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[7:6]));

  SB_RAM2048x2 #(
    .INIT_0(256'h1c73400240702b282002222801490b3e2e0a411c005e301e222146640b70654e),
    .INIT_1(256'h2000205e55304848517d226a7319082a0b09242c00082442421840481818380a),
    .INIT_2(256'h446808542e4a661c624a1011494a00162442047a495a480a0862210211074a0a),
    .INIT_3(256'h62562029060264356206232128350e022001601a2c3c7c68101c3c426e4a303c),
    .INIT_4(256'h297a0a757c581c0020122b6c06483c7a0c22262060010010606352323e212c11),
    .INIT_5(256'h3c694b3f07310a7d04791418545a64546d7a786e715610464805404c00401a45),
    .INIT_6(256'h284d19314218444c090d4241424c0a00343c4c2004031d07263602010c3c2068),
    .INIT_7(256'h01211018103040243c3c000c682c3046503f0431441016311e780a10241c440c),
    .INIT_8(256'h10701058082c3d1808050428507c4428346c480861252c20040c082014156821),
    .INIT_9(256'h082c1424001c00280400483c096d081c04204000042804204c1804201c140034),
    .INIT_A(256'h0029281914313000080828081d1800153010142c01200128000900381d181c38),
    .INIT_B(256'h0018381d3c3c0114201904082925101c2c38181430342809383c1439283d2009),
    .INIT_C(256'h082700390c2b0d3f2839000910263d30303b3b323a381e2a0e390602023b100c),
    .INIT_D(256'h122a0b2a0506003d1211002502123511141c101d30180203303b062b083a0533),
    .INIT_E(256'h0e1908030c3a0a1f190e1c31083a2e180602380e0c3830070d25120720330821),
    .INIT_F(256'h020a142218070a182e3a050f0f2834170c1210150d200212021c0812110d000d)
  ) _bn04 (
    .RDATA(insn0[9:8]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[9:8]));

  SB_RAM2048x2 #(
    .INIT_0(256'h10180044025406072202203100110b212204304c203020141034282a240d442d),
    .INIT_1(256'h2125200000404850552431252040080000072228023422120040015908282010),
    .INIT_2(256'h44000040282030403160240043010220261026384b0d12042208220504050054),
    .INIT_3(256'h2204100664600440221041432010001814013040044038500010000038400100),
    .INIT_4(256'h2124100030001412005620511108014140481010201000123002004010102508),
    .INIT_5(256'h20000040010149000020504000004400401109286002004010400004080a042c),
    .INIT_6(256'h7344012e00404450405003030a1a1c4c644810400106050c0400101404000060),
    .INIT_7(256'h04341030181850404c50000020400a0a03620829024001015062001804041454),
    .INIT_8(256'h48285000406c1010101810004030004000200040405400300018001004257048),
    .INIT_9(256'h0020042000000130000000640038000000200000007008280048407000041028),
    .INIT_A(256'h0021002110200000202000181131202830000c00002001390800080800000018),
    .INIT_B(256'h080414011109100530200010011000003c050400100000243030102010010029),
    .INIT_C(256'h0121002004000100000000000001100030001001102010221029000102220008),
    .INIT_D(256'h0a2a042c10101030000802301000000000110008100000081818183000381101),
    .INIT_E(256'h1a0a1a1010381001000018201028300002000804160e10050525000212000426),
    .INIT_F(256'h02000020001018001a0004110000141010000000003200001200021001081002)
  ) _bn05 (
    .RDATA(insn0[11:10]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[11:10]));

  SB_RAM2048x2 #(
    .INIT_0(256'h671156007a0027200200210159002f300e007d0036600e0077436a224e123400),
    .INIT_1(256'h21010a5061004a0075106b0041003c001f006e042a02430174007b203e001800),
    .INIT_2(256'h76000c006f215c006b0025006b212e0016007e007f014b01720007006f047620),
    .INIT_3(256'h36042b20670075004a400300390c5610652158004410780014007b214a000d00),
    .INIT_4(256'h631077001100171072427f404908692832003200111012122302230039085500),
    .INIT_5(256'h69001f0233017d00415039000900441051003b10570110100500060a420a2560),
    .INIT_6(256'h4705430254004448450043405f426d402c000c080f0927002e121d0034002400),
    .INIT_7(256'h050110083c1044213d004c0024004c000528091062106302530050011d005c00),
    .INIT_8(256'h4900580004007100140068005c00240074084000650024000c0008080d086100),
    .INIT_9(256'h200004001100050004003d404100140004001000300019000010040004002908),
    .INIT_A(256'h05003100380010003c08202031203c0010003c00110119000c0018000d002000),
    .INIT_B(256'h2c101d081504190028002120292020200d002500140030103120150009003901),
    .INIT_C(256'h210010080500350011000308370133011402170216021602210107011e021904),
    .INIT_D(256'h03090501150318001b02130004000d00070908001a000b021f00190016102100),
    .INIT_E(256'h0f001b083200210115011c08070037040700371c062413012701321407000702),
    .INIT_F(256'h2e00321013101a002b011f01070136000200350033001800220c12001d101e10)
  ) _bn06 (
    .RDATA(insn0[13:12]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[13:12]));

  SB_RAM2048x2 #(
    .INIT_0(256'h10660014007a5037005e403d004d007f4006003f015e000e0076104a005d0035),
    .INIT_1(256'h0278005a003f015a006c006b0009107c4017017e403a004a0038006f413e4018),
    .INIT_2(256'h316e005c004e001c046b422d1462007e0056017a007e006a0072004710690026),
    .INIT_3(256'h4036002b006f007e005e040322350052026504180254217e421c007c004e420d),
    .INIT_4(256'h00730877005408030072007f004d006d10260036421d055a044b006744300051),
    .INIT_5(256'h1065007f013f007d005d001c00290076007f005d085700562845006e205b0075),
    .INIT_6(256'h204f0863305c407c205f2047005d016c012c102a007f1067403e403d0074007f),
    .INIT_7(256'h00754438002c012c003c106d012c106c003d007f003e007f107f2950407c003b),
    .INIT_8(256'h007d315c000400752814006c007d1168017c3408006d0874205c4538005d1461),
    .INIT_9(256'h00141924003c000d2110005d0075215408556419014c0075205500112954100d),
    .INIT_A(256'h002d003900180034003d00240030003c081c003d00340008001c003c00291124),
    .INIT_B(256'h013c003d0035001900280429003d003c100d0134101d00302039000d0025203d),
    .INIT_C(256'h0806003a001f003f043b001f003d0837001e001f2116003a08050023023e003f),
    .INIT_D(256'h1409100500140418001f0c33000c200d102d041a301e042b003f001d00360021),
    .INIT_E(256'h002b201700060025001c0200002700370826002f0022003308060826002f0807),
    .INIT_F(256'h002e001b0837201f002f201f0026003e0826003d0817003d002f003e201e003e)
  ) _bn07 (
    .RDATA(insn0[15:14]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[15:14]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn10 (
    .RDATA(insn1[1:0]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[1:0]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn11 (
    .RDATA(insn1[3:2]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[3:2]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn12 (
    .RDATA(insn1[5:4]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[5:4]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn13 (
    .RDATA(insn1[7:6]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[7:6]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn14 (
    .RDATA(insn1[9:8]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[9:8]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn15 (
    .RDATA(insn1[11:10]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[11:10]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn16 (
    .RDATA(insn1[13:12]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[13:12]));

  SB_RAM2048x2 #(
    .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
  ) _bn17 (
    .RDATA(insn1[15:14]),
    .RADDR(code_addr[10:0]),
    .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
    .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]),
    .WADDR(mem_addr[11:1]),
    .MASK(16'h0000), .WDATA(dout[15:14]));

    reg c11;
    always @(posedge clk) c11 <= code_addr[11];
    wire [15:0] cm = {16{c11}};
    assign insn = (cm & insn1) | (~cm & insn0);
    // assign insn = c11 ? insn1 : insn0;

  j1 _j1(
    .clk(clk),
    .resetq(resetq),
    .io_rd(io_rd),
    .io_wr(io_wr),
    .mem_wr(mem_wr),
    .dout(dout),
    .io_din(io_din),
    .mem_addr(mem_addr),
    .code_addr(code_addr),
    .insn(insn));

  /*
  // ######   TICKS   #########################################

  reg [15:0] ticks;
  always @(posedge clk)
    ticks <= ticks + 16'd1;
  */

  // ######   IO SIGNALS   ####################################

`define EASE_IO_TIMING
`ifdef EASE_IO_TIMING
  reg io_wr_, io_rd_;
  reg [15:0] dout_;
  reg [15:0] io_addr_;

  always @(posedge clk) begin
    {io_rd_, io_wr_, dout_} <= {io_rd, io_wr, dout};
    if (io_rd | io_wr)
      io_addr_ <= mem_addr;
  end
`else
  wire io_wr_ = io_wr, io_rd_ = io_rd;
  wire [15:0] dout_ = dout;
  wire [15:0] io_addr_ = mem_addr;
`endif

  // ######   PMOD   ##########################################

  reg [7:0] pmod_dir;   // 1:output, 0:input
  wire [7:0] pmod_in;

  ioport _mod (.clk(clk),
               .pins({PIO1_09, PIO1_08, PIO1_07, PIO1_06, PIO1_05, PIO1_04, PIO1_03, PIO1_02}),
               .we(io_wr_ & io_addr_[0]),
               .wd(dout_),
               .rd(pmod_in),
               .dir(pmod_dir));

  // ######   HDR1   ##########################################

  reg [7:0] hdr1_dir;   // 1:output, 0:input
  wire [7:0] hdr1_in;

  ioport _hdr1 (.clk(clk),
               .pins({PIO0_09, PIO0_08, PIO0_07, PIO0_06, PIO0_05, PIO0_04, PIO0_03, PIO0_02}),
               .we(io_wr_ & io_addr_[4]),
               .wd(dout_[7:0]),
               .rd(hdr1_in),
               .dir(hdr1_dir));

  // ######   HDR2   ##########################################

  reg [7:0] hdr2_dir;   // 1:output, 0:input
  wire [7:0] hdr2_in;

  ioport _hdr2 (.clk(clk),
               .pins({PIO2_17, PIO2_16, PIO2_15, PIO2_14, PIO2_13, PIO2_12, PIO2_11, PIO2_10}),
               .we(io_wr_ & io_addr_[6]),
               .wd(dout_[7:0]),
               .rd(hdr2_in),
               .dir(hdr2_dir));

  // ######   UART   ##########################################

  wire uart0_valid, uart0_busy;
  wire [7:0] uart0_data;
  wire uart0_wr = io_wr_ & io_addr_[12];
  wire uart0_rd = io_rd_ & io_addr_[12];
  wire uart_RXD;
  inpin _rcxd(.clk(clk), .pin(RXD), .rd(uart_RXD));
  buart _uart0 (
     .clk(clk),
     .resetq(1'b1),
     .rx(uart_RXD),
     .tx(TXD),
     .rd(uart0_rd),
     .wr(uart0_wr),
     .valid(uart0_valid),
     .busy(uart0_busy),
     .tx_data(dout_[7:0]),
     .rx_data(uart0_data));

  wire [4:0] LEDS;
  wire w4 = io_wr_ & io_addr_[2];

  outpin led0 (.clk(clk), .we(w4), .pin(D5), .wd(dout_[0]), .rd(LEDS[0]));
  outpin led1 (.clk(clk), .we(w4), .pin(D4), .wd(dout_[1]), .rd(LEDS[1]));
  outpin led2 (.clk(clk), .we(w4), .pin(D3), .wd(dout_[2]), .rd(LEDS[2]));
  outpin led3 (.clk(clk), .we(w4), .pin(D2), .wd(dout_[3]), .rd(LEDS[3]));
  outpin led4 (.clk(clk), .we(w4), .pin(D1), .wd(dout_[4]), .rd(LEDS[4]));

  wire [4:0] PIOS;
  wire w8 = io_wr_ & io_addr_[3];

  outpin pio0 (.clk(clk), .we(w8), .pin(PIOS_03), .wd(dout_[0]), .rd(PIOS[0]));
  outpin pio1 (.clk(clk), .we(w8), .pin(PIOS_02), .wd(dout_[1]), .rd(PIOS[1]));
  outpin pio2 (.clk(clk), .we(w8), .pin(PIOS_00), .wd(dout_[2]), .rd(PIOS[2]));
  outpin pio3 (.clk(clk), .we(w8), .pin(PIO1_18), .wd(dout_[3]), .rd(PIOS[3]));
  outpin pio4 (.clk(clk), .we(w8), .pin(PIO1_20), .wd(dout_[4]), .rd(PIOS[4]));

  // ######   RING OSCILLATOR   ###############################

  wire [1:0] buffers_in, buffers_out;
  assign buffers_in = {buffers_out[0:0], ~buffers_out[1]};
  SB_LUT4 #(
          .LUT_INIT(16'd2)
  ) buffers [1:0] (
          .O(buffers_out),
          .I0(buffers_in),
          .I1(1'b0),
          .I2(1'b0),
          .I3(1'b0)
  );
  wire random = 0; // ~buffers_out[1];

  // ######   IO PORTS   ######################################

  /*        bit   mode    device
      0001  0     r/w     PMOD GPIO
      0002  1     r/w     PMOD direction
      0004  2     r/w     LEDS
      0008  3     r/w     misc.out
      0010  4     r/w     HDR1 GPIO
      0020  5     r/w     HDR1 direction
      0040  6     r/w     HDR2 GPIO
      0080  7     r/w     HDR2 direction
      0800  11      w     sb_warmboot
      1000  12    r/w     UART RX, UART TX
      2000  13    r       misc.in
  */

  assign io_din =
    (io_addr_[ 0] ? {8'd0, pmod_in}                                     : 16'd0) |
    (io_addr_[ 1] ? {8'd0, pmod_dir}                                    : 16'd0) |
    (io_addr_[ 2] ? {11'd0, LEDS}                                       : 16'd0) |
    (io_addr_[ 3] ? {11'd0, PIOS}                                       : 16'd0) |
    (io_addr_[ 4] ? {8'd0, hdr1_in}                                     : 16'd0) |
    (io_addr_[ 5] ? {8'd0, hdr1_dir}                                    : 16'd0) |
    (io_addr_[ 6] ? {8'd0, hdr2_in}                                     : 16'd0) |
    (io_addr_[ 7] ? {8'd0, hdr2_dir}                                    : 16'd0) |
    (io_addr_[12] ? {8'd0, uart0_data}                                  : 16'd0) |
    (io_addr_[13] ? {11'd0, random, PIO1_19, PIOS_01, uart0_valid, !uart0_busy} : 16'd0);

  reg boot, s0, s1;

  SB_WARMBOOT _sb_warmboot (
    .BOOT(boot),
    .S0(s0),
    .S1(s1)
    );

  always @(posedge clk) begin
    if (io_wr_ & io_addr_[1])
      pmod_dir <= dout_[7:0];
    if (io_wr_ & io_addr_[5])
      hdr1_dir <= dout_[7:0];
    if (io_wr_ & io_addr_[7])
      hdr2_dir <= dout_[7:0];
    if (io_wr_ & io_addr_[11])
      {boot, s1, s0} <= dout_[2:0];
  end

  always @(negedge resetq or posedge clk)
    if (!resetq)
      unlocked <= 0;
    else
      unlocked <= unlocked | io_wr_;

endmodule // top
`default_nettype none

`define CLKFREQ   12000000    // frequency of incoming signal 'clk'
`define BAUD      115200

// Simple baud generator for transmitter
// ser_clk pulses at 115200 Hz

module baudgen(
  input wire clk,
  output wire ser_clk);

  localparam lim = (`CLKFREQ / `BAUD) - 1; 
  localparam w = $clog2(lim);
  wire [w-1:0] limit = lim;
  reg [w-1:0] counter;
  assign ser_clk = (counter == limit);

  always @(posedge clk)
    counter <= ser_clk ? 0 : (counter + 1);
endmodule

// For receiver, a similar baud generator.
//
// Need to restart the counter when the transmission starts
// Generate 2X the baud rate to allow sampling on bit boundary
// So ser_clk pulses at 2*115200 Hz

module baudgen2(
  input wire clk,
  input wire restart,
  output wire ser_clk);

  localparam lim = (`CLKFREQ / (2 * `BAUD)) - 1; 
  localparam w = $clog2(lim);
  wire [w-1:0] limit = lim;
  reg [w-1:0] counter;
  assign ser_clk = (counter == limit);

  always @(posedge clk)
    if (restart)
      counter <= 0;
    else
      counter <= ser_clk ? 0 : (counter + 1);

endmodule

/*

-----+     +-----+-----+-----+-----+-----+-----+-----+-----+-----+-----+----
     |     |     |     |     |     |     |     |     |     |     |     |
     |start|  1  |  2  |  3  |  4  |  5  |  6  |  7  |  8  |stop1|stop2|
     |     |     |     |     |     |     |     |     |     |     |  ?  |
     +-----+-----+-----+-----+-----+-----+-----+-----+-----+           +

*/

module uart(
   input wire clk,
   input wire resetq,

   output wire uart_busy,       // High means UART is transmitting
   output reg uart_tx,          // UART transmit wire

   input wire uart_wr_i,        // Raise to transmit byte
   input wire [7:0] uart_dat_i
);
  reg [3:0] bitcount;           // 0 means idle, so this is a 1-based counter
  reg [8:0] shifter;

  assign uart_busy = |bitcount;
  wire sending = |bitcount;

  wire ser_clk;

  baudgen _baudgen(
    .clk(clk),
    .ser_clk(ser_clk));

  always @(negedge resetq or posedge clk)
  begin
    if (!resetq) begin
      uart_tx <= 1;
      bitcount <= 0;
      shifter <= 0;
    end else begin
      if (uart_wr_i) begin
        { shifter, uart_tx } <= { uart_dat_i[7:0], 1'b0, 1'b1 };
        bitcount <= 1 + 8 + 1;    // 1 start, 8 data, 1 stop
      end else if (ser_clk & sending) begin
        { shifter, uart_tx } <= { 1'b1, shifter };
        bitcount <= bitcount - 4'd1;
      end
    end
  end

endmodule

module rxuart(
   input wire clk,
   input wire resetq,
   input wire uart_rx,      // UART recv wire
   input wire rd,           // read strobe
   output wire valid,       // has data 
   output wire [7:0] data); // data
  reg [4:0] bitcount;
  reg [7:0] shifter;

  // bitcount == 11111: idle
  //             0-17:  sampling incoming bits
  //             18:    character received

  // On starting edge, wait 3 half-bits then sample, and sample every 2 bits thereafter

  wire idle = &bitcount;
  assign valid = (bitcount == 18);

  wire sample;
  reg [2:0] hh = 3'b111;
  wire [2:0] hhN = {hh[1:0], uart_rx};
  wire startbit = idle & (hhN[2:1] == 2'b10);
  wire [7:0] shifterN = sample ? {hh[1], shifter[7:1]} : shifter;

  wire ser_clk;

  baudgen2 _baudgen(
    .clk(clk),
    .restart(startbit),
    .ser_clk(ser_clk));

  reg [4:0] bitcountN;
  always @*
    if (startbit)
      bitcountN = 0;
    else if (!idle & !valid & ser_clk)
      bitcountN = bitcount + 5'd1;
    else if (valid & rd)
      bitcountN = 5'b11111;
    else
      bitcountN = bitcount;

  // 3,5,7,9,11,13,15,17
  assign sample = (|bitcount[4:1]) & bitcount[0] & ser_clk;
  assign data = shifter;

  always @(negedge resetq or posedge clk)
  begin
    if (!resetq) begin
      hh <= 3'b111;
      bitcount <= 5'b11111;
      shifter <= 0;
    end else begin
      hh <= hhN;
      bitcount <= bitcountN;
      shifter <= shifterN;
    end
  end
endmodule

module buart(
   input wire clk,
   input wire resetq,
   input wire rx,           // recv wire
   output wire tx,          // xmit wire
   input wire rd,           // read strobe
   input wire wr,           // write strobe
   output wire valid,       // has recv data 
   output wire busy,        // is transmitting
   input wire [7:0] tx_data,
   output wire [7:0] rx_data // data
);
  rxuart _rx (
     .clk(clk),
     .resetq(resetq),
     .uart_rx(rx),
     .rd(rd),
     .valid(valid),
     .data(rx_data));
  uart _tx (
     .clk(clk),
     .resetq(resetq),
     .uart_busy(busy),
     .uart_tx(tx),
     .uart_wr_i(wr),
     .uart_dat_i(tx_data));
endmodule
`default_nettype none
`define WIDTH 16

module j1(
  input wire clk,
  input wire resetq,

  output wire io_rd,
  output wire io_wr,
  output wire [15:0] mem_addr,
  output wire mem_wr,
  output wire [`WIDTH-1:0] dout,

  input  wire [`WIDTH-1:0] io_din,

  output wire [12:0] code_addr,
  input  wire [15:0] insn);

  reg [3:0] dsp, dspN;          // data stack pointer
  reg [`WIDTH-1:0] st0, st0N;   // top of data stack
  reg dstkW;                    // data stack write

  reg [12:0] pc /* verilator public_flat */, pcN;           // program counter
  wire [12:0] pc_plus_1 = pc + 13'd1;
  reg rstkW;                    // return stack write
  wire [`WIDTH-1:0] rstkD;      // return stack write value
  reg reboot = 1;

  assign mem_addr = st0[15:0];
  assign code_addr = pcN;

  // The D and R stacks
  wire [`WIDTH-1:0] st1, rst0;
  reg [1:0] dspI, rspI;
  stack2 #(.DEPTH(15)) dstack(.clk(clk), .rd(st1),  .we(dstkW), .wd(st0),   .delta(dspI));
  stack2 #(.DEPTH(17)) rstack(.clk(clk), .rd(rst0), .we(rstkW), .wd(rstkD), .delta(rspI));

  wire [16:0] minus = {1'b1, ~st0} + st1 + 1;
  wire signedless = st0[15] ^ st1[15] ? st1[15] : minus[16];

  always @*
  begin
    // Compute the new value of st0
    casez ({pc[12], insn[15:8]})
      9'b1_???_?????: st0N = insn;                    // literal
      9'b0_1??_?????: st0N = { {(`WIDTH - 15){1'b0}}, insn[14:0] };    // literal
      9'b0_000_?????: st0N = st0;                     // jump
      9'b0_010_?????: st0N = st0;                     // call
      9'b0_001_?????: st0N = st1;                     // conditional jump
      9'b0_011_?0000: st0N = st0;                     // ALU operations...
      9'b0_011_?0001: st0N = st1;
      9'b0_011_?0010: st0N = st0 + st1;
      9'b0_011_?0011: st0N = st0 & st1;
      9'b0_011_?0100: st0N = st0 | st1;
      9'b0_011_?0101: st0N = st0 ^ st1;
      9'b0_011_?0110: st0N = ~st0;

      9'b0_011_?0111: st0N = {`WIDTH{(minus == 0)}};                //  =
      9'b0_011_?1000: st0N = {`WIDTH{(signedless)}};                //  <

      9'b0_011_?1001: st0N = {st0[`WIDTH - 1], st0[`WIDTH - 1:1]};
      9'b0_011_?1010: st0N = {st0[`WIDTH - 2:0], 1'b0};
      9'b0_011_?1011: st0N = rst0;
      9'b0_011_?1100: st0N = minus[15:0];
      9'b0_011_?1101: st0N = io_din;
      9'b0_011_?1110: st0N = {{(`WIDTH - 4){1'b0}}, dsp};
      9'b0_011_?1111: st0N = {`WIDTH{(minus[16])}};                 // u<
      default: st0N = {`WIDTH{1'bx}};
    endcase
  end

  wire func_T_N =   (insn[6:4] == 1);
  wire func_T_R =   (insn[6:4] == 2);
  wire func_write = (insn[6:4] == 3);
  wire func_iow =   (insn[6:4] == 4);
  wire func_ior =   (insn[6:4] == 5);

  wire is_alu = !pc[12] & (insn[15:13] == 3'b011);
  assign mem_wr = !reboot & is_alu & func_write;
  assign dout = st1;
  assign io_wr = !reboot & is_alu & func_iow;
  assign io_rd = !reboot & is_alu & func_ior;

  assign rstkD = (insn[13] == 1'b0) ? {{(`WIDTH - 14){1'b0}}, pc_plus_1, 1'b0} : st0;

  always @*
  begin
    casez ({pc[12], insn[15:13]})
    4'b1_???,
    4'b0_1??:   {dstkW, dspI} = {1'b1,      2'b01};
    4'b0_001:   {dstkW, dspI} = {1'b0,      2'b11};
    4'b0_011:   {dstkW, dspI} = {func_T_N,  {insn[1:0]}};
    default:    {dstkW, dspI} = {1'b0,      2'b00};
    endcase
    dspN = dsp + {dspI[1], dspI[1], dspI};

    casez ({pc[12], insn[15:13]})
    4'b1_???:   {rstkW, rspI} = {1'b0,      2'b11};
    4'b0_010:   {rstkW, rspI} = {1'b1,      2'b01};
    4'b0_011:   {rstkW, rspI} = {func_T_R,  insn[3:2]};
    default:    {rstkW, rspI} = {1'b0,      2'b00};
    endcase

    casez ({reboot, pc[12], insn[15:13], insn[7], |st0})
    7'b1_0_???_?_?:   pcN = 0;
    7'b0_0_000_?_?,
    7'b0_0_010_?_?,
    7'b0_0_001_?_0:   pcN = insn[12:0];
    7'b0_1_???_?_?,
    7'b0_0_011_1_?:   pcN = rst0[13:1];
    default:          pcN = pc_plus_1;
    endcase
  end

  always @(negedge resetq or posedge clk)
  begin
    if (!resetq) begin
      reboot <= 1'b1;
      { pc, dsp, st0} <= 0;
    end else begin
      reboot <= 0;
      { pc, dsp, st0} <= { pcN, dspN, st0N };
    end
  end

endmodule
`default_nettype none
`define WIDTH 16

module stack2( 
  input wire clk,
  output wire [`WIDTH-1:0] rd,
  input wire we,
  input wire [1:0] delta,
  input wire [`WIDTH-1:0] wd);
  parameter DEPTH = 18;
  localparam BITS = (`WIDTH * DEPTH) - 1;

  wire move = delta[0];

  reg [15:0] head;
  reg [BITS:0] tail;
  wire [15:0] headN;
  wire [BITS:0] tailN;

  assign headN = we ? wd : tail[15:0];
  assign tailN = delta[1] ? {16'h55aa, tail[BITS:16]} : {tail[BITS-16:0], head};

  always @(posedge clk) begin
    if (we | move)
      head <= headN;
    if (move)
      tail <= tailN;
  end

  assign rd = head;

`ifdef VERILATOR
  int depth /* verilator public_flat */;
  always @(posedge clk) begin
    if (delta == 2'b11)
      depth <= depth - 1;
    if (delta == 2'b01)
      depth <= depth + 1;
  end
`endif

endmodule

