module top;
   int a [int];
   assign a[5] = 5;

   int b [string];
   assign b["HERE"] = 5;
endmodule
