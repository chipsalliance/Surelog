/*
:name: class_member_test_18
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function void subroutine(input bool x);
endclass