module top ();

endmodule

