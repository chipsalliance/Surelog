/*
:name: real-token
:description: Testing the real variable type
:should_fail: 0
:tags: 5.7.2
*/
module top();
  real a;
endmodule
