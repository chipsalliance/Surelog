/*
:name: class_test_2
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class static Foo; endclass