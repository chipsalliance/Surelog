/*
:name: stime_task
:description: $stime test
:should_fail: 0
:tags: 20.3
*/
module top();

initial
	$display($stime);

endmodule
