
module r5p_soc_top #(
  
  int unsigned GW = 32,

  int unsigned XLEN = 32
)(
  
);
endmodule
