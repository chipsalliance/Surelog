/*
:name: string_atoreal
:description: string.atoreal()  tests
:should_fail: 0
:tags: 6.16.10
*/
module top();
	string a = "4.76";
	real b = a.atoreal();
endmodule
