/*
:name: 22.12--line-illegal-1
:description: The level parameter shall be 0, 1, or 2
:should_fail: 1
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 3
