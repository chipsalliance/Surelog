/*
:name: class_member_test_25
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern virtual function integer subroutine;
endclass