// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: parameter_aggregate
:description: parameter aggregate type tests
:tags: 6.20.2
*/
module top();
	parameter logic [31:0] p [3:0] = '{1, 2, 3, 4};
endmodule
