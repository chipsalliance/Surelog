/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 13446
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_dqs_rcvr_no_esd_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath,
//View - schematic
// LAST TIME SAVED: Dec  7 16:22:35 2020
// NETLIST TIME: Dec 12 00:59:10 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath (out_cb, out_tb, vdda, vddq, vss, ena, 
    enb, in_c, in_t, se_ena, se_enb);

output  out_cb, out_tb;

inout  vdda, vddq, vss;

input  ena, enb, in_c, in_t, se_ena, se_enb;


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel INV4 ( .in(net1), .vss(vss), .out(net033), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel INV3 ( .in(net033), .vss(vss), .out(net1), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel INV2 ( .in(clk_b), .vss(vss), .out(clk), 
    .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel INV1 ( .in(clk), .vss(vss), .out(clk_b), 
    .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT PD ( .vss(vss), .enb(enb), .y(clk));

wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT PU0 ( .vdd(vddq), .en(ena), .y(clk_b));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV6 ( .in(net033), .vss(vss), .out(net2), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV5 ( .in(net1), .vss(vss), .out(net031), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT I1 ( .in(net034), .vss(vss), .out(net033), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV0 ( .in(net032), .vss(vss), .out(net1), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT6_2 ( .out(out_cb), .en(ena), .enb(enb), 
    .vss(vss), .in(net031), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT6_1 ( .out(out_cb), .en(ena), .enb(enb), 
    .vss(vss), .in(net031), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT6_0 ( .out(out_cb), .en(ena), .enb(enb), 
    .vss(vss), .in(net031), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT2 ( .out(net79), .en(se_ena), .enb(se_enb), 
    .vss(vss), .in(net80), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT4_1 ( .out(clk), .en(ena), .enb(enb), .vss(vss), 
    .in(net80), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT4_0 ( .out(clk), .en(ena), .enb(enb), .vss(vss), 
    .in(net80), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_1 ( .out(clk_b), .en(ena), .enb(enb), .vss(vss), 
    .in(net79), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_0 ( .out(clk_b), .en(ena), .enb(enb), .vss(vss), 
    .in(net79), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT5_2 ( .out(out_tb), .en(ena), .enb(enb), 
    .vss(vss), .in(net2), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT5_1 ( .out(out_tb), .en(ena), .enb(enb), 
    .vss(vss), .in(net2), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT5_0 ( .out(out_tb), .en(ena), .enb(enb), 
    .vss(vss), .in(net2), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_INVT INVT3 ( .out(net80), .en(vdda), .enb(vss), .vss(vss), 
    .in(in_t), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_INVT INVT0 ( .out(net79), .en(se_enb), .enb(se_ena), 
    .vss(vss), .in(in_c), .vdd(vddq));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT I0 ( .tielo(vss), .tiehi(vdda), .in(o_h_b), .vss(vss), 
    .out(net034), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT I2 ( .tielo(vss), .tiehi(vdda), .in(o_h), .vss(vss), 
    .out(net032), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath_lvlshift LVLSHIFT ( .out_cb(o_h), 
    .out_tb(o_h_b), .in_c(clk_b), .in_t(clk), .vss(vss), .vdda(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det, View -
//schematic
// LAST TIME SAVED: Dec 11 13:53:24 2020
// NETLIST TIME: Dec 12 00:59:10 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det (edge_det, edge_det_b, vdda, vddq, vss, byp, 
    ena, in, refsel);

output  edge_det, edge_det_b;

inout  vdda, vddq, vss;

input  byp, ena, in, refsel;


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det_sf Filter ( .out(net1), .ena(ena), .in(in), 
    .refsel(refsel), .vss(vss), .vddq(vddq), .vdda(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT PU0_1 ( .vdd(vdda), .en(pullupctrl), .y(net6));

wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT PU0_0 ( .vdd(vdda), .en(pullupctrl), .y(net6));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_LVT NOR1 ( .tielo(vss), .tiehi(vdda), .y(net4), .vss(vss), 
    .vdd(vdda), .b(byp), .a(ena));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_LVT NOR0 ( .tielo(vss), .tiehi(vdda), .y(net12), 
    .vss(vss), .vdd(vdda), .b(net1), .a(byp));

wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT PD0_1 ( .vss(vss), .enb(endge_det), .y(net6));

wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT PD0_0 ( .vss(vss), .enb(endge_det), .y(net6));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV13_1 ( .in(net3), .vss(vss), .out(edge_det_b), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV13_0 ( .in(net3), .vss(vss), .out(edge_det_b), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV12 ( .in(net4), .vss(vss), .out(pullupctrl), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV15_1 ( .in(edge_det_b), .vss(vss), .out(edge_det), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV15_0 ( .in(edge_det_b), .vss(vss), .out(edge_det), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_timing INV5 ( .in(net6), .vss(vss), .out(net3), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV2 ( .in(net12), .vss(vss), .out(endge_det), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT_timing INV4 ( .tielo(vss), .tiehi(vdda), .in(net3), .vss(vss), 
    .out(net6), .vdd(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell -
//wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay, View - schematic
// LAST TIME SAVED: Dec  7 15:38:07 2020
// NETLIST TIME: Dec 12 00:59:11 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay (out_c, out_t, vdda, vss, cal_ena, 
    cal_enb, dly_ctrl_c, dly_ctrl_t, ena, enb, in_c, in_t);

output  out_c, out_t;

inout  vdda, vss;

input  cal_ena, cal_enb, ena, enb, in_c, in_t;

input [3:0]  dly_ctrl_c;
input [3:0]  dly_ctrl_t;


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV1 ( .in(net6), .vss(vss), .out(out_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT INV0 ( .in(net2), .vss(vss), .out(out_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_5 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_4 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_3 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_2 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_1 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT0_0 ( .out(net8), .en(ena), .enb(enb), .vss(vss), 
    .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_5 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_4 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_3 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_2 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_1 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT INVT1_0 ( .out(net1), .en(ena), .enb(enb), .vss(vss), 
    .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT PU0 ( .vdd(vdda), .en(ena), .y(net1));

wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT PD0 ( .vss(vss), .enb(enb), .y(net8));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay_capdac CAPDAC_T ( .out(net2), 
    .dly_ctrl(dly_ctrl_t), .in(net8), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay_capdac CAPDAC_C ( .out(net6), 
    .dly_ctrl(dly_ctrl_c), .in(net1), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT_Mmod_nomodel INV5 ( .out(net1), .en(cal_enb), 
    .enb(cal_ena), .vss(vss), .in(net8), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT_Mmod_nomodel INV4 ( .out(net8), .en(cal_enb), 
    .enb(cal_ena), .vss(vss), .in(net1), .vdd(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath,
//View - schematic
// LAST TIME SAVED: Dec 11 22:28:06 2020
// NETLIST TIME: Dec 12 00:59:11 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath (out_cb, out_tb, vdda, vss, cal_cn, 
    cal_cp, cal_tn, cal_tp, dqs_in_c, dqs_in_t, ena, enb, fbctrl, 
    fbctrlb);

output  out_cb, out_tb;

inout  vdda, vss;

input  dqs_in_c, dqs_in_t, ena, enb;

input [2:0]  fbctrl;
input [3:0]  cal_tp;
input [3:0]  cal_tn;
input [2:0]  fbctrlb;
input [3:0]  cal_cp;
input [3:0]  cal_cn;


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_6 ( .out(out_tb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_5 ( .out(out_tb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_4 ( .out(out_tb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_3 ( .out(out_tb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_2 ( .out(out_tb), .ena(fbctrl[1]), 
    .enb(fbctrlb[1]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_1 ( .out(out_tb), .ena(fbctrl[1]), 
    .enb(fbctrlb[1]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_T_0 ( .out(out_tb), .ena(fbctrl[0]), 
    .enb(fbctrlb[0]), .in(in_t), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_6 ( .out(out_cb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_5 ( .out(out_cb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_4 ( .out(out_cb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_3 ( .out(out_cb), .ena(fbctrl[2]), 
    .enb(fbctrlb[2]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_2 ( .out(out_cb), .ena(fbctrl[1]), 
    .enb(fbctrlb[1]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_1 ( .out(out_cb), .ena(fbctrl[1]), 
    .enb(fbctrlb[1]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res FBRES_C_0 ( .out(out_cb), .ena(fbctrl[0]), 
    .enb(fbctrlb[0]), .in(in_c), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath_caps ACCAPS ( .out_t(in_t), .out_c(in_c), 
    .in_t(dqs_in_t), .in_c(dqs_in_c));

wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT PU0 ( .vdd(vdda), .en(ena), .y(out_tb));

wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT PD ( .vss(vss), .enb(enb), .y(out_cb));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf I64_4 ( .en(cal_cn), .out(out_cb), 
    .enb(cal_cp), .vss(vss), .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf I64_3 ( .en(cal_cn), .out(out_cb), 
    .enb(cal_cp), .vss(vss), .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf I64_2 ( .en(cal_cn), .out(out_cb), 
    .enb(cal_cp), .vss(vss), .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf I64_1 ( .en(cal_cn), .out(out_cb), 
    .enb(cal_cp), .vss(vss), .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf I64_0 ( .en(cal_cn), .out(out_cb), 
    .enb(cal_cp), .vss(vss), .in(in_c), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf INBUF_T_4 ( .en(cal_tn), .out(out_tb), 
    .enb(cal_tp), .vss(vss), .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf INBUF_T_3 ( .en(cal_tn), .out(out_tb), 
    .enb(cal_tp), .vss(vss), .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf INBUF_T_2 ( .en(cal_tn), .out(out_tb), 
    .enb(cal_tp), .vss(vss), .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf INBUF_T_1 ( .en(cal_tn), .out(out_tb), 
    .enb(cal_tp), .vss(vss), .in(in_t), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf INBUF_T_0 ( .en(cal_tn), .out(out_tb), 
    .enb(cal_tp), .vss(vss), .in(in_t), .vdd(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_core_v2,
//View - schematic
// LAST TIME SAVED: Dec 11 14:04:51 2020
// NETLIST TIME: Dec 12 00:59:11 2020
`timescale 1ps / 1ps 




 

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_core_v2 (dqs_out_c, dqs_out_t, vdda, vddq, 
    vss, cal_c_n, cal_c_p, cal_t_n, cal_t_p, dcpath_ena, dly_ctrl_c, 
    dly_ctrl_t, dqs_in_c, dqs_in_t, edge_det_byp, edge_det_ena, 
    edge_det_refsel, ena, fb_ena, rxcal_ena, se_mode);

output  dqs_out_c, dqs_out_t;

inout  vdda, vddq, vss;

input  dcpath_ena, dqs_in_c, dqs_in_t, edge_det_byp, edge_det_ena, 
    edge_det_refsel, ena, rxcal_ena, se_mode;

input [2:0]  fb_ena;
input [3:0]  cal_t_p;
input [3:0]  cal_t_n;
input [7:0]  dly_ctrl_t;
input [3:0]  cal_c_n;
input [7:0]  dly_ctrl_c;
input [3:0]  cal_c_p;

// Buses in the design

wire  [2:0]  fbNen;

wire  [3:0]  cal_tp;

wire  [3:0]  cal_tn;

wire  [3:0]  cal_cn;

wire  [3:0]  net095;

wire  [3:0]  cal_cp;

wire  [3:0]  net092;

wire  [2:0]  fbNen_b;


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath LOWSPEED_PATH ( .out_cb(acdc_nb), 
    .out_tb(acdc_tb), .in_t(dqs_in_t), .ena(dcena), .enb(dcenb), 
    .in_c(dqs_in_c), .se_ena(se_ena), .se_enb(se_enb), .vddq(vddq), 
    .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det SI ( .byp(edge_det_byp), .edge_det(frx_ena_dly), 
    .edge_det_b(frx_enb_dly), .in(dqs_in_c), .refsel(edge_det_refsel), 
    .ena(edge_det_ena), .vddq(vddq), .vdda(vdda), .vss(vss));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND12 ( .tielo(vss), .vdd(vdda), .y(dcenb), 
    .vss(vss), .tiehi(vdda), .b(ena_buf), .a(dcpath));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND9_3 ( .tielo(vss), .vdd(vdda), .y(cal_tp[3]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_p[3]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND9_2 ( .tielo(vss), .vdd(vdda), .y(cal_tp[2]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_p[2]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND9_1 ( .tielo(vss), .vdd(vdda), .y(cal_tp[1]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_p[1]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND9_0 ( .tielo(vss), .vdd(vdda), .y(cal_tp[0]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_p[0]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND0_2 ( .tielo(vss), .vdd(vdda), .y(fbNen_b[2]), 
    .vss(vss), .tiehi(vdda), .b(dcpath_b), .a(fb_ena[2]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND0_1 ( .tielo(vss), .vdd(vdda), .y(fbNen_b[1]), 
    .vss(vss), .tiehi(vdda), .b(dcpath_b), .a(fb_ena[1]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND0_0 ( .tielo(vss), .vdd(vdda), .y(fbNen_b[0]), 
    .vss(vss), .tiehi(vdda), .b(dcpath_b), .a(fb_ena[0]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND6_3 ( .tielo(vss), .vdd(vdda), .y(net092[3]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_n[3]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND6_2 ( .tielo(vss), .vdd(vdda), .y(net092[2]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_n[2]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND6_1 ( .tielo(vss), .vdd(vdda), .y(net092[1]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_n[1]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND6_0 ( .tielo(vss), .vdd(vdda), .y(net092[0]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_t_n[0]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND4 ( .tielo(vss), .vdd(vdda), .y(frx_enb), 
    .vss(vss), .tiehi(vdda), .b(ena_buf), .a(dcpath_b));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND7_3 ( .tielo(vss), .vdd(vdda), .y(net095[3]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_n[3]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND7_2 ( .tielo(vss), .vdd(vdda), .y(net095[2]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_n[2]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND7_1 ( .tielo(vss), .vdd(vdda), .y(net095[1]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_n[1]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND7_0 ( .tielo(vss), .vdd(vdda), .y(net095[0]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_n[0]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND8_3 ( .tielo(vss), .vdd(vdda), .y(cal_cp[3]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_p[3]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND8_2 ( .tielo(vss), .vdd(vdda), .y(cal_cp[2]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_p[2]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND8_1 ( .tielo(vss), .vdd(vdda), .y(cal_cp[1]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_p[1]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND8_0 ( .tielo(vss), .vdd(vdda), .y(cal_cp[0]), 
    .vss(vss), .tiehi(vdda), .b(frx_ena), .a(cal_c_p[0]));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND3 ( .tielo(vss), .vdd(vdda), .y(fp_enb_c), 
    .vss(vss), .tiehi(vdda), .b(net058), .a(net059));

wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT NAND2 ( .tielo(vss), .vdd(vdda), .y(fp_enb_t), 
    .vss(vss), .tiehi(vdda), .b(net051), .a(net052));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_course_delay COURSE_DELAY ( .fp_ena_c(fp_ena_c), 
    .fp_ena_t(fp_ena_t), .fp_enb_c(fp_enb_c), .fp_enb_t(fp_enb_t), 
    .in_cb(fine_c), .in_tb(fine_t), .out_c(dqs_out_c), 
    .out_t(dqs_out_t), .dly_ctrl_c(dly_ctrl_c[7:4]), 
    .dly_ctrl_t(dly_ctrl_t[7:4]), .vss(vss), .vdda(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV32_3 ( .in(net095[3]), .vss(vss), .out(cal_cn[3]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV32_2 ( .in(net095[2]), .vss(vss), .out(cal_cn[2]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV32_1 ( .in(net095[1]), .vss(vss), .out(cal_cn[1]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV32_0 ( .in(net095[0]), .vss(vss), .out(cal_cn[0]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV45 ( .in(dcenb), .vss(vss), .out(dcena), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV35 ( .in(cal_enb), .vss(vss), .out(cal_ena), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV31 ( .in(fp_enb_t), .vss(vss), .out(fp_ena_t), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV28 ( .in(enb), .vss(vss), .out(ena_buf), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV27 ( .in(dcpath_b), .vss(vss), .out(dcpath), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV26 ( .in(se_enb), .vss(vss), .out(se_ena), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV25 ( .in(se_mode), .vss(vss), .out(se_enb), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV29 ( .in(frx_enb), .vss(vss), .out(frx_ena), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV9_2 ( .in(fbNen_b[2]), .vss(vss), .out(fbNen[2]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV9_1 ( .in(fbNen_b[1]), .vss(vss), .out(fbNen[1]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV9_0 ( .in(fbNen_b[0]), .vss(vss), .out(fbNen[0]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV34 ( .in(rxcal_ena), .vss(vss), .out(cal_enb), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV30_3 ( .in(net092[3]), .vss(vss), .out(cal_tn[3]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV30_2 ( .in(net092[2]), .vss(vss), .out(cal_tn[2]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV30_1 ( .in(net092[1]), .vss(vss), .out(cal_tn[1]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV30_0 ( .in(net092[0]), .vss(vss), .out(cal_tn[0]), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV13 ( .in(dcpath_ena), .vss(vss), .out(dcpath_b), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV8 ( .in(ena), .vss(vss), .out(enb), .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT INV24 ( .in(fp_enb_c), .vss(vss), .out(fp_ena_c), 
    .vdd(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT NOR0 ( .tielo(vss), .tiehi(vdda), .y(net051), 
    .vss(vss), .vdd(vdda), .b(dly_ctrl_t[4]), .a(dly_ctrl_t[5]));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT NOR001 ( .tielo(vss), .tiehi(vdda), .y(net052), 
    .vss(vss), .vdd(vdda), .b(dly_ctrl_t[6]), .a(dly_ctrl_t[7]));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT NOR2 ( .tielo(vss), .tiehi(vdda), .y(net059), 
    .vss(vss), .vdd(vdda), .b(dly_ctrl_c[6]), .a(dly_ctrl_c[7]));

wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT NOR3 ( .tielo(vss), .tiehi(vdda), .y(net058), 
    .vss(vss), .vdd(vdda), .b(dly_ctrl_c[4]), .a(dly_ctrl_c[5]));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay FINE_DELAY ( .out_c(fine_c), 
    .out_t(fine_t), .cal_ena(cal_ena), .cal_enb(cal_enb), 
    .dly_ctrl_c(dly_ctrl_c[3:0]), .dly_ctrl_t(dly_ctrl_t[3:0]), 
    .ena(frx_ena_dly), .enb(frx_enb_dly), .in_c(acdc_nb), 
    .in_t(acdc_tb), .vss(vss), .vdda(vdda));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath HIGHSPEED_PATH ( .fbctrlb(fbNen_b[2:0]), 
    .fbctrl(fbNen[2:0]), .out_cb(acdc_nb), .out_tb(acdc_tb), 
    .cal_cn(cal_cn[3:0]), .cal_cp(cal_cp[3:0]), .cal_tn(cal_tn[3:0]), 
    .cal_tp(cal_tp[3:0]), .dqs_in_c(dqs_in_c), .dqs_in_t(dqs_in_t), 
    .ena(ena_buf), .enb(enb), .vss(vss), .vdda(vdda));

endmodule
// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_dqs_rcvr_no_esd,
//View - schematic
// LAST TIME SAVED: Dec 11 10:22:08 2020
// NETLIST TIME: Dec 12 00:59:11 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_dqs_rcvr_no_esd (d_dqs_out_c, d_dqs_out_t,  
      d_cal_n_c, d_cal_n_t, d_cal_p_c, d_cal_p_t, 
    d_dcpath_ena, d_dly_ctrl_c, d_dly_ctrl_t, d_edge_det_byp, 
    d_edge_det_ena, d_edge_det_refsel, d_ena, d_fb_ena, d_rxcal_ena, 
    d_se_mode, dqs_in_c, dqs_in_t
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vddq  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vddq;
assign vddq=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vddq;
inout vss;
`endif


output  d_dqs_out_c, d_dqs_out_t;



input  d_dcpath_ena, d_edge_det_byp, d_edge_det_ena, d_edge_det_refsel, 
    d_ena, d_rxcal_ena, d_se_mode, dqs_in_c, dqs_in_t;

input [3:0]  d_cal_p_c;
input [7:0]  d_dly_ctrl_t;
input [3:0]  d_cal_n_t;
input [7:0]  d_dly_ctrl_c;
input [3:0]  d_cal_n_c;
input [3:0]  d_cal_p_t;
input [2:0]  d_fb_ena;

`ifdef SYNTHESIS
`else 

logic dqs_in_t_channel;
logic dqs_in_c_channel;

wphy_lp4x5_dqs_rcvr_no_esd_wphy_real_channel_model #(
     //parameters
     .COEFF_FILE         ( "channel_coeffs_10ps.txt"),
     .TIMESTEP_PS        ( 7        ),
     .NUM_OF_COEFFS      ( 20        ),
     .DELAY              ( 0        ),         // in ps
     .AMP_RATIO          ( 1        )         // 0<=value<=1,
   ) CH_T (
     .rx_in(dqs_in_t),
     .rxp_out(dqs_in_t_channel));

wphy_lp4x5_dqs_rcvr_no_esd_wphy_real_channel_model #(
     //parameters
     .COEFF_FILE         ( "channel_coeffs_10ps.txt"),
     .TIMESTEP_PS        ( 7        ),
     .NUM_OF_COEFFS      ( 20        ),
     .DELAY              ( 0        ),         // in ps
     .AMP_RATIO          ( 1        )         // 0<=value<=1,
   ) CH_C (
     .rx_in(dqs_in_c),
     .rxp_out(dqs_in_c_channel));


wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_core_v2 DQS_RCVR ( .edge_det_byp(d_edge_det_byp), 
    .edge_det_ena(d_edge_det_ena), .edge_det_refsel(d_edge_det_refsel), 
    .dqs_in_t(dqs_in_t_channel), .rxcal_ena(d_rxcal_ena), 
    .cal_c_n(d_cal_n_c[3:0]), .cal_c_p(d_cal_p_c[3:0]), 
    .cal_t_n(d_cal_n_t[3:0]), .fb_ena(d_fb_ena[2:0]), .vddq(vddq), 
    .cal_t_p(d_cal_p_t[3:0]), .dqs_out_c(d_dqs_out_c), 
    .dqs_out_t(d_dqs_out_t), .vss(vss), .vdda(vdda), 
    .dqs_in_c(dqs_in_c_channel), .se_mode(d_se_mode), 
    .dly_ctrl_c(d_dly_ctrl_c[7:0]), .dly_ctrl_t(d_dly_ctrl_t[7:0]), 
    .ena(d_ena), .dcpath_ena(d_dcpath_ena));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell -
//wphy_lp4x5_dqs_rcvr_no_esd_tb, View - schematic
// LAST TIME SAVED: Dec 11 22:01:46 2020
// NETLIST TIME: Dec 12 00:59:12 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_inbuf ( in, vdd, vss, out, en, enb );

  input in;
  output out;
  input  [3:0] en;
  inout vdd;
  input  [3:0] enb;
  inout vss;

  assign out = (|en) ? ~in : 1'bz;

endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath_caps"
//"systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_acpath_caps ( out_c, out_t, in_c, in_t );

  input in_t;
  output reg out_t;
  input in_c;
  output reg out_c;

  real ac_delay = 35.0;

  initial begin
    out_c = in_c;
    out_t = in_t;
  end

  always @(*) begin
    out_c <= #(ac_delay) in_c;
  end

  always @(*) begin
    out_t <= #(ac_delay) in_t;
  end

endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res"
//"systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_fb_mos_res ( in, out, vdda, vss, ena, enb );

  inout in;
  inout vdda;
  inout out;
  input ena;
  input enb;
  inout vss;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT_Mmod_delay"
//"systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT_Mmod_nomodel( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
  input en;
  input enb;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG


endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay_capdac"
//"systemVerilog"

`timescale 1ps/1fs

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_fine_delay_capdac ( out, vss, dly_ctrl, in );

  input in;
  output out;
  input  [3:0] dly_ctrl;
  inout vss;

  reg out_reg;

  wire power_ok;
  assign power_ok = ~vss;
  real fine_delay = 0.85;
  real total_fine_delay;

  initial begin
    total_fine_delay=dly_ctrl*fine_delay;
    out_reg <= #(total_fine_delay) in;
  end

  always @(*) begin
    total_fine_delay=dly_ctrl*fine_delay;
    out_reg <= #(total_fine_delay) in;
  end
 
  assign out = (power_ok) ? out_reg : 1'bx; 

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_course_delay"
//"systemVerilog"

`timescale 1ps/1fs

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_course_delay ( out_c, out_t, vdda, vss, dly_ctrl_c,
dly_ctrl_t, fp_ena_c, fp_ena_t, fp_enb_c, fp_enb_t, in_cb, in_tb );

  input  [3:0] dly_ctrl_t;
  input in_cb;
  input fp_enb_t;
  input in_tb;
  inout vdda;
  output out_t;
  output out_c;
  input  [3:0] dly_ctrl_c;
  input fp_enb_c;
  input fp_ena_t;
  input fp_ena_c;
  inout vss;


  reg out_t_reg;
  reg out_c_reg;

  wire power_ok;
  assign power_ok = ~vss & vdda;
  real coarse_t_delay = 13.6;
  real coarse_c_delay = 13.6;
  real total_coarse_t_delay;
  real total_coarse_c_delay;

  initial begin
    total_coarse_t_delay=dly_ctrl_t*coarse_t_delay;
    out_t_reg <= #(total_coarse_t_delay) ~in_tb;

    total_coarse_c_delay=dly_ctrl_c*coarse_c_delay;
    out_c_reg <= #(total_coarse_c_delay) ~in_cb;
  end

  always @(*) begin
    total_coarse_t_delay=dly_ctrl_t*coarse_t_delay;
    out_t_reg <= #(total_coarse_t_delay) ~in_tb;
  end

  always @(*) begin
    total_coarse_c_delay=dly_ctrl_c*coarse_c_delay;
    out_c_reg <= #(total_coarse_c_delay) ~in_cb;
  end
 
  assign out_t = (power_ok) ? out_t_reg : 1'bx;
  assign out_c = (power_ok) ? out_c_reg : 1'bx;



endmodule



module wphy_lp4x5_dqs_rcvr_no_esd_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT_timing( in, out
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign out = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign (weak1,weak0) #(3) out =  ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_timing( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

    assign (weak1,weak0) #(3)  out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_LVT" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_NOR2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);


endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det_sf" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_hc_tst_dqs_edge_det_sf ( out, vdda, vddq, vss, ena, in, refsel );

  input refsel;
  input in;
  inout vdda;
  output out;
  input ena;
  inout vddq;
  inout vss;


wire power_ok;
assign power_ok = vdda & vddq & (~vss);

assign out = ena & in;

endmodule
//systemVerilog HDL for "wphy_gf12lp_lp4x5_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath_lvlshift"
//"systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rx_dcpath_lvlshift ( out_cb, out_tb, vdda, vss, in_c,
in_t );

  input in_t;
  inout vdda;
  output out_tb;
  input in_c;
  output out_cb;
  inout vss;

  reg out_tb_reg;
  reg out_cb_reg;

  real dc_path_delay=225.0;

  wire power_ok;
  assign power_ok = vdda & (~vss);

  initial begin
    out_tb_reg =  ~in_t;
    out_cb_reg =  ~in_c;
  end

  always @(*) begin
    out_tb_reg <= #(dc_path_delay)  ~in_t;
  end

  always @(*) begin
    out_cb_reg <= #(dc_path_delay)  ~in_c;
  end

  assign out_tb = (power_ok) ? out_tb_reg : 1'bx;
  assign out_cb = (power_ok) ? out_cb_reg : 1'bx;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D1_GL16_LVT( in, out
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign out = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

    assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT" "systemVerilog"

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_INVT( in, out, en, enb 
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG



assign out = (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT" "systemVerilog"

module wphy_lp4x5_dqs_rcvr_no_esd_INVT_D2_GL16_LVT( in, out, en, enb 
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG



assign out = (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT" "systemVerilog"

`timescale 1ps/1ps

module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

    assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_PU_D2_GL16_LVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign  y = en ? 1'bz : 1'b1;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT" "systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_PD_D2_GL16_LVT ( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel"
//"systemVerilog"


module wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_wphy_lp4x5_dqs_rcvr_no_esd_INV_D2_GL16_LVT_Mmod_nomodel( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG


endmodule

`timescale 1ps/1ps
module wphy_lp4x5_dqs_rcvr_no_esd_wphy_real_channel_model #(
  parameter     NUM_OF_COEFFS   = 200,
  parameter     TIMESTEP_PS     = 10,
  parameter     COEFF_FILE      = "channel_coeffs_10ps.txt",
  parameter     DELAY           = 0,
  parameter     AMP_RATIO       = 1
)(  rx_in, rxp_out);
 
input   rx_in;
output  rxp_out;

`ifdef WCHANNEL_EN
reg rxp_out_reg;
integer skew=0;
integer max_c2c_jit=0;
integer max_accum_jit=0;

initial begin
   rxp_out_reg = rx_in;
end

initial begin
    if ($value$plusargs("RCVR_SKEW=%d", skew)) begin
    end
    if ($value$plusargs("RCVR_MAX_C2C_JIT=%d", max_c2c_jit)) begin
    end
    if ($value$plusargs("RCVR_MAX_ACCUM_JIT=%d", max_accum_jit)) begin
    end

end


always @(rx_in) begin
  rxp_out_reg <= #(30) rx_in;  //the delay matches SA channel model delay
end

//assign rxp_out = rxp_out_reg;

ddr_jitter_buf u_jitter_buf (
   .i_clk(rxp_out_reg),
   .i_skew(skew),
   .i_max_c2c_jit(max_c2c_jit),
   .i_max_accum_jit(max_accum_jit),
   .o_clk(rxp_out)
);
`else

assign rxp_out = rx_in;

`endif


endmodule

`endif //SYNTHESIS
