module libmodule;
endmodule
