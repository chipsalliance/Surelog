/*
:name: empty_test_5
:description: Test
:type: preprocessing
:tags: 5.3 5.4
*/
/* comment */
