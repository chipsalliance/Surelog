/*
:name: typedef_test_24
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef struct {
  int sample;
  int tile;
} tuple_t;