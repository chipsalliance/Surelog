/*
:name: 22.11--pragma-invalid
:description: Test
:should_fail_because: pragma macro takes name as an argument
:tags: 22.11
:type: preprocessing
*/
`pragma
