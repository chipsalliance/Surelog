
 //pragma translate_off

class a;

endclass

 //pragma translate_on

module top ();

assign a = b;

//pragma translate_off

  ggggll
  
//pragma translate_on

assign c = d;


endmodule
