/*
:name: string_atobin
:description: string.atobin()  tests
:tags: 6.16.9
*/
module top();
	string a = "10101";
	int b = a.atobin();
endmodule
