/*
:name: class_test_42
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class macros_as_class_item;
 `uvm_object_utils_begin(foobar)
 `uvm_object_utils(blah)
 `uvm_object_utils_end
endclass