/*
:name: specparam
:description: specparam tests
:should_fail: 0
:tags: 6.20.5
*/
module top();
	specparam delay = 50;
endmodule
