/*
:name: 22.11--pragma-number-multi
:description: Test
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_number_other a = 123, b = 4
