module dut;

   function [1:0] foo;
   
   endfunction

   function bar;
   
   endfunction

endmodule

