/*
:name: class_test_59
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
`ifdef DEBUGGER
`endif
endclass