module top ();
   middleman #(.invert(1)) mdl1();
   middleman #(.invert(0)) mdl0();
endmodule


