/*
:name: global_constant
:description: class with global constant variable
:should_fail: 0
:tags: 8.19
*/
module class_tb ();
	class a_cls;
		const int c = 12;
	endclass
endmodule
