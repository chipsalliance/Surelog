/*
:name: string_len
:description: string.len()  tests
:should_fail: 0
:tags: 6.16.1
*/
module top();
	string a = "Test";
	int b = a.len();
endmodule
