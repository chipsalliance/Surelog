/*
:name: attributes-module
:description: Assing attributes to a module
:should_fail: 0
:tags: 5.12
*/

(* optimize_power *)
module topa();
endmodule

(* optimize_power=0 *)
module topb();
endmodule

(* optimize_power=1 *)
module topc();
endmodule
