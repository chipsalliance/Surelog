// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: number_test_3
:description: Test
:tags: 5.6.4 5.7.1 5.7.2
*/
parameter int foo = '1;

module test;
endmodule
