/*
:name: class_member_test_19
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subr(bool x[N]);
endclass