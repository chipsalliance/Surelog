/*
:name: iface_class_test_3
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic extends basebase;
endclass