/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

uvm_resource_db#(bit)::set(.scope("REG::*WDDR_CMN_PLL_CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1"), .name("NO_REG_TESTS"), .val(1), .accessor(this));
uvm_resource_db#(bit)::set(.scope("REG::*WDDR_CMN_PLL_CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1"), .name("NO_REG_TESTS"), .val(1), .accessor(this));
uvm_resource_db#(bit)::set(.scope("REG::*WDDR_CMN_PLL_CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1"), .name("NO_REG_TESTS"), .val(1), .accessor(this));
uvm_resource_db#(bit)::set(.scope("REG::*WDDR_INTF_INTF_MODE"), .name("NO_REG_TESTS"), .val(1), .accessor(this));
uvm_resource_db#(bit)::set(.scope("REG::*WDDR_CTRL_CTRL_CLK_CFG"), .name("NO_REG_TESTS"), .val(1), .accessor(this));

uvm_resource_db#(bit)::set(.scope("REG::*_CFG_7"), .name("NO_REG_TESTS"), .val(1), .accessor(this));
