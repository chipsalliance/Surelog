// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: struct_test_0
:description: Test
:tags: 7.2
*/
typedef struct mystruct_fwd;

typedef struct { logic a; logic b; } mystruct_fwd;

module test;
endmodule
