/*
:name: preproc_test_1
:description: Test
:should_fail: 0
:tags: 5.6.4
*/
`define FOO BAR-1
