module top(b);
input b;
reg N=0.0/0'H0;
endmodule

