/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s001
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 15762
// Design library name: wphy_gf12lp_lp4x5_sim_lib
// Design cell name: wphy_lp4x5_cke_drvr_w_lpbk_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_lp4x5_lib, Cell - wphy_lp4x5_cke_drvr_w_lpbk,
//View - schematic
// LAST TIME SAVED: Sep 22 07:33:55 2020
// NETLIST TIME: Oct 29 04:02:09 2020
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_lp4x5_cke_drvr_w_lpbk (d_lpbk_out, pad_cke_out,  
      d_bs_din, d_bs_ena, d_in_c, d_lpbk_ena, d_ovrd, 
    d_ovrd_val, freeze_n_hv
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vdda1p2  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vdda1p2;
assign vdda1p2=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vdda1p2;
inout vss;
`endif


output  d_lpbk_out;

inout  pad_cke_out;

input  d_bs_din, d_bs_ena, d_in_c, d_lpbk_ena, d_ovrd_val, freeze_n_hv;

input [2:0]  d_ovrd;

`ifdef SYNTHESIS
`else 

wphy_lp4x5_cke_drvr_w_lpbk_MUXT2_D2_GL16_RVT MUX1 ( .vss(vss), .sb(bs_enb), .s(bs_ena), 
    .b(d_bs_din), .a(d_ovrd_val), .yb(ovrd_b_input), .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_MUXT2_D2_GL16_RVT MUX0 ( .vss(vss), .sb(ovrdORbs), .s(ovrdNORbs), 
    .b(d_in_c), .a(ovrd_b_input), .yb(in_t), .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT INV3 ( .in(ovrdNORbs), .vss(vss), .out(ovrdORbs), 
    .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT INV6 ( .in(d_bs_ena), .vss(vss), .out(bs_enb), 
    .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT INV7 ( .in(bs_enb), .vss(vss), .out(bs_ena), 
    .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT INV0 ( .in(ovrd_b), .vss(vss), .out(ovrd), .vdd(vdda));

wphy_lp4x5_cke_drvr_w_lpbk_NOR2_D1_GL16_LVT NOR1 ( .tielo(vss), .tiehi(vdda), .y(ovrdNORbs), 
    .vss(vss), .vdd(vdda), .b(bs_ena), .a(ovrd));

wphy_lp4x5_cke_drvr_w_lpbk_wphy_lp4x5_cke_drv_core DRV ( .vdda1p2(vdda1p2), .out_h(pad_cke_out), 
    .inb_h(inb_h), .vss(vss));

wphy_lp4x5_cke_drvr_w_lpbk_INV_D1_GL150_EGU INV2 ( .vdda1p2(vdda), .in(net014), .vss(vss), 
    .out(d_lpbk_out));

wphy_lp4x5_cke_drvr_w_lpbk_LVLHC0_D1_GL16_RVT LVLSFT0 ( .freezeb_hv(freeze_n_hv), 
    .outn(lpbk_enb_h), .in(d_lpbk_ena), .outp(lpbk_ena_h), 
    .vdda1p8(vdda1p2), .vdd(vdda), .vss(vss));

wphy_lp4x5_cke_drvr_w_lpbk_LVLHC0_D1_GL16_RVT LS0 ( .freezeb_hv(freeze_n_hv), .outn(inb_h), 
    .in(in_t), .outp(net015), .vdda1p8(vdda1p2), .vdd(vdda), 
    .vss(vss));

wphy_lp4x5_cke_drvr_w_lpbk_NOR3_D1_GL16_RVT NOR0 ( .vdd(vdda), .c(d_ovrd[0]), .y(ovrd_b), 
    .vss(vss), .b(d_ovrd[1]), .a(d_ovrd[2]));

wphy_lp4x5_cke_drvr_w_lpbk_wphy_esd_prim_diodes PRIM_ESD0 ( .vss(vss), .vddq(vdda1p2), 
    .pad(pad_cke_out));

wphy_lp4x5_cke_drvr_w_lpbk_wphy_esd_sec_diodes SEC_ESD1 ( .vdd(vdda1p2), .vss(vss), .out(rxin_h), 
    .in(pad_cke_out));

wphy_lp4x5_cke_drvr_w_lpbk_NAND2_D1_GL150_EGU NAND0 ( .y(net014), .vss(vss), .vdda1p2(vdda1p2), 
    .b(lpbk_ena_h), .a(rxin_h));

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_lp4x5_sim_lib, Cell -
//wphy_lp4x5_cke_drvr_w_lpbk_tb, View - schematic
// LAST TIME SAVED: Oct 29 03:29:57 2020
// NETLIST TIME: Oct 29 04:02:09 2020
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "NAND2_D1_GL150_UD12" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_NAND2_D1_GL150_EGU ( y, a, b
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdda1p2 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p2;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdda1p2;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y = ~(a&b);


endmodule

module wphy_lp4x5_cke_drvr_w_lpbk_wphy_esd_sec_diodes( out, in, vdd, vss );

  input reg in;
  inout vdd;
`ifdef WPIN_EN
  output integer out;
`else
  output reg out;
`endif
  inout vss;

initial begin
  if (in === 1'bx) begin
    out = 1'bx;
  end else if (in === 1'bz) begin
    out = 1'bz;
  end else if (in == 1'b1) begin
`ifdef WPIN_EN
    out = 1000;
`else
    out = 1;
`endif
  end else if (in == 1'b0) begin
    out = 0;
  end
end

always @(*) begin
  if (in === 1'bx) begin
    out = 1'bx;
  end else if (in === 1'bz) begin
    out = 1'bz;
  end else if (in == 1'b1) begin
`ifdef WPIN_EN
    out = 1000;
`else
    out = 1;
`endif
  end else if (in == 1'b0) begin
    out = 0;
  end 
end

endmodule
//Verilog HDL for "aic_shared", "esd_prim_diodes" "functional"


module wphy_lp4x5_cke_drvr_w_lpbk_wphy_esd_prim_diodes( pad, vddq, vss );

  inout pad;
  inout vddq;
  inout vss;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cke_drvr_w_lpbk_NOR3_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_NOR3_D1_GL16_RVT ( y, a, b, c
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input c;
  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y = ~(a|b|c);



endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cke_drvr_w_lpbk_LVLHC0_D1_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_LVLHC0_D1_GL16_RVT ( outn, outp, in, freezeb_hv
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd, vdda1p8 
`endif //WLOGIC_MODEL_NO_PG
); 

  input freezeb_hv;
  input in;
  output outn;
  output outp;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p8;
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
  assign outp = ~freezeb_hv ? 1'b0 : in;
  assign outn = ~freezeb_hv ? 1'b1 : ~in;
`else

  assign outp = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b0 : in)  : 1'b0;
  assign outn = (vdd & vdda1p8 & ~vss) ? (~freezeb_hv ? 1'b1 : ~in) : 1'b0;

`endif //WLOGIC_MODEL_NO_PG



endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "INV_D1_GL150_UD12" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_INV_D1_GL150_EGU ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdda1p2, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdda1p2;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdda1p2;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//Verilog HDL for "wphy_lp4x5_lib", "wphy_lp4x5_cke_drvr_w_lpbk_wphy_lp4x5_cke_drv_core" "functional"


module wphy_lp4x5_cke_drvr_w_lpbk_wphy_lp4x5_cke_drv_core ( out_h, vdda1p2, vss, inb_h );

  output out_h;
  inout vdda1p2;
  input inb_h;
  inout vss;

	wire pwr_ok;
	assign pwr_ok = vdda1p2 & ~vss;
	assign out_h = pwr_ok ? ~inb_h : 1'bx;
endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cke_drvr_w_lpbk_NOR2_D1_GL16_LVT" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_NOR2_D1_GL16_LVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


  assign y=~(a|b);


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_lp4x5_cke_drvr_w_lpbk_MUXT2_D2_GL16_RVT" "systemVerilog"


module wphy_lp4x5_cke_drvr_w_lpbk_MUXT2_D2_GL16_RVT( yb, a, b, s, sb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input a; 
  input sb;
  input s;
  output yb;
  input b;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire yb;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign yb = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign yb = (s && ~sb) ? ~b:~a;



endmodule
`endif //SYNTHESIS
