package my_pkg;
   function automatic void assign_1();
   endfunction 
   function automatic logic assign_2();
   endfunction 
   function automatic assign_3();
   endfunction 

endpackage 
