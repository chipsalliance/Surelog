
`ifndef BP_FE_ICACHE_VH
`define BP_FE_ICACHE_VH

`include "bp_common_me_if.vh"

`endif
