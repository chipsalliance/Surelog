module top();
  always @(posedge clock) begin

     if (_GEN_4174 & _T_3461) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:1321 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%x, expected %%x\", hartExceptionId, 0.U)\n"); // @[Debug.scala 1321:15:boom.system.TestHarness.SmallBoomConfig.fir@94896.14]
        end
     end

































































































































































































































































































































































































class toto;
endclass































                
















































































































 always @(posedge clock) begin

     if (_GEN_4174 & _T_3461) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected 'EXCEPTION' hart\n    at Debug.scala:1321 assert(hartExceptionId === 0.U, \"Unexpected 'EXCEPTION' hart\")//Chisel3 #540, %%x, expected %%x\", hartExceptionId, 0.U)\n"); // @[Debug.scala 1321:15:boom.system.TestHarness.SmallBoomConfig.fir@94896.14]
        end
     end


endmodule