/*
:name: desc_test_1
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
`ifdef VERBOSE
`else
`endif
`endif
