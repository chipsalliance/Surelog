/*
:name: 22.11--pragma-basic
:description: Test
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_name "pragma_value"
