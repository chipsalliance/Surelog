/*
:name: parameter_type
:description: parameter type tests
:tags: 6.20.3
*/
module top #(type T = real);
endmodule
