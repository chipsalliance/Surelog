/*
:name: 22.7--timescale-basic-3
:description: Test
:should_fail_because: the valid integers in this type of expression are 1, 10, and 100
:tags: 22.7
:type: simulation
*/
`timescale 9 ns / 1 ps
