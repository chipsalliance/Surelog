/*
:name: event
:description: event type tests
:tags: 6.17
*/
module top();
	event a;
endmodule
