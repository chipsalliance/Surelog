/*
:name: queues-basic
:description: Test queues support
:tags: 7.10
*/
module top ();

int q[$];

endmodule
