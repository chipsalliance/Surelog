// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: iface_class_test_10
:description: Test
:tags: 8.3 8.26
*/
interface class base_ic;
pure virtual function void pure_task1;
pure virtual function string concatenator(string arg);
endclass

module test;
endmodule
