module wire_top(inp, xn);
    input wire signed inp;
    output reg [4:0] xn;

    assign xn = inp;
endmodule
