// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: enum_anon
:description: anonymous enum tests
:tags: 6.19
*/
module top();
	enum {a, b, c} val;
endmodule
