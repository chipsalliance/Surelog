// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: cast_op
:description: cast operator
:tags: 6.24.1
*/
module top();
	int a = int'(2.1 * 3.7);
endmodule
