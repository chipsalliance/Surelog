/*
:name: cast_op
:description: cast operator
:tags: 6.24.1
*/
module top();
	int a = int'(2.1 * 3.7);
endmodule
