
module top();

   for (i = 3; i > 0 ; i--) begin
      assign tmp[i] = 1'b1;
   end

endmodule