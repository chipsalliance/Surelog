/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/
`include "APB/APB_agent/wav_APB_vif.sv"
`include "APB/APB_agent/wav_APB_Agent_config.sv"
`include "APB/APB_agent/wav_APB_transfer.sv"
`include "APB/APB_agent/wav_APB_monitor.sv"
`include "APB/APB_agent/wav_APB_sequencer.sv"
`include "APB/APB_agent/wav_APB_driver.sv"
`include "APB/APB_agent/wav_APB_agent.sv"
`include "APB/APB_agent/wav_APB_seq_lib.sv"
`include "APB/APB_agent/reg_to_apb_adapter.sv"
