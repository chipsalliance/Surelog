/*
:name: net_decl_assignment
:description: net declaration assignment test
:should_fail: 0
:tags: 10.3.1
*/
module top(input a, input b);

wire w = a & b;

endmodule
