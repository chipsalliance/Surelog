module top(b);inout b;reg c;assign+0-c=b;endmodule

