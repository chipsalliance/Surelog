/*
:name: class_member_test_39
:description: Test
:should_fail: 0
:tags: 8.3
*/
class constructible;
function new;
endfunction
endclass