module top;
   byte b[] = {1, 1, 1};
  
endmodule
