/*
:name: associative-arrays-class
:description: Test associative arrays support
:should_fail: 0
:tags: 7.8.3 7.8
*/
module top ();

class C;
    int x;
endclass

int arr [ C ];

endmodule
