// This file exists for preproc_test_2.sv
`define SUCCESS
