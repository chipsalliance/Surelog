// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: min_max_avg_delay
:description: minimum, typical and maximum delay expressions test
:tags: 11.11
*/
module top();

initial begin
	#(100:200:300) $display("Done");
end

endmodule
