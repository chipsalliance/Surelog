/*
:name: class_member_test_18
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subroutine(input bool x);
endclass