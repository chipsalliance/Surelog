/*********************************************************************************
Copyright (c) 2021 Wavious LLC

This program is free software: you can redistribute it and/or modify
it under the terms of the GNU General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

This program is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU General Public License for more details.

You should have received a copy of the GNU General Public License
along with this program.  If not, see <http://www.gnu.org/licenses/>.

*********************************************************************************/

`define MCUTOP_SWI_RSVD                                                        'h00000000
`define MCUTOP_SWI_RSVD__RSVD                                                        31:0
`define MCUTOP_SWI_RSVD___POR                                                32'h00000000

`define MCUTOP_SWI_CFG                                                         'h00000004
`define MCUTOP_SWI_CFG__FETCH_EN                                                        0
`define MCUTOP_SWI_CFG__DEBUG_EN                                                        1
`define MCUTOP_SWI_CFG___POR                                                 32'h00000000

`define MCUTOP_SWI_STA                                                         'h00000008
`define MCUTOP_SWI_STA__RESERVED0                                                    31:0
`define MCUTOP_SWI_STA___POR                                                 32'h00000000

`define MCUINTF_SWI_HOST2MCU_MSG_DATA                                          'h00000000
`define MCUINTF_SWI_HOST2MCU_MSG_DATA__DATA                                          31:0
`define MCUINTF_SWI_HOST2MCU_MSG_DATA___POR                                  32'h00000000

`define MCUINTF_SWI_HOST2MCU_MSG_ID                                            'h00000004
`define MCUINTF_SWI_HOST2MCU_MSG_ID__ID                                              31:0
`define MCUINTF_SWI_HOST2MCU_MSG_ID___POR                                    32'h00000000

`define MCUINTF_SWI_HOST2MCU_MSG_REQ                                           'h00000008
`define MCUINTF_SWI_HOST2MCU_MSG_REQ__REQ                                               0
`define MCUINTF_SWI_HOST2MCU_MSG_REQ___POR                                   32'h00000000

`define MCUINTF_SWI_HOST2MCU_MSG_ACK                                           'h0000000C
`define MCUINTF_SWI_HOST2MCU_MSG_ACK__ACK                                               0
`define MCUINTF_SWI_HOST2MCU_MSG_ACK___POR                                   32'h00000000

`define MCUINTF_SWI_MCU2HOST_MSG_DATA                                          'h00000010
`define MCUINTF_SWI_MCU2HOST_MSG_DATA__DATA                                          31:0
`define MCUINTF_SWI_MCU2HOST_MSG_DATA___POR                                  32'h00000000

`define MCUINTF_SWI_MCU2HOST_MSG_ID                                            'h00000014
`define MCUINTF_SWI_MCU2HOST_MSG_ID__ID                                              31:0
`define MCUINTF_SWI_MCU2HOST_MSG_ID___POR                                    32'h00000000

`define MCUINTF_SWI_MCU2HOST_MSG_REQ                                           'h00000018
`define MCUINTF_SWI_MCU2HOST_MSG_REQ__REQ                                               0
`define MCUINTF_SWI_MCU2HOST_MSG_REQ___POR                                   32'h00000000

`define MCUINTF_SWI_MCU2HOST_MSG_ACK                                           'h0000001C
`define MCUINTF_SWI_MCU2HOST_MSG_ACK__ACK                                               0
`define MCUINTF_SWI_MCU2HOST_MSG_ACK___POR                                   32'h00000000

`define MCU_SWI_IRQ_FAST_CLR_CFG                                               'h00000000
`define MCU_SWI_IRQ_FAST_CLR_CFG__CLR                                                31:0
`define MCU_SWI_IRQ_FAST_CLR_CFG___POR                                       32'h00000000

`define MCU_SWI_IRQ_FAST_STICKY_CFG                                            'h00000004
`define MCU_SWI_IRQ_FAST_STICKY_CFG__EN                                              31:0
`define MCU_SWI_IRQ_FAST_STICKY_CFG___POR                                    32'h00000000

`define MCU_SWI_IRQ_FAST_MSK_CFG                                               'h00000008
`define MCU_SWI_IRQ_FAST_MSK_CFG__MSK                                                31:0
`define MCU_SWI_IRQ_FAST_MSK_CFG___POR                                       32'h00000000

`define MCU_SWI_IRQ_FAST_SYNC_CFG                                              'h0000000C
`define MCU_SWI_IRQ_FAST_SYNC_CFG__EN                                                31:0
`define MCU_SWI_IRQ_FAST_SYNC_CFG___POR                                      32'h00000000

`define MCU_SWI_IRQ_FAST_EDGE_CFG                                              'h00000010
`define MCU_SWI_IRQ_FAST_EDGE_CFG__EN                                                31:0
`define MCU_SWI_IRQ_FAST_EDGE_CFG___POR                                      32'h00000000

`define MCU_SWI_IRQ_FAST_STA                                                   'h00000014
`define MCU_SWI_IRQ_FAST_STA__IRQ_STA                                                31:0
`define MCU_SWI_IRQ_FAST_STA___POR                                           32'h00000000

`define MCU_SWI_MSIP_CFG                                                       'h00000018
`define MCU_SWI_MSIP_CFG__INTERRUPT                                                     0
`define MCU_SWI_MSIP_CFG___POR                                               32'h00000000

`define MCU_SWI_MTIME_LO_STA                                                   'h0000001C
`define MCU_SWI_MTIME_LO_STA__TIME_LO                                                31:0
`define MCU_SWI_MTIME_LO_STA___POR                                           32'h00000000

`define MCU_SWI_MTIME_HI_STA                                                   'h00000020
`define MCU_SWI_MTIME_HI_STA__TIME_HI                                                31:0
`define MCU_SWI_MTIME_HI_STA___POR                                           32'h00000000

`define MCU_SWI_MTIMECMP_LO_CFG                                                'h00000024
`define MCU_SWI_MTIMECMP_LO_CFG__TIMECMP_LO                                          31:0
`define MCU_SWI_MTIMECMP_LO_CFG___POR                                        32'h00000000

`define MCU_SWI_MTIMECMP_HI_CFG                                                'h00000028
`define MCU_SWI_MTIMECMP_HI_CFG__TIMECMP_HI                                          31:0
`define MCU_SWI_MTIMECMP_HI_CFG___POR                                        32'h00000000

`define MCU_SWI_MTIMECMP_CFG                                                   'h0000002C
`define MCU_SWI_MTIMECMP_CFG__LOAD                                                      0
`define MCU_SWI_MTIMECMP_CFG___POR                                           32'h00000000

`define MCU_SWI_MTIME_CFG                                                      'h00000030
`define MCU_SWI_MTIME_CFG__ENABLE                                                       0
`define MCU_SWI_MTIME_CFG___POR                                              32'h00000001

`define MCU_SWI_GP0_CFG                                                        'h00000034
`define MCU_SWI_GP0_CFG__RESERVED0                                                   31:0
`define MCU_SWI_GP0_CFG___POR                                                32'h00000000

`define MCU_SWI_GP1_CFG                                                        'h00000038
`define MCU_SWI_GP1_CFG__RESERVED0                                                   31:0
`define MCU_SWI_GP1_CFG___POR                                                32'h00000000

`define MCU_SWI_GP2_CFG                                                        'h0000003C
`define MCU_SWI_GP2_CFG__RESERVED0                                                   31:0
`define MCU_SWI_GP2_CFG___POR                                                32'h00000000

`define MCU_SWI_GP3_CFG                                                        'h00000040
`define MCU_SWI_GP3_CFG__RESERVED0                                                   31:0
`define MCU_SWI_GP3_CFG___POR                                                32'h00000000

`define MCU_SWI_DEBUG_CFG                                                      'h00000044
`define MCU_SWI_DEBUG_CFG__STEP                                                         2
`define MCU_SWI_DEBUG_CFG__INTR                                                         0
`define MCU_SWI_DEBUG_CFG__EXIT                                                         4
`define MCU_SWI_DEBUG_CFG___POR                                              32'h00000000

`define MCU_SWI_ITCM_CFG                                                       'h00000048
`define MCU_SWI_ITCM_CFG__TIMING_PARAM                                                7:0
`define MCU_SWI_ITCM_CFG___POR                                               32'h0000003F

`define MCU_SWI_DTCM_CFG                                                       'h0000004C
`define MCU_SWI_DTCM_CFG__TIMING_PARAM                                                7:0
`define MCU_SWI_DTCM_CFG___POR                                               32'h0000003F

`define CMN_SWI_VREF_M0_CFG                                                    'h00000008
`define CMN_SWI_VREF_M0_CFG__PWR                                                    12:11
`define CMN_SWI_VREF_M0_CFG__HIZ                                                       10
`define CMN_SWI_VREF_M0_CFG__EN                                                         9
`define CMN_SWI_VREF_M0_CFG__CTRL                                                     7:0
`define CMN_SWI_VREF_M0_CFG___POR                                            32'h00000000

`define CMN_SWI_VREF_M1_CFG                                                    'h0000000C
`define CMN_SWI_VREF_M1_CFG__PWR                                                    12:11
`define CMN_SWI_VREF_M1_CFG__HIZ                                                       10
`define CMN_SWI_VREF_M1_CFG__EN                                                         9
`define CMN_SWI_VREF_M1_CFG__CTRL                                                     7:0
`define CMN_SWI_VREF_M1_CFG___POR                                            32'h00000000

`define CMN_SWI_ZQCAL_CFG                                                      'h00000010
`define CMN_SWI_ZQCAL_CFG__PCAL                                                      13:8
`define CMN_SWI_ZQCAL_CFG__VOL_0P6_SEL                                                  7
`define CMN_SWI_ZQCAL_CFG__PD_SEL                                                       6
`define CMN_SWI_ZQCAL_CFG__CAL_EN                                                       5
`define CMN_SWI_ZQCAL_CFG__NCAL                                                       4:0
`define CMN_SWI_ZQCAL_CFG___POR                                              32'h00000000

`define CMN_SWI_ZQCAL_STA                                                      'h00000014
`define CMN_SWI_ZQCAL_STA__COMP                                                         0
`define CMN_SWI_ZQCAL_STA___POR                                              32'h00000000

`define CMN_SWI_IBIAS_CFG                                                      'h00000018
`define CMN_SWI_IBIAS_CFG__EN                                                           0
`define CMN_SWI_IBIAS_CFG___POR                                              32'h00000000

`define CMN_SWI_TEST_CFG                                                       'h0000001C
`define CMN_SWI_TEST_CFG__DTST_DIV_EN                                                  17
`define CMN_SWI_TEST_CFG__DTST_EXT_SEL                                              16:12
`define CMN_SWI_TEST_CFG__DTST_DRVR_IMPD                                             10:8
`define CMN_SWI_TEST_CFG__ATST_SEL                                                    5:2
`define CMN_SWI_TEST_CFG__ATB_MODE                                                    1:0
`define CMN_SWI_TEST_CFG___POR                                               32'h00000000

`define CMN_SWI_LDO_M0_CFG                                                     'h00000020
`define CMN_SWI_LDO_M0_CFG__HIZ                                                        13
`define CMN_SWI_LDO_M0_CFG__ATST_SEL                                                12:10
`define CMN_SWI_LDO_M0_CFG__TRAN_ENH_EN                                                 9
`define CMN_SWI_LDO_M0_CFG__EN                                                          8
`define CMN_SWI_LDO_M0_CFG__VREF_CTRL                                                 7:0
`define CMN_SWI_LDO_M0_CFG___POR                                             32'h00000000

`define CMN_SWI_LDO_M1_CFG                                                     'h00000024
`define CMN_SWI_LDO_M1_CFG__HIZ                                                        13
`define CMN_SWI_LDO_M1_CFG__ATST_SEL                                                12:10
`define CMN_SWI_LDO_M1_CFG__TRAN_ENH_EN                                                 9
`define CMN_SWI_LDO_M1_CFG__EN                                                          8
`define CMN_SWI_LDO_M1_CFG__VREF_CTRL                                                 7:0
`define CMN_SWI_LDO_M1_CFG___POR                                             32'h00000000

`define CMN_SWI_CLK_CTRL_CFG                                                   'h00000028
`define CMN_SWI_CLK_CTRL_CFG__GFCM_EN                                                   3
`define CMN_SWI_CLK_CTRL_CFG__PLL0_DIV_CLK_EN                                           2
`define CMN_SWI_CLK_CTRL_CFG__PLL0_DIV_CLK_RST                                          1
`define CMN_SWI_CLK_CTRL_CFG__PLL0_DIV_CLK_BYP                                          0
`define CMN_SWI_CLK_CTRL_CFG___POR                                           32'h00000002

`define CMN_SWI_PMON_ANA_CFG                                                   'h00000038
`define CMN_SWI_PMON_ANA_CFG__NOR_EN                                                    1
`define CMN_SWI_PMON_ANA_CFG__NAND_EN                                                   0
`define CMN_SWI_PMON_ANA_CFG___POR                                           32'h00000000

`define CMN_SWI_PMON_DIG_CFG                                                   'h0000003C
`define CMN_SWI_PMON_DIG_CFG__REFCLK_RST                                                8
`define CMN_SWI_PMON_DIG_CFG__INITWAIT                                                7:0
`define CMN_SWI_PMON_DIG_CFG___POR                                           32'h00000100

`define CMN_SWI_PMON_DIG_NAND_CFG                                              'h00000040
`define CMN_SWI_PMON_DIG_NAND_CFG__COUNT_EN                                            12
`define CMN_SWI_PMON_DIG_NAND_CFG__REFCOUNT                                          11:0
`define CMN_SWI_PMON_DIG_NAND_CFG___POR                                      32'h00000000

`define CMN_SWI_PMON_DIG_NOR_CFG                                               'h00000044
`define CMN_SWI_PMON_DIG_NOR_CFG__COUNT_EN                                             12
`define CMN_SWI_PMON_DIG_NOR_CFG__REFCOUNT                                           11:0
`define CMN_SWI_PMON_DIG_NOR_CFG___POR                                       32'h00000000

`define CMN_SWI_PMON_NAND_STA                                                  'h00000048
`define CMN_SWI_PMON_NAND_STA__DONE                                                    24
`define CMN_SWI_PMON_NAND_STA__COUNT                                                 23:0
`define CMN_SWI_PMON_NAND_STA___POR                                          32'h00000000

`define CMN_SWI_PMON_NOR_STA                                                   'h0000004C
`define CMN_SWI_PMON_NOR_STA__DONE                                                     24
`define CMN_SWI_PMON_NOR_STA__COUNT                                                  23:0
`define CMN_SWI_PMON_NOR_STA___POR                                           32'h00000000

`define CMN_SWI_CLK_STA                                                        'h00000050
`define CMN_SWI_CLK_STA__GFCM1_CLKB_SEL                                                 3
`define CMN_SWI_CLK_STA__GFCM1_CLKA_SEL                                                 2
`define CMN_SWI_CLK_STA__GFCM0_CLKB_SEL                                                 1
`define CMN_SWI_CLK_STA__GFCM0_CLKA_SEL                                                 0
`define CMN_SWI_CLK_STA___POR                                                32'h00000000

`define CMN_SWI_RSTN_CFG                                                       'h00000054
`define CMN_SWI_RSTN_CFG__RSTN_BS_ENA                                                   4
`define CMN_SWI_RSTN_CFG__RSTN_BS_DIN                                                   3
`define CMN_SWI_RSTN_CFG__RSTN_LPBK_ENA                                                 2
`define CMN_SWI_RSTN_CFG__RSTN_OVR_VAL                                                  1
`define CMN_SWI_RSTN_CFG__RSTN_OVR_SEL                                                  0
`define CMN_SWI_RSTN_CFG___POR                                               32'h00000000

`define CMN_SWI_RSTN_STA                                                       'h00000058
`define CMN_SWI_RSTN_STA__RSTN_LPBK                                                     0
`define CMN_SWI_RSTN_STA___POR                                               32'h00000000

`define CMN_PLL_MVP_PLL_CORE_OVERRIDES                                         'h00000000
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_GFCM_SEL_MUX                               6
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_GFCM_SEL                                   5
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_VCO_SEL_MUX                                4
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_VCO_SEL                                  3:2
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_RESET_MUX                                  1
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES__CORE_RESET                                      0
`define CMN_PLL_MVP_PLL_CORE_OVERRIDES___POR                                 32'h00000000

`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO                                        'h00000004
`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO__CORE_SWITCH_VCO                                0
`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO___POR                                32'h00000000

`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO_HW                                     'h00000008
`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO_HW__CORE_SWITCH_VCO_HW_MUX                      1
`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO_HW__CORE_SWITCH_VCO_HW                          0
`define CMN_PLL_MVP_PLL_CORE_SWTICH_VCO_HW___POR                             32'h00000000

`define CMN_PLL_MVP_PLL_CORE_STATUS                                            'h0000000C
`define CMN_PLL_MVP_PLL_CORE_STATUS__FSM_STATE                                      24:21
`define CMN_PLL_MVP_PLL_CORE_STATUS__FREQ_DETECT_CYCLES                              20:4
`define CMN_PLL_MVP_PLL_CORE_STATUS__FREQ_DETECT_LOCK                                   3
`define CMN_PLL_MVP_PLL_CORE_STATUS__CORE_INITIAL_SWITCH_DONE                           2
`define CMN_PLL_MVP_PLL_CORE_STATUS__CORE_FASTLOCK_READY                                1
`define CMN_PLL_MVP_PLL_CORE_STATUS__CORE_READY                                         0
`define CMN_PLL_MVP_PLL_CORE_STATUS___POR                                    32'h00000000

`define CMN_PLL_MVP_PLL_CORE_STATUS_INT                                        'h00000010
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO2_FLL_THRESHOLD                             8
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO2_FLL_LOCKED                                7
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO1_FLL_THRESHOLD                             6
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO1_FLL_LOCKED                                5
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO0_FLL_THRESHOLD                             4
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__VCO0_FLL_LOCKED                                3
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__INITIAL_SWITCH_DONE                            2
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__CORE_LOCKED                                    1
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT__LOSS_OF_LOCK                                   0
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT___POR                                32'h00000000

`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN                                     'h00000014
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO2_FLL_THRESHOLD_INT_EN                    8
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO2_FLL_LOCKED_INT_EN                      7
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO1_FLL_THRESHOLD_INT_EN                    6
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO1_FLL_LOCKED_INT_EN                      5
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO0_FLL_THRESHOLD_INT_EN                    4
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__VCO0_FLL_LOCKED_INT_EN                      3
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__INITIAL_SWITCH_DONE_INT_EN                    2
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__CORE_LOCKED_INT_EN                          1
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN__LOSS_OF_LOCK_INT_EN                         0
`define CMN_PLL_MVP_PLL_CORE_STATUS_INT_EN___POR                             32'h00000000

`define CMN_PLL_MVP_PLL_VCO0_BAND                                              'h00000018
`define CMN_PLL_MVP_PLL_VCO0_BAND__VCO0_FINE_MUX                                       14
`define CMN_PLL_MVP_PLL_VCO0_BAND__VCO0_FINE                                         13:8
`define CMN_PLL_MVP_PLL_VCO0_BAND__RESERVED0                                            7
`define CMN_PLL_MVP_PLL_VCO0_BAND__VCO0_BAND_MUX                                        6
`define CMN_PLL_MVP_PLL_VCO0_BAND__VCO0_BAND                                          5:0
`define CMN_PLL_MVP_PLL_VCO0_BAND___POR                                      32'h00005F40

`define CMN_PLL_MVP_PLL_VCO0_CONTROL                                           'h0000001C
`define CMN_PLL_MVP_PLL_VCO0_CONTROL__VCO0_BYP_CLK_SEL                                  2
`define CMN_PLL_MVP_PLL_VCO0_CONTROL__VCO0_ENA_MUX                                      1
`define CMN_PLL_MVP_PLL_VCO0_CONTROL__VCO0_ENA                                          0
`define CMN_PLL_MVP_PLL_VCO0_CONTROL___POR                                   32'h00000000

`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1                                      'h00000020
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_LOCKED                                 28
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_TOO_SLOW_STATUS                        27
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_TOO_FAST_STATUS                        26
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FLL_PERSISTENT_MODE                    25
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FLL_BYPASS_FINE                        24
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FLL_BYPASS_BAND                        23
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_LOCKED_COUNT_THRESHOLD                22:19
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_USE_DEMETED_CHECK                      18
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_DELAY_COUNT                         17:14
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FINE_START                           13:8
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_BAND_START                            7:2
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FLL_MANUAL_MODE                         1
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1__VCO0_FLL_ENABLE                              0
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL1___POR                              32'h02A49F7C

`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL2                                      'h00000024
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL2__VCO0_FLL_RANGE                           28:24
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL2__VCO0_FLL_VCO_COUNT_TARGET                 23:8
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL2__VCO0_FLL_REFCLK_COUNT                      7:0
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL2___POR                              32'h0400D008

`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL3                                      'h00000028
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL3__VCO0_FLL_BAND_THRESH                       5:0
`define CMN_PLL_MVP_PLL_VCO0_FLL_CONTROL3___POR                              32'h0000003C

`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS                                   'h0000002C
`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS__VCO0_FINE_PREV_STATUS                 23:18
`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS__VCO0_FINE_STATUS                      17:12
`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS__VCO0_BAND_PREV_STATUS                  11:6
`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS__VCO0_BAND_STATUS                        5:0
`define CMN_PLL_MVP_PLL_VCO0_FLL_BAND_STATUS___POR                           32'h00000000

`define CMN_PLL_MVP_PLL_VCO0_FLL_COUNT_STATUS                                  'h00000030
`define CMN_PLL_MVP_PLL_VCO0_FLL_COUNT_STATUS__VCO0_VCO_COUNT                        15:0
`define CMN_PLL_MVP_PLL_VCO0_FLL_COUNT_STATUS___POR                          32'h00000000

`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS                                 'h00000034
`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS__VCO0_FRAC_EN_AUTO                      26
`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS__VCO0_FRAC_EN                           25
`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS__VCO0_FRAC                            24:9
`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS__VCO0_INT                              8:0
`define CMN_PLL_MVP_PLL_VCO0_INT_FRAC_SETTINGS___POR                         32'h0400000A

`define CMN_PLL_MVP_PLL_VCO0_PROP_GAINS                                        'h00000038
`define CMN_PLL_MVP_PLL_VCO0_PROP_GAINS__VCO0_PROP_GAIN                               4:0
`define CMN_PLL_MVP_PLL_VCO0_PROP_GAINS___POR                                32'h0000000A

`define CMN_PLL_MVP_PLL_VCO1_BAND                                              'h0000003C
`define CMN_PLL_MVP_PLL_VCO1_BAND__VCO1_FINE_MUX                                       14
`define CMN_PLL_MVP_PLL_VCO1_BAND__VCO1_FINE                                         13:8
`define CMN_PLL_MVP_PLL_VCO1_BAND__RESERVED0                                            7
`define CMN_PLL_MVP_PLL_VCO1_BAND__VCO1_BAND_MUX                                        6
`define CMN_PLL_MVP_PLL_VCO1_BAND__VCO1_BAND                                          5:0
`define CMN_PLL_MVP_PLL_VCO1_BAND___POR                                      32'h00000000

`define CMN_PLL_MVP_PLL_VCO1_CONTROL                                           'h00000040
`define CMN_PLL_MVP_PLL_VCO1_CONTROL__VCO1_POST_DIV                                   4:3
`define CMN_PLL_MVP_PLL_VCO1_CONTROL__VCO1_BYP_CLK_SEL                                  2
`define CMN_PLL_MVP_PLL_VCO1_CONTROL__VCO1_ENA_MUX                                      1
`define CMN_PLL_MVP_PLL_VCO1_CONTROL__VCO1_ENA                                          0
`define CMN_PLL_MVP_PLL_VCO1_CONTROL___POR                                   32'h00000000

`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1                                      'h00000044
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_LOCKED                                 28
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_TOO_SLOW_STATUS                        27
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_TOO_FAST_STATUS                        26
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FLL_PERSISTENT_MODE                    25
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FLL_BYPASS_FINE                        24
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FLL_BYPASS_BAND                        23
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_LOCKED_COUNT_THRESHOLD                22:19
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_USE_DEMETED_CHECK                      18
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_DELAY_COUNT                         17:14
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FINE_START                           13:8
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_BAND_START                            7:2
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FLL_MANUAL_MODE                         1
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1__VCO1_FLL_ENABLE                              0
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL1___POR                              32'h00249F00

`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL2                                      'h00000048
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL2__VCO1_FLL_RANGE                           28:24
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL2__VCO1_FLL_VCO_COUNT_TARGET                 23:8
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL2__VCO1_FLL_REFCLK_COUNT                      7:0
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL2___POR                              32'h0400D008

`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL3                                      'h0000004C
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL3__VCO1_FLL_BAND_THRESH                       5:0
`define CMN_PLL_MVP_PLL_VCO1_FLL_CONTROL3___POR                              32'h0000003C

`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS                                   'h00000050
`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS__VCO1_FINE_PREV_STATUS                 23:18
`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS__VCO1_FINE_STATUS                      17:12
`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS__VCO1_BAND_PREV_STATUS                  11:6
`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS__VCO1_BAND_STATUS                        5:0
`define CMN_PLL_MVP_PLL_VCO1_FLL_BAND_STATUS___POR                           32'h00000000

`define CMN_PLL_MVP_PLL_VCO1_FLL_COUNT_STATUS                                  'h00000054
`define CMN_PLL_MVP_PLL_VCO1_FLL_COUNT_STATUS__VCO1_VCO_COUNT                        15:0
`define CMN_PLL_MVP_PLL_VCO1_FLL_COUNT_STATUS___POR                          32'h00000000

`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS                                 'h00000058
`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS__VCO1_FRAC_EN_AUTO                      26
`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS__VCO1_FRAC_EN                           25
`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS__VCO1_FRAC                            24:9
`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS__VCO1_INT                              8:0
`define CMN_PLL_MVP_PLL_VCO1_INT_FRAC_SETTINGS___POR                         32'h0400000A

`define CMN_PLL_MVP_PLL_VCO1_PROP_GAINS                                        'h0000005C
`define CMN_PLL_MVP_PLL_VCO1_PROP_GAINS__VCO1_PROP_GAIN                               4:0
`define CMN_PLL_MVP_PLL_VCO1_PROP_GAINS___POR                                32'h0000000A

`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS                                      'h00000060
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS__VCO1_SSC_CENTER_SPREAD                      29
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS__VCO1_SSC_COUNT_CYCLES                       28
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS__VCO1_SSC_AMP                             27:11
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS__VCO1_SSC_STEPSIZE                         10:1
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS__VCO1_SSC_ENABLE                              0
`define CMN_PLL_MVP_PLL_VCO1_SSC_CONTROLS___POR                              32'h00000000

`define CMN_PLL_MVP_PLL_VCO2_BAND                                              'h00000064
`define CMN_PLL_MVP_PLL_VCO2_BAND__VCO2_FINE_MUX                                       14
`define CMN_PLL_MVP_PLL_VCO2_BAND__VCO2_FINE                                         13:8
`define CMN_PLL_MVP_PLL_VCO2_BAND__RESERVED0                                            7
`define CMN_PLL_MVP_PLL_VCO2_BAND__VCO2_BAND_MUX                                        6
`define CMN_PLL_MVP_PLL_VCO2_BAND__VCO2_BAND                                          5:0
`define CMN_PLL_MVP_PLL_VCO2_BAND___POR                                      32'h00000000

`define CMN_PLL_MVP_PLL_VCO2_CONTROL                                           'h00000068
`define CMN_PLL_MVP_PLL_VCO2_CONTROL__VCO2_POST_DIV                                   4:3
`define CMN_PLL_MVP_PLL_VCO2_CONTROL__VCO2_BYP_CLK_SEL                                  2
`define CMN_PLL_MVP_PLL_VCO2_CONTROL__VCO2_ENA_MUX                                      1
`define CMN_PLL_MVP_PLL_VCO2_CONTROL__VCO2_ENA                                          0
`define CMN_PLL_MVP_PLL_VCO2_CONTROL___POR                                   32'h00000000

`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1                                      'h0000006C
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_LOCKED                                 28
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_TOO_SLOW_STATUS                        27
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_TOO_FAST_STATUS                        26
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FLL_PERSISTENT_MODE                    25
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FLL_BYPASS_FINE                        24
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FLL_BYPASS_BAND                        23
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_LOCKED_COUNT_THRESHOLD                22:19
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_USE_DEMETED_CHECK                      18
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_DELAY_COUNT                         17:14
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FINE_START                           13:8
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_BAND_START                            7:2
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FLL_MANUAL_MODE                         1
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1__VCO2_FLL_ENABLE                              0
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL1___POR                              32'h00249F00

`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL2                                      'h00000070
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL2__VCO2_FLL_RANGE                           28:24
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL2__VCO2_FLL_VCO_COUNT_TARGET                 23:8
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL2__VCO2_FLL_REFCLK_COUNT                      7:0
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL2___POR                              32'h0400D008

`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL3                                      'h00000074
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL3__VCO2_FLL_BAND_THRESH                       5:0
`define CMN_PLL_MVP_PLL_VCO2_FLL_CONTROL3___POR                              32'h0000003C

`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS                                   'h00000078
`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS__VCO2_FINE_PREV_STATUS                 23:18
`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS__VCO2_FINE_STATUS                      17:12
`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS__VCO2_BAND_PREV_STATUS                  11:6
`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS__VCO2_BAND_STATUS                        5:0
`define CMN_PLL_MVP_PLL_VCO2_FLL_BAND_STATUS___POR                           32'h00000000

`define CMN_PLL_MVP_PLL_VCO2_FLL_COUNT_STATUS                                  'h0000007C
`define CMN_PLL_MVP_PLL_VCO2_FLL_COUNT_STATUS__VCO2_VCO_COUNT                        15:0
`define CMN_PLL_MVP_PLL_VCO2_FLL_COUNT_STATUS___POR                          32'h00000000

`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS                                 'h00000080
`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS__VCO2_FRAC_EN_AUTO                      26
`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS__VCO2_FRAC_EN                           25
`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS__VCO2_FRAC                            24:9
`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS__VCO2_INT                              8:0
`define CMN_PLL_MVP_PLL_VCO2_INT_FRAC_SETTINGS___POR                         32'h0400000A

`define CMN_PLL_MVP_PLL_VCO2_PROP_GAINS                                        'h00000084
`define CMN_PLL_MVP_PLL_VCO2_PROP_GAINS__VCO2_PROP_GAIN                               4:0
`define CMN_PLL_MVP_PLL_VCO2_PROP_GAINS___POR                                32'h0000000A

`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS                                      'h00000088
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS__VCO2_SSC_CENTER_SPREAD                      29
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS__VCO2_SSC_COUNT_CYCLES                       28
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS__VCO2_SSC_AMP                             27:11
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS__VCO2_SSC_STEPSIZE                         10:1
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS__VCO2_SSC_ENABLE                              0
`define CMN_PLL_MVP_PLL_VCO2_SSC_CONTROLS___POR                              32'h00000000

`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS                                 'h0000008C
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS__FLL_INITIAL_SETTLE                  24:21
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS__DISABLE_LOCK_DET_AFTER_LOCK                   20
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS__SWITCH_COUNT                        19:16
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS__PRE_LOCKING_COUNT                    15:8
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS__BIAS_SETTLE_COUNT                     7:0
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS___POR                         32'h00810408

`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2                                'h00000090
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2__SWITCH_2_TIME                      23:16
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2__SWITCH_1_TIME                       15:8
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2__SWITCH_RESET_TIME                    7:4
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2__PRE_SWITCH_TIME                      3:0
`define CMN_PLL_MVP_PLL_STATE_MACHINE_CONTROLS2___POR                        32'h00010311

`define CMN_PLL_MVP_PLL_INTR_GAINS                                             'h00000094
`define CMN_PLL_MVP_PLL_INTR_GAINS__NORMAL_INT_GAIN                                   4:0
`define CMN_PLL_MVP_PLL_INTR_GAINS___POR                                     32'h0000000F

`define CMN_PLL_MVP_PLL_INTR_PROP_FL_GAINS                                     'h00000098
`define CMN_PLL_MVP_PLL_INTR_PROP_FL_GAINS__FL_PROP_GAIN                              9:5
`define CMN_PLL_MVP_PLL_INTR_PROP_FL_GAINS__FL_INT_GAIN                               4:0
`define CMN_PLL_MVP_PLL_INTR_PROP_FL_GAINS___POR                             32'h000003DE

`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE                               'h0000009C
`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE__PROP_GAIN_MUX                        11
`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE__PROP_GAIN                          10:6
`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE__INT_GAIN_MUX                          5
`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE__INT_GAIN                            4:0
`define CMN_PLL_MVP_PLL_INTR_PROP_GAINS_OVERRIDE___POR                       32'h0000024F

`define CMN_PLL_MVP_PLL_LOCK_DET_SETTINGS                                      'h000000A0
`define CMN_PLL_MVP_PLL_LOCK_DET_SETTINGS__LD_RANGE                                 21:16
`define CMN_PLL_MVP_PLL_LOCK_DET_SETTINGS__LD_REFCLK_CYCLES                          15:0
`define CMN_PLL_MVP_PLL_LOCK_DET_SETTINGS___POR                              32'h00040200

`define CMN_PLL_MVP_PLL_FASTLOCK_DET_SETTINGS                                  'h000000A4
`define CMN_PLL_MVP_PLL_FASTLOCK_DET_SETTINGS__FASTLD_RANGE                         21:16
`define CMN_PLL_MVP_PLL_FASTLOCK_DET_SETTINGS__FASTLD_REFCLK_CYCLES                  15:0
`define CMN_PLL_MVP_PLL_FASTLOCK_DET_SETTINGS___POR                          32'h00080100

`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET                                        'h000000A8
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__VCO_SEL_MUX                                   16
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__VCO_SEL                                    15:14
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__FBDIV_SEL_MUX                                 13
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__FBDIV_SEL                                   12:4
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__PLL_RESET_MUX                                  3
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__PLL_RESET                                      2
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__PLL_EN_MUX                                     1
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET__PLL_EN                                         0
`define CMN_PLL_MVP_PLL_ANALOG_EN_RESET___POR                                32'h00000000

`define CMN_PLL_MVP_PLL_MODE_DTST_MISC                                         'h000000AC
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__BIAS_SEL                                        8
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__DIV16EN                                         7
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__EN_LOCK_DET_MUX                                 6
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__EN_LOCK_DET                                     5
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__CP_INT_MODE                                     4
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC__BIAS_LVL                                      3:0
`define CMN_PLL_MVP_PLL_MODE_DTST_MISC___POR                                 32'h00000008

`define CMN_PLL_MVP_PLL_PROP_CTRLS                                             'h000000B0
`define CMN_PLL_MVP_PLL_PROP_CTRLS__PROP_R_CTRL                                       3:2
`define CMN_PLL_MVP_PLL_PROP_CTRLS__PROP_C_CTRL                                       1:0
`define CMN_PLL_MVP_PLL_PROP_CTRLS___POR                                     32'h00000000

`define CMN_PLL_MVP_PLL_REFCLK_CONTROLS                                        'h000000B4
`define CMN_PLL_MVP_PLL_REFCLK_CONTROLS__SEL_REFCLK_ALT                                 2
`define CMN_PLL_MVP_PLL_REFCLK_CONTROLS__PFD_MODE                                     1:0
`define CMN_PLL_MVP_PLL_REFCLK_CONTROLS___POR                                32'h00000000

`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES                                       'h000000B8
`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES__FORCE_VCO2_CLK_GATE                           3
`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES__FORCE_VCO1_CLK_GATE                           2
`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES__FORCE_VCO0_CLK_GATE                           1
`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES__FORCE_FBCLK_GATE                              0
`define CMN_PLL_MVP_PLL_CLKGATE_DISABLES___POR                               32'h00000000

`define CMN_PLL_MVP_PLL_DEBUG_BUS_CTRL                                         'h000000BC
`define CMN_PLL_MVP_PLL_DEBUG_BUS_CTRL__DEBUG_BUS_CTRL_SEL                            5:0
`define CMN_PLL_MVP_PLL_DEBUG_BUS_CTRL___POR                                 32'h00000000

`define CMN_PLL_MVP_PLL_DEBUG_BUS_STATUS                                       'h000000C0
`define CMN_PLL_MVP_PLL_DEBUG_BUS_STATUS__DEBUG_BUS_CTRL_STATUS                      31:0
`define CMN_PLL_MVP_PLL_DEBUG_BUS_STATUS___POR                               32'h00000000

`define FSW_SWI_CTRL_CFG                                                       'h00000000
`define FSW_SWI_CTRL_CFG__POST_GFMSEL_WAIT                                          19:16
`define FSW_SWI_CTRL_CFG__SWITCH_DONE_STICKY_CLR                                       12
`define FSW_SWI_CTRL_CFG__SWITCH_DONE_OVR                                              11
`define FSW_SWI_CTRL_CFG__PSTWORK_DONE_OVR                                             10
`define FSW_SWI_CTRL_CFG__PSTWORK_DONE                                                  9
`define FSW_SWI_CTRL_CFG__PREP_DONE                                                     8
`define FSW_SWI_CTRL_CFG__MSR_OVR_VAL                                                   7
`define FSW_SWI_CTRL_CFG__MSR_OVR                                                       6
`define FSW_SWI_CTRL_CFG__MSR_TOGGLE_EN                                                 5
`define FSW_SWI_CTRL_CFG__VCO_TOGGLE_EN                                                 4
`define FSW_SWI_CTRL_CFG__VCO_SEL_OVR_VAL                                             2:1
`define FSW_SWI_CTRL_CFG__VCO_SEL_OVR                                                   0
`define FSW_SWI_CTRL_CFG___POR                                               32'h00040C31

`define FSW_SWI_CTRL_STA                                                       'h00000004
`define FSW_SWI_CTRL_STA__CORE_READY                                                    4
`define FSW_SWI_CTRL_STA__CMN_MSR                                                       3
`define FSW_SWI_CTRL_STA__SWITCH_DONE                                                   2
`define FSW_SWI_CTRL_STA__VCO_SEL                                                     1:0
`define FSW_SWI_CTRL_STA___POR                                               32'h00000000

`define FSW_SWI_DEBUG_CFG                                                      'h00000008
`define FSW_SWI_DEBUG_CFG__DEBUG_BUS_SEL                                              3:0
`define FSW_SWI_DEBUG_CFG___POR                                              32'h00000000

`define FSW_SWI_CSP_0_CFG                                                      'h0000002C
`define FSW_SWI_CSP_0_CFG__PSTPIEN_WAIT                                             23:20
`define FSW_SWI_CSP_0_CFG__PSTCLKEN_WAIT                                            19:16
`define FSW_SWI_CSP_0_CFG__PSTRST_WAIT                                              15:12
`define FSW_SWI_CSP_0_CFG__RST_PULSE_WIDTH                                           11:8
`define FSW_SWI_CSP_0_CFG__PRERST_WAIT                                                7:4
`define FSW_SWI_CSP_0_CFG__PRECLKDIS_WAIT                                             3:0
`define FSW_SWI_CSP_0_CFG___POR                                              32'h00333333

`define FSW_SWI_CSP_1_CFG                                                      'h00000030
`define FSW_SWI_CSP_1_CFG__REQ_COMPLETE_STA_CLR                                         9
`define FSW_SWI_CSP_1_CFG__CLK_DISABLE_OVR_VAL                                          8
`define FSW_SWI_CSP_1_CFG__DIV_RST_OVR_VAL                                              7
`define FSW_SWI_CSP_1_CFG__PI_DISABLE_OVR_VAL                                           6
`define FSW_SWI_CSP_1_CFG__CGC_EN_OVR_VAL                                               5
`define FSW_SWI_CSP_1_CFG__REQ_COMPLETE_OVR_VAL                                         4
`define FSW_SWI_CSP_1_CFG__REQ_OVR_VAL                                                  3
`define FSW_SWI_CSP_1_CFG__CGC_EN_OVR                                                   2
`define FSW_SWI_CSP_1_CFG__REQ_COMPLETE_OVR                                             1
`define FSW_SWI_CSP_1_CFG__REQ_OVR                                                      0
`define FSW_SWI_CSP_1_CFG___POR                                              32'h00000100

`define FSW_SWI_CSP_STA                                                        'h00000034
`define FSW_SWI_CSP_STA__REQ_COMPLETE                                                   0
`define FSW_SWI_CSP_STA___POR                                                32'h00000000

`define CTRL_SWI_CLK_CFG                                                       'h00000000
`define CTRL_SWI_CLK_CFG__REF_CLK_SEL                                                   1
`define CTRL_SWI_CLK_CFG__REF_CLK_ON                                                    5
`define CTRL_SWI_CLK_CFG__REF_CLK_CGC_EN                                                9
`define CTRL_SWI_CLK_CFG__PLL_CLK_EN                                                    0
`define CTRL_SWI_CLK_CFG__MCU_GFM_SEL                                                   2
`define CTRL_SWI_CLK_CFG__MCU_CLK_CGC_EN                                                8
`define CTRL_SWI_CLK_CFG__AHB_CLK_ON                                                    4
`define CTRL_SWI_CLK_CFG__AHBCLK_DIV2_EN                                                3
`define CTRL_SWI_CLK_CFG___POR                                               32'h00000308

`define CTRL_SWI_CLK_STA                                                       'h00000004
`define CTRL_SWI_CLK_STA__MCU_GFM_SEL1                                                  1
`define CTRL_SWI_CLK_STA__MCU_GFM_SEL0                                                  0
`define CTRL_SWI_CLK_STA__DFI_CLK_ON                                                    2
`define CTRL_SWI_CLK_STA___POR                                               32'h00000000

`define CTRL_SWI_AHB_SNOOP_CFG                                                 'h00000008
`define CTRL_SWI_AHB_SNOOP_CFG__TS_RESET                                                1
`define CTRL_SWI_AHB_SNOOP_CFG__TS_ENABLE                                               0
`define CTRL_SWI_AHB_SNOOP_CFG__SNOOP_MODE                                             12
`define CTRL_SWI_AHB_SNOOP_CFG__RDATA_UPDATE                                           10
`define CTRL_SWI_AHB_SNOOP_CFG__RDATA_CLR                                               8
`define CTRL_SWI_AHB_SNOOP_CFG___POR                                         32'h00000000

`define CTRL_SWI_AHB_SNOOP_STA                                                 'h0000000C
`define CTRL_SWI_AHB_SNOOP_STA__FULL                                                    1
`define CTRL_SWI_AHB_SNOOP_STA__EMPTY                                                   0
`define CTRL_SWI_AHB_SNOOP_STA___POR                                         32'h00000000

`define CTRL_SWI_AHB_SNOOP_DATA_STA                                            'h00000010
`define CTRL_SWI_AHB_SNOOP_DATA_STA__RDATA                                           31:0
`define CTRL_SWI_AHB_SNOOP_DATA_STA___POR                                    32'h00000000

`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG                                         'h00000014
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_1_POLARITY                                  9
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_1_MODE                                  11:10
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_1_EN                                        8
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_0_POLARITY                                  1
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_0_MODE                                    3:2
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG__PAT_0_EN                                        0
`define CTRL_SWI_AHB_SNOOP_PATTERN_CFG___POR                                 32'h00000000

`define CTRL_SWI_AHB_SNOOP_PATTERN_0_CFG                                       'h00000018
`define CTRL_SWI_AHB_SNOOP_PATTERN_0_CFG__PAT_VAL                                    31:0
`define CTRL_SWI_AHB_SNOOP_PATTERN_0_CFG___POR                               32'h00000000

`define CTRL_SWI_AHB_SNOOP_PATTERN_1_CFG                                       'h0000001C
`define CTRL_SWI_AHB_SNOOP_PATTERN_1_CFG__PAT_VAL                                    31:0
`define CTRL_SWI_AHB_SNOOP_PATTERN_1_CFG___POR                               32'h00000000

`define CTRL_SWI_AHB_SNOOP_PATTERN_STA                                         'h00000020
`define CTRL_SWI_AHB_SNOOP_PATTERN_STA__PAT_1_DETECT                                    1
`define CTRL_SWI_AHB_SNOOP_PATTERN_STA__PAT_0_DETECT                                    0
`define CTRL_SWI_AHB_SNOOP_PATTERN_STA___POR                                 32'h00000000

`define CTRL_SWI_DEBUG_CFG                                                     'h00000024
`define CTRL_SWI_DEBUG_CFG__VAL                                                      31:0
`define CTRL_SWI_DEBUG_CFG___POR                                             32'h00000000

`define CTRL_SWI_DEBUG1_CFG                                                    'h00000028
`define CTRL_SWI_DEBUG1_CFG__OVR_SEL                                                    0
`define CTRL_SWI_DEBUG1_CFG___POR                                            32'h00000000

`define DFI_SWI_TOP_0_CFG                                                      'h00000000
`define DFI_SWI_TOP_0_CFG__CA_LPBK_SEL                                                  0
`define DFI_SWI_TOP_0_CFG___POR                                              32'h00000000

`define DFI_SWI_DATA_BIT_ENABLE_CFG                                            'h00000004
`define DFI_SWI_DATA_BIT_ENABLE_CFG__VAL                                             31:0
`define DFI_SWI_DATA_BIT_ENABLE_CFG___POR                                    32'h000001FF

`define DFI_SWI_PHYFREQ_RANGE_CFG                                              'h00000008
`define DFI_SWI_PHYFREQ_RANGE_CFG__VAL                                               31:0
`define DFI_SWI_PHYFREQ_RANGE_CFG___POR                                      32'h0000EFB5

`define DFI_SWI_STATUS_IF_CFG                                                  'h0000000C
`define DFI_SWI_STATUS_IF_CFG__SW_REQ_VAL                                               1
`define DFI_SWI_STATUS_IF_CFG__SW_REQ_OVR                                               0
`define DFI_SWI_STATUS_IF_CFG__SW_FREQ_RATIO_VAL                                    15:14
`define DFI_SWI_STATUS_IF_CFG__SW_FREQ_OVR                                              8
`define DFI_SWI_STATUS_IF_CFG__SW_FREQ_FSP_VAL                                      13:12
`define DFI_SWI_STATUS_IF_CFG__SW_FREQUENCY_VAL                                     20:16
`define DFI_SWI_STATUS_IF_CFG__SW_EVENT_1_VAL                                           7
`define DFI_SWI_STATUS_IF_CFG__SW_EVENT_1_OVR                                           6
`define DFI_SWI_STATUS_IF_CFG__SW_EVENT_0_VAL                                           5
`define DFI_SWI_STATUS_IF_CFG__SW_EVENT_0_OVR                                           4
`define DFI_SWI_STATUS_IF_CFG__SW_ACK_VAL                                               3
`define DFI_SWI_STATUS_IF_CFG__SW_ACK_OVR                                               2
`define DFI_SWI_STATUS_IF_CFG___POR                                          32'h0000000D

`define DFI_SWI_STATUS_IF_STA                                                  'h00000010
`define DFI_SWI_STATUS_IF_STA__REQ                                                      0
`define DFI_SWI_STATUS_IF_STA__FREQ_RATIO                                             7:6
`define DFI_SWI_STATUS_IF_STA__FREQ_FSP                                               5:4
`define DFI_SWI_STATUS_IF_STA__FREQUENCY                                             12:8
`define DFI_SWI_STATUS_IF_STA__ACK                                                      1
`define DFI_SWI_STATUS_IF_STA___POR                                          32'h00000000

`define DFI_SWI_STATUS_IF_EVENT_0_CFG                                          'h00000014
`define DFI_SWI_STATUS_IF_EVENT_0_CFG__SW_EVENT_CNT_SEL                                31
`define DFI_SWI_STATUS_IF_EVENT_0_CFG__SW_EVENT_CNT                                  19:0
`define DFI_SWI_STATUS_IF_EVENT_0_CFG___POR                                  32'h00000000

`define DFI_SWI_STATUS_IF_EVENT_1_CFG                                          'h00000018
`define DFI_SWI_STATUS_IF_EVENT_1_CFG__SW_EVENT_CNT_SEL                                31
`define DFI_SWI_STATUS_IF_EVENT_1_CFG__SW_EVENT_CNT                                  19:0
`define DFI_SWI_STATUS_IF_EVENT_1_CFG___POR                                  32'h00000000

`define DFI_SWI_CTRLUPD_IF_CFG                                                 'h0000001C
`define DFI_SWI_CTRLUPD_IF_CFG__SW_REQ_VAL                                              1
`define DFI_SWI_CTRLUPD_IF_CFG__SW_REQ_OVR                                              0
`define DFI_SWI_CTRLUPD_IF_CFG__SW_EVENT_1_VAL                                          7
`define DFI_SWI_CTRLUPD_IF_CFG__SW_EVENT_1_OVR                                          6
`define DFI_SWI_CTRLUPD_IF_CFG__SW_EVENT_0_VAL                                          5
`define DFI_SWI_CTRLUPD_IF_CFG__SW_EVENT_0_OVR                                          4
`define DFI_SWI_CTRLUPD_IF_CFG__SW_ACK_VAL                                              3
`define DFI_SWI_CTRLUPD_IF_CFG__SW_ACK_OVR                                              2
`define DFI_SWI_CTRLUPD_IF_CFG___POR                                         32'h00000000

`define DFI_SWI_CTRLUPD_IF_STA                                                 'h00000020
`define DFI_SWI_CTRLUPD_IF_STA__REQ                                                     0
`define DFI_SWI_CTRLUPD_IF_STA__ACK                                                     1
`define DFI_SWI_CTRLUPD_IF_STA___POR                                         32'h00000000

`define DFI_SWI_CTRLUPD_IF_EVENT_0_CFG                                         'h00000024
`define DFI_SWI_CTRLUPD_IF_EVENT_0_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_CTRLUPD_IF_EVENT_0_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_CTRLUPD_IF_EVENT_0_CFG___POR                                 32'h00000000

`define DFI_SWI_CTRLUPD_IF_EVENT_1_CFG                                         'h00000028
`define DFI_SWI_CTRLUPD_IF_EVENT_1_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_CTRLUPD_IF_EVENT_1_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_CTRLUPD_IF_EVENT_1_CFG___POR                                 32'h00000000

`define DFI_SWI_LP_CTRL_IF_CFG                                                 'h0000002C
`define DFI_SWI_LP_CTRL_IF_CFG__SW_REQ_VAL                                              1
`define DFI_SWI_LP_CTRL_IF_CFG__SW_REQ_OVR                                              0
`define DFI_SWI_LP_CTRL_IF_CFG__SW_EVENT_1_VAL                                          7
`define DFI_SWI_LP_CTRL_IF_CFG__SW_EVENT_1_OVR                                          6
`define DFI_SWI_LP_CTRL_IF_CFG__SW_EVENT_0_VAL                                          5
`define DFI_SWI_LP_CTRL_IF_CFG__SW_EVENT_0_OVR                                          4
`define DFI_SWI_LP_CTRL_IF_CFG__SW_ACK_VAL                                              3
`define DFI_SWI_LP_CTRL_IF_CFG__SW_ACK_OVR                                              2
`define DFI_SWI_LP_CTRL_IF_CFG___POR                                         32'h00000000

`define DFI_SWI_LP_CTRL_IF_STA                                                 'h00000030
`define DFI_SWI_LP_CTRL_IF_STA__WAKEUP                                                9:4
`define DFI_SWI_LP_CTRL_IF_STA__REQ                                                     0
`define DFI_SWI_LP_CTRL_IF_STA__ACK                                                     1
`define DFI_SWI_LP_CTRL_IF_STA___POR                                         32'h00000000

`define DFI_SWI_LP_CTRL_IF_EVENT_0_CFG                                         'h00000034
`define DFI_SWI_LP_CTRL_IF_EVENT_0_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_LP_CTRL_IF_EVENT_0_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_LP_CTRL_IF_EVENT_0_CFG___POR                                 32'h00000000

`define DFI_SWI_LP_CTRL_IF_EVENT_1_CFG                                         'h00000038
`define DFI_SWI_LP_CTRL_IF_EVENT_1_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_LP_CTRL_IF_EVENT_1_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_LP_CTRL_IF_EVENT_1_CFG___POR                                 32'h00000000

`define DFI_SWI_LP_DATA_IF_CFG                                                 'h0000003C
`define DFI_SWI_LP_DATA_IF_CFG__SW_REQ_VAL                                              1
`define DFI_SWI_LP_DATA_IF_CFG__SW_REQ_OVR                                              0
`define DFI_SWI_LP_DATA_IF_CFG__SW_EVENT_1_VAL                                          7
`define DFI_SWI_LP_DATA_IF_CFG__SW_EVENT_1_OVR                                          6
`define DFI_SWI_LP_DATA_IF_CFG__SW_EVENT_0_VAL                                          5
`define DFI_SWI_LP_DATA_IF_CFG__SW_EVENT_0_OVR                                          4
`define DFI_SWI_LP_DATA_IF_CFG__SW_ACK_VAL                                              3
`define DFI_SWI_LP_DATA_IF_CFG__SW_ACK_OVR                                              2
`define DFI_SWI_LP_DATA_IF_CFG___POR                                         32'h00000000

`define DFI_SWI_LP_DATA_IF_STA                                                 'h00000040
`define DFI_SWI_LP_DATA_IF_STA__WAKEUP                                                9:4
`define DFI_SWI_LP_DATA_IF_STA__REQ                                                     0
`define DFI_SWI_LP_DATA_IF_STA__ACK                                                     1
`define DFI_SWI_LP_DATA_IF_STA___POR                                         32'h00000000

`define DFI_SWI_LP_DATA_IF_EVENT_0_CFG                                         'h00000044
`define DFI_SWI_LP_DATA_IF_EVENT_0_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_LP_DATA_IF_EVENT_0_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_LP_DATA_IF_EVENT_0_CFG___POR                                 32'h00000000

`define DFI_SWI_LP_DATA_IF_EVENT_1_CFG                                         'h00000048
`define DFI_SWI_LP_DATA_IF_EVENT_1_CFG__SW_EVENT_CNT_SEL                               31
`define DFI_SWI_LP_DATA_IF_EVENT_1_CFG__SW_EVENT_CNT                                 19:0
`define DFI_SWI_LP_DATA_IF_EVENT_1_CFG___POR                                 32'h00000000

`define DFI_SWI_PHYUPD_IF_CFG                                                  'h0000004C
`define DFI_SWI_PHYUPD_IF_CFG__SW_TYPE                                                9:8
`define DFI_SWI_PHYUPD_IF_CFG__SW_REQ_VAL                                               1
`define DFI_SWI_PHYUPD_IF_CFG__SW_REQ_OVR                                               0
`define DFI_SWI_PHYUPD_IF_CFG__SW_EVENT_VAL                                             5
`define DFI_SWI_PHYUPD_IF_CFG__SW_EVENT_OVR                                             4
`define DFI_SWI_PHYUPD_IF_CFG__SW_ACK_VAL                                               3
`define DFI_SWI_PHYUPD_IF_CFG__SW_ACK_OVR                                               2
`define DFI_SWI_PHYUPD_IF_CFG___POR                                          32'h00000000

`define DFI_SWI_PHYUPD_IF_STA                                                  'h00000050
`define DFI_SWI_PHYUPD_IF_STA__REQ                                                      0
`define DFI_SWI_PHYUPD_IF_STA__EVENT                                                    2
`define DFI_SWI_PHYUPD_IF_STA__ACK                                                      1
`define DFI_SWI_PHYUPD_IF_STA___POR                                          32'h00000000

`define DFI_SWI_PHYMSTR_IF_CFG                                                 'h00000054
`define DFI_SWI_PHYMSTR_IF_CFG__SW_TYPE                                              10:9
`define DFI_SWI_PHYMSTR_IF_CFG__SW_STATE_SEL                                            6
`define DFI_SWI_PHYMSTR_IF_CFG__SW_REQ_VAL                                              1
`define DFI_SWI_PHYMSTR_IF_CFG__SW_REQ_OVR                                              0
`define DFI_SWI_PHYMSTR_IF_CFG__SW_EVENT_VAL                                            5
`define DFI_SWI_PHYMSTR_IF_CFG__SW_EVENT_OVR                                            4
`define DFI_SWI_PHYMSTR_IF_CFG__SW_CS_STATE                                           8:7
`define DFI_SWI_PHYMSTR_IF_CFG__SW_ACK_VAL                                              3
`define DFI_SWI_PHYMSTR_IF_CFG__SW_ACK_OVR                                              2
`define DFI_SWI_PHYMSTR_IF_CFG___POR                                         32'h00000000

`define DFI_SWI_PHYMSTR_IF_STA                                                 'h00000058
`define DFI_SWI_PHYMSTR_IF_STA__REQ                                                     0
`define DFI_SWI_PHYMSTR_IF_STA__EVENT                                                   2
`define DFI_SWI_PHYMSTR_IF_STA__ACK                                                     1
`define DFI_SWI_PHYMSTR_IF_STA___POR                                         32'h00000000

`define DFI_SWI_DEBUG_CFG                                                      'h0000005C
`define DFI_SWI_DEBUG_CFG__DEBUG_BUS_SEL                                              3:0
`define DFI_SWI_DEBUG_CFG___POR                                              32'h00000000

`define DFICH0_SWI_TOP_1_CFG                                                   'h00000000
`define DFICH0_SWI_TOP_1_CFG__WDATA_UPDATE                                              7
`define DFICH0_SWI_TOP_1_CFG__WDATA_HOLD                                                5
`define DFICH0_SWI_TOP_1_CFG__WDATA_ENABLE                                              6
`define DFICH0_SWI_TOP_1_CFG__WDATA_CLR                                                 4
`define DFICH0_SWI_TOP_1_CFG__WCK_MODE                                                 16
`define DFICH0_SWI_TOP_1_CFG__TS_RESET                                                  1
`define DFICH0_SWI_TOP_1_CFG__TS_ENABLE                                                 0
`define DFICH0_SWI_TOP_1_CFG__RDOUT_EN_OVR_SEL                                         18
`define DFICH0_SWI_TOP_1_CFG__RDOUT_EN_OVR                                             19
`define DFICH0_SWI_TOP_1_CFG__RDATA_UPDATE                                             10
`define DFICH0_SWI_TOP_1_CFG__RDATA_ENABLE                                              9
`define DFICH0_SWI_TOP_1_CFG__RDATA_CLR                                                 8
`define DFICH0_SWI_TOP_1_CFG__DQBYTE_RDVALID_MASK                                   31:28
`define DFICH0_SWI_TOP_1_CFG__CA_RDDATA_EN                                             17
`define DFICH0_SWI_TOP_1_CFG__BUF_MODE                                                 12
`define DFICH0_SWI_TOP_1_CFG__BUF_CLK_EN                                               13
`define DFICH0_SWI_TOP_1_CFG___POR                                           32'h00002000

`define DFICH0_SWI_TOP_2_CFG                                                   'h00000004
`define DFICH0_SWI_TOP_2_CFG__IG_STOP_PTR                                            13:8
`define DFICH0_SWI_TOP_2_CFG__IG_START_PTR                                          21:16
`define DFICH0_SWI_TOP_2_CFG__IG_NUM_LOOPS                                            7:4
`define DFICH0_SWI_TOP_2_CFG__IG_LOOP_MODE                                              0
`define DFICH0_SWI_TOP_2_CFG__IG_LOAD_PTR                                               1
`define DFICH0_SWI_TOP_2_CFG___POR                                           32'h00000010

`define DFICH0_SWI_TOP_3_CFG                                                   'h00000008
`define DFICH0_SWI_TOP_3_CFG__TS_BRKPT_VAL                                           15:0
`define DFICH0_SWI_TOP_3_CFG__TS_BRKPT_EN                                              16
`define DFICH0_SWI_TOP_3_CFG___POR                                           32'h00000000

`define DFICH0_SWI_TOP_STA                                                     'h0000000C
`define DFICH0_SWI_TOP_STA__IG_STATE_UPD                                                2
`define DFICH0_SWI_TOP_STA__IG_STATE                                                  1:0
`define DFICH0_SWI_TOP_STA__EG_STATE_UPD                                                6
`define DFICH0_SWI_TOP_STA__EG_STATE                                                  5:4
`define DFICH0_SWI_TOP_STA___POR                                             32'h00000000

`define DFICH0_SWI_IG_DATA_CFG                                                 'h00000010
`define DFICH0_SWI_IG_DATA_CFG__WDATA                                                31:0
`define DFICH0_SWI_IG_DATA_CFG___POR                                         32'h00000000

`define DFICH0_SWI_EG_DATA_STA                                                 'h00000014
`define DFICH0_SWI_EG_DATA_STA__RDATA                                                31:0
`define DFICH0_SWI_EG_DATA_STA___POR                                         32'h00000000

`define DFICH0_SWI_WRC_M0_CFG                                                  'h00000018
`define DFICH0_SWI_WRC_M0_CFG__POST_GB_FC_DLY                                         5:4
`define DFICH0_SWI_WRC_M0_CFG__PIPE_EN                                                  0
`define DFICH0_SWI_WRC_M0_CFG__GB_MODE                                              15:12
`define DFICH0_SWI_WRC_M0_CFG___POR                                          32'h00005000

`define DFICH0_SWI_WRC_M1_CFG                                                  'h0000001C
`define DFICH0_SWI_WRC_M1_CFG__POST_GB_FC_DLY                                         5:4
`define DFICH0_SWI_WRC_M1_CFG__PIPE_EN                                                  0
`define DFICH0_SWI_WRC_M1_CFG__GB_MODE                                              15:12
`define DFICH0_SWI_WRC_M1_CFG___POR                                          32'h00005000

`define DFICH0_SWI_WRCCTRL_M0_CFG                                              'h00000020
`define DFICH0_SWI_WRCCTRL_M0_CFG__POST_GB_FC_DLY                                     5:4
`define DFICH0_SWI_WRCCTRL_M0_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WRCCTRL_M0_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WRCCTRL_M0_CFG___POR                                      32'h00005000

`define DFICH0_SWI_WRCCTRL_M1_CFG                                              'h00000024
`define DFICH0_SWI_WRCCTRL_M1_CFG__POST_GB_FC_DLY                                     5:4
`define DFICH0_SWI_WRCCTRL_M1_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WRCCTRL_M1_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WRCCTRL_M1_CFG___POR                                      32'h00005000

`define DFICH0_SWI_CKCTRL_M0_CFG                                               'h00000028
`define DFICH0_SWI_CKCTRL_M0_CFG__POST_GB_FC_DLY                                      5:4
`define DFICH0_SWI_CKCTRL_M0_CFG__PIPE_EN                                               0
`define DFICH0_SWI_CKCTRL_M0_CFG__GB_MODE                                           15:12
`define DFICH0_SWI_CKCTRL_M0_CFG___POR                                       32'h00005000

`define DFICH0_SWI_CKCTRL_M1_CFG                                               'h0000002C
`define DFICH0_SWI_CKCTRL_M1_CFG__POST_GB_FC_DLY                                      5:4
`define DFICH0_SWI_CKCTRL_M1_CFG__PIPE_EN                                               0
`define DFICH0_SWI_CKCTRL_M1_CFG__GB_MODE                                           15:12
`define DFICH0_SWI_CKCTRL_M1_CFG___POR                                       32'h00005000

`define DFICH0_SWI_RDC_M0_CFG                                                  'h00000030
`define DFICH0_SWI_RDC_M0_CFG__GB_MODE                                                3:0
`define DFICH0_SWI_RDC_M0_CFG___POR                                          32'h00000006

`define DFICH0_SWI_RDC_M1_CFG                                                  'h00000034
`define DFICH0_SWI_RDC_M1_CFG__GB_MODE                                                3:0
`define DFICH0_SWI_RDC_M1_CFG___POR                                          32'h00000006

`define DFICH0_SWI_RCTRL_M0_CFG                                                'h00000038
`define DFICH0_SWI_RCTRL_M0_CFG__POST_GB_FC_DLY                                       6:4
`define DFICH0_SWI_RCTRL_M0_CFG__PIPE_EN                                                0
`define DFICH0_SWI_RCTRL_M0_CFG__GB_MODE                                            15:12
`define DFICH0_SWI_RCTRL_M0_CFG___POR                                        32'h00005000

`define DFICH0_SWI_RCTRL_M1_CFG                                                'h0000003C
`define DFICH0_SWI_RCTRL_M1_CFG__POST_GB_FC_DLY                                       6:4
`define DFICH0_SWI_RCTRL_M1_CFG__PIPE_EN                                                0
`define DFICH0_SWI_RCTRL_M1_CFG__GB_MODE                                            15:12
`define DFICH0_SWI_RCTRL_M1_CFG___POR                                        32'h00005000

`define DFICH0_SWI_WCTRL_M0_CFG                                                'h00000040
`define DFICH0_SWI_WCTRL_M0_CFG__POST_GB_FC_DLY                                       6:4
`define DFICH0_SWI_WCTRL_M0_CFG__PIPE_EN                                                0
`define DFICH0_SWI_WCTRL_M0_CFG__GB_MODE                                            15:12
`define DFICH0_SWI_WCTRL_M0_CFG___POR                                        32'h00005000

`define DFICH0_SWI_WCTRL_M1_CFG                                                'h00000044
`define DFICH0_SWI_WCTRL_M1_CFG__POST_GB_FC_DLY                                       6:4
`define DFICH0_SWI_WCTRL_M1_CFG__PIPE_EN                                                0
`define DFICH0_SWI_WCTRL_M1_CFG__GB_MODE                                            15:12
`define DFICH0_SWI_WCTRL_M1_CFG___POR                                        32'h00005000

`define DFICH0_SWI_WENCTRL_M0_CFG                                              'h00000048
`define DFICH0_SWI_WENCTRL_M0_CFG__POST_GB_FC_DLY                                     7:4
`define DFICH0_SWI_WENCTRL_M0_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WENCTRL_M0_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WENCTRL_M0_CFG___POR                                      32'h00005000

`define DFICH0_SWI_WENCTRL_M1_CFG                                              'h0000004C
`define DFICH0_SWI_WENCTRL_M1_CFG__POST_GB_FC_DLY                                     7:4
`define DFICH0_SWI_WENCTRL_M1_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WENCTRL_M1_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WENCTRL_M1_CFG___POR                                      32'h00005000

`define DFICH0_SWI_WCKCTRL_M0_CFG                                              'h00000050
`define DFICH0_SWI_WCKCTRL_M0_CFG__POST_GB_FC_DLY                                     6:4
`define DFICH0_SWI_WCKCTRL_M0_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WCKCTRL_M0_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WCKCTRL_M0_CFG___POR                                      32'h00005000

`define DFICH0_SWI_WCKCTRL_M1_CFG                                              'h00000054
`define DFICH0_SWI_WCKCTRL_M1_CFG__POST_GB_FC_DLY                                     6:4
`define DFICH0_SWI_WCKCTRL_M1_CFG__PIPE_EN                                              0
`define DFICH0_SWI_WCKCTRL_M1_CFG__GB_MODE                                          15:12
`define DFICH0_SWI_WCKCTRL_M1_CFG___POR                                      32'h00005000

`define DFICH0_SWI_WRD_M0_CFG                                                  'h00000058
`define DFICH0_SWI_WRD_M0_CFG__POST_GB_FC_DLY                                         5:4
`define DFICH0_SWI_WRD_M0_CFG__PIPE_EN                                                  0
`define DFICH0_SWI_WRD_M0_CFG__GB_MODE                                              15:12
`define DFICH0_SWI_WRD_M0_CFG___POR                                          32'h00005000

`define DFICH0_SWI_WRD_M1_CFG                                                  'h0000005C
`define DFICH0_SWI_WRD_M1_CFG__POST_GB_FC_DLY                                         5:4
`define DFICH0_SWI_WRD_M1_CFG__PIPE_EN                                                  0
`define DFICH0_SWI_WRD_M1_CFG__GB_MODE                                              15:12
`define DFICH0_SWI_WRD_M1_CFG___POR                                          32'h00005000

`define DFICH0_SWI_RDD_M0_CFG                                                  'h00000060
`define DFICH0_SWI_RDD_M0_CFG__GB_MODE                                                3:0
`define DFICH0_SWI_RDD_M0_CFG___POR                                          32'h00000006

`define DFICH0_SWI_RDD_M1_CFG                                                  'h00000064
`define DFICH0_SWI_RDD_M1_CFG__GB_MODE                                                3:0
`define DFICH0_SWI_RDD_M1_CFG___POR                                          32'h00000006

`define DFICH0_SWI_CTRL0_M0_CFG                                                'h00000068
`define DFICH0_SWI_CTRL0_M0_CFG__WR_INTF_PIPE_EN                                        0
`define DFICH0_SWI_CTRL0_M0_CFG__RD_INTF_PIPE_EN                                        1
`define DFICH0_SWI_CTRL0_M0_CFG___POR                                        32'h00000003

`define DFICH0_SWI_CTRL0_M1_CFG                                                'h0000006C
`define DFICH0_SWI_CTRL0_M1_CFG__WR_INTF_PIPE_EN                                        0
`define DFICH0_SWI_CTRL0_M1_CFG__RD_INTF_PIPE_EN                                        1
`define DFICH0_SWI_CTRL0_M1_CFG___POR                                        32'h00000003

`define DFICH0_SWI_CTRL1_M0_CFG                                                'h00000070
`define DFICH0_SWI_CTRL1_M0_CFG__DQ_WRTRAFFIC_OVR_SEL                                   0
`define DFICH0_SWI_CTRL1_M0_CFG__DQ_WRTRAFFIC_OVR                                       4
`define DFICH0_SWI_CTRL1_M0_CFG__DQ_RDTRAFFIC_OVR_SEL                                   8
`define DFICH0_SWI_CTRL1_M0_CFG__DQ_RDTRAFFIC_OVR                                       9
`define DFICH0_SWI_CTRL1_M0_CFG__DQS_WRTRAFFIC_OVR_SEL                                  1
`define DFICH0_SWI_CTRL1_M0_CFG__DQS_WRTRAFFIC_OVR                                      5
`define DFICH0_SWI_CTRL1_M0_CFG__CK_TRAFFIC_OVR_SEL                                     3
`define DFICH0_SWI_CTRL1_M0_CFG__CK_TRAFFIC_OVR                                         7
`define DFICH0_SWI_CTRL1_M0_CFG__CA_TRAFFIC_OVR_SEL                                     2
`define DFICH0_SWI_CTRL1_M0_CFG__CA_TRAFFIC_OVR                                         6
`define DFICH0_SWI_CTRL1_M0_CFG___POR                                        32'h000000FF

`define DFICH0_SWI_CTRL1_M1_CFG                                                'h00000074
`define DFICH0_SWI_CTRL1_M1_CFG__DQ_WRTRAFFIC_OVR_SEL                                   0
`define DFICH0_SWI_CTRL1_M1_CFG__DQ_WRTRAFFIC_OVR                                       4
`define DFICH0_SWI_CTRL1_M1_CFG__DQ_RDTRAFFIC_OVR_SEL                                   8
`define DFICH0_SWI_CTRL1_M1_CFG__DQ_RDTRAFFIC_OVR                                       9
`define DFICH0_SWI_CTRL1_M1_CFG__DQS_WRTRAFFIC_OVR_SEL                                  1
`define DFICH0_SWI_CTRL1_M1_CFG__DQS_WRTRAFFIC_OVR                                      5
`define DFICH0_SWI_CTRL1_M1_CFG__CK_TRAFFIC_OVR_SEL                                     3
`define DFICH0_SWI_CTRL1_M1_CFG__CK_TRAFFIC_OVR                                         7
`define DFICH0_SWI_CTRL1_M1_CFG__CA_TRAFFIC_OVR_SEL                                     2
`define DFICH0_SWI_CTRL1_M1_CFG__CA_TRAFFIC_OVR                                         6
`define DFICH0_SWI_CTRL1_M1_CFG___POR                                        32'h000000FF

`define DFICH0_SWI_CTRL2_M0_CFG                                                'h00000078
`define DFICH0_SWI_CTRL2_M0_CFG__RDCLK_EN_PULSE_EXT                                 19:16
`define DFICH0_SWI_CTRL2_M0_CFG__DQ_WRCLK_EN_PULSE_EXT                                3:0
`define DFICH0_SWI_CTRL2_M0_CFG__DQS_WRCLK_EN_PULSE_EXT                               7:4
`define DFICH0_SWI_CTRL2_M0_CFG__CK_CLK_EN_PULSE_EXT                                15:12
`define DFICH0_SWI_CTRL2_M0_CFG__CA_CLK_EN_PULSE_EXT                                 11:8
`define DFICH0_SWI_CTRL2_M0_CFG___POR                                        32'h000F0033

`define DFICH0_SWI_CTRL2_M1_CFG                                                'h0000007C
`define DFICH0_SWI_CTRL2_M1_CFG__RDCLK_EN_PULSE_EXT                                 19:16
`define DFICH0_SWI_CTRL2_M1_CFG__DQ_WRCLK_EN_PULSE_EXT                                3:0
`define DFICH0_SWI_CTRL2_M1_CFG__DQS_WRCLK_EN_PULSE_EXT                               7:4
`define DFICH0_SWI_CTRL2_M1_CFG__CK_CLK_EN_PULSE_EXT                                15:12
`define DFICH0_SWI_CTRL2_M1_CFG__CA_CLK_EN_PULSE_EXT                                 11:8
`define DFICH0_SWI_CTRL2_M1_CFG___POR                                        32'h000F0033

`define DFICH0_SWI_CTRL3_M0_CFG                                                'h00000080
`define DFICH0_SWI_CTRL3_M0_CFG__WRD_OE_PHASE_EXT                                   21:16
`define DFICH0_SWI_CTRL3_M0_CFG__WRD_EN_PHASE_EXT                                    13:8
`define DFICH0_SWI_CTRL3_M0_CFG__WRD_CS_PHASE_EXT                                     5:0
`define DFICH0_SWI_CTRL3_M0_CFG___POR                                        32'h00020200

`define DFICH0_SWI_CTRL3_M1_CFG                                                'h00000084
`define DFICH0_SWI_CTRL3_M1_CFG__WRD_OE_PHASE_EXT                                   21:16
`define DFICH0_SWI_CTRL3_M1_CFG__WRD_EN_PHASE_EXT                                    13:8
`define DFICH0_SWI_CTRL3_M1_CFG__WRD_CS_PHASE_EXT                                     5:0
`define DFICH0_SWI_CTRL3_M1_CFG___POR                                        32'h00020200

`define DFICH0_SWI_CTRL4_M0_CFG                                                'h00000088
`define DFICH0_SWI_CTRL4_M0_CFG__WCK_OE_PHASE_EXT                                     5:0
`define DFICH0_SWI_CTRL4_M0_CFG__WCK_CS_PHASE_EXT                                    13:8
`define DFICH0_SWI_CTRL4_M0_CFG___POR                                        32'h00000002

`define DFICH0_SWI_CTRL4_M1_CFG                                                'h0000008C
`define DFICH0_SWI_CTRL4_M1_CFG__WCK_OE_PHASE_EXT                                     5:0
`define DFICH0_SWI_CTRL4_M1_CFG__WCK_CS_PHASE_EXT                                    13:8
`define DFICH0_SWI_CTRL4_M1_CFG___POR                                        32'h00000002

`define DFICH0_SWI_CTRL5_M0_CFG                                                'h00000090
`define DFICH0_SWI_CTRL5_M0_CFG__RE_PHASE_EXT                                       21:16
`define DFICH0_SWI_CTRL5_M0_CFG__REN_PHASE_EXT                                      29:24
`define DFICH0_SWI_CTRL5_M0_CFG__RCS_PHASE_EXT                                        5:0
`define DFICH0_SWI_CTRL5_M0_CFG__IE_PHASE_EXT                                        13:8
`define DFICH0_SWI_CTRL5_M0_CFG___POR                                        32'h00000000

`define DFICH0_SWI_CTRL5_M1_CFG                                                'h00000094
`define DFICH0_SWI_CTRL5_M1_CFG__RE_PHASE_EXT                                       21:16
`define DFICH0_SWI_CTRL5_M1_CFG__REN_PHASE_EXT                                      29:24
`define DFICH0_SWI_CTRL5_M1_CFG__RCS_PHASE_EXT                                        5:0
`define DFICH0_SWI_CTRL5_M1_CFG__IE_PHASE_EXT                                        13:8
`define DFICH0_SWI_CTRL5_M1_CFG___POR                                        32'h00000000

`define CH0_DQ0_SWI_TOP_CFG                                                    'h00000000
`define CH0_DQ0_SWI_TOP_CFG__WCS_SW_OVR_VAL                                             1
`define CH0_DQ0_SWI_TOP_CFG__WCS_SW_OVR                                                 0
`define CH0_DQ0_SWI_TOP_CFG__TRAINING_MODE                                              9
`define CH0_DQ0_SWI_TOP_CFG__RCS_SW_OVR_VAL                                             3
`define CH0_DQ0_SWI_TOP_CFG__RCS_SW_OVR                                                 2
`define CH0_DQ0_SWI_TOP_CFG__FIFO_CLR                                                   8
`define CH0_DQ0_SWI_TOP_CFG___POR                                            32'h00000000

`define CH0_DQ0_SWI_TOP_STA                                                    'h00000004
`define CH0_DQ0_SWI_TOP_STA__WCS                                                        0
`define CH0_DQ0_SWI_TOP_STA__RCS                                                        1
`define CH0_DQ0_SWI_TOP_STA___POR                                            32'h00000000

`define CH0_DQ0_SWI_DQ_RX_BSCAN_STA                                            'h00000008
`define CH0_DQ0_SWI_DQ_RX_BSCAN_STA__VAL                                              8:0
`define CH0_DQ0_SWI_DQ_RX_BSCAN_STA___POR                                    32'h00000000

`define CH0_DQ0_SWI_DQ_RX_M0_CFG                                               'h0000000C
`define CH0_DQ0_SWI_DQ_RX_M0_CFG__RGB_MODE                                            2:0
`define CH0_DQ0_SWI_DQ_RX_M0_CFG__FGB_MODE                                            7:4
`define CH0_DQ0_SWI_DQ_RX_M0_CFG___POR                                       32'h00000074

`define CH0_DQ0_SWI_DQ_RX_M1_CFG                                               'h00000010
`define CH0_DQ0_SWI_DQ_RX_M1_CFG__RGB_MODE                                            2:0
`define CH0_DQ0_SWI_DQ_RX_M1_CFG__FGB_MODE                                            7:4
`define CH0_DQ0_SWI_DQ_RX_M1_CFG___POR                                       32'h00000074

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0                                       'h00000014
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1                                       'h00000018
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2                                       'h0000001C
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3                                       'h00000020
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4                                       'h00000024
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5                                       'h00000028
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6                                       'h0000002C
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7                                       'h00000030
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8                                       'h00000034
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0                                       'h00000038
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1                                       'h0000003C
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2                                       'h00000040
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3                                       'h00000044
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4                                       'h00000048
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5                                       'h0000004C
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6                                       'h00000050
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7                                       'h00000054
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8                                       'h00000058
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0                                       'h0000005C
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1                                       'h00000060
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2                                       'h00000064
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3                                       'h00000068
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4                                       'h0000006C
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5                                       'h00000070
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6                                       'h00000074
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7                                       'h00000078
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8                                       'h0000007C
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0                                       'h00000080
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1                                       'h00000084
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2                                       'h00000088
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3                                       'h0000008C
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4                                       'h00000090
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5                                       'h00000094
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6                                       'h00000098
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7                                       'h0000009C
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8                                       'h000000A0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                   7:0
`define CH0_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_IO_STA                                               'h000000A4
`define CH0_DQ0_SWI_DQ_RX_IO_STA__CORE_IG                                            31:0
`define CH0_DQ0_SWI_DQ_RX_IO_STA___POR                                       32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0                                       'h000000A8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1                                       'h000000AC
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2                                       'h000000B0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3                                       'h000000B4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4                                       'h000000B8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5                                       'h000000BC
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6                                       'h000000C0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7                                       'h000000C4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8                                       'h000000C8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0                                       'h000000CC
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1                                       'h000000D0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2                                       'h000000D4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3                                       'h000000D8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4                                       'h000000DC
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5                                       'h000000E0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6                                       'h000000E4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7                                       'h000000E8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8                                       'h000000EC
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0                                       'h000000F0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1                                       'h000000F4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2                                       'h000000F8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3                                       'h000000FC
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4                                       'h00000100
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5                                       'h00000104
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6                                       'h00000108
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7                                       'h0000010C
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8                                       'h00000110
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0                                       'h00000114
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1                                       'h00000118
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2                                       'h0000011C
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3                                       'h00000120
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4                                       'h00000124
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5                                       'h00000128
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6                                       'h0000012C
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7                                       'h00000130
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8                                       'h00000134
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                   'h00000138
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                   'h0000013C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                   'h00000140
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                   'h00000144
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                   'h00000148
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                   'h0000014C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                   'h00000150
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                   'h00000154
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                   'h00000158
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                   'h0000015C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                   'h00000160
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                   'h00000164
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                   'h00000168
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                   'h0000016C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                   'h00000170
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                   'h00000174
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                   'h00000178
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                   'h0000017C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                   'h00000180
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                   'h00000184
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                   'h00000188
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                   'h0000018C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                   'h00000190
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                   'h00000194
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                   'h00000198
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                   'h0000019C
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                   'h000001A0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                   'h000001A4
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                   'h000001A8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                   'h000001AC
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                   'h000001B0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                   'h000001B4
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                   'h000001B8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                   'h000001BC
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                   'h000001C0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                   'h000001C4
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                 9:8
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                              25:24
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                              17:16
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                  1:0
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                               15:10
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                              31:26
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                              23:18
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                  7:2
`define CH0_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                           32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_0                                             'h000001C8
`define CH0_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_0___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_1                                             'h000001CC
`define CH0_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_1___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_2                                             'h000001D0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_2___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_3                                             'h000001D4
`define CH0_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_3___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_4                                             'h000001D8
`define CH0_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_4___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_5                                             'h000001DC
`define CH0_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_5___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_6                                             'h000001E0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_6___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_7                                             'h000001E4
`define CH0_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_7___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_RX_SA_STA_8                                             'h000001E8
`define CH0_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                           1
`define CH0_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                          3
`define CH0_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                          2
`define CH0_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                            0
`define CH0_DQ0_SWI_DQ_RX_SA_STA_8___POR                                     32'h00000000

`define CH0_DQ0_SWI_DQ_TX_BSCAN_CFG                                            'h000001EC
`define CH0_DQ0_SWI_DQ_TX_BSCAN_CFG__VAL                                              8:0
`define CH0_DQ0_SWI_DQ_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                  'h000001F0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                  'h000001F4
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                  'h000001F8
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                  'h000001FC
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                  'h00000200
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                  'h00000204
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                  'h00000208
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                  'h0000020C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                  'h00000210
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                  'h00000214
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                  'h00000218
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                  'h0000021C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                  'h00000220
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                  'h00000224
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                  'h00000228
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                  'h0000022C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                  'h00000230
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                  'h00000234
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                            5:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                          32'h00000001

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                  'h00000238
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                  'h0000023C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                  'h00000240
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                  'h00000244
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                  'h00000248
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                  'h0000024C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                  'h00000250
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                  'h00000254
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                  'h00000258
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                  'h0000025C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                  'h00000260
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                  'h00000264
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                  'h00000268
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                  'h0000026C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                  'h00000270
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                  'h00000274
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                  'h00000278
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                  'h0000027C
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                            6:0
`define CH0_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                          32'h00000002

`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                     'h00000280
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                     'h00000284
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                     'h00000288
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                     'h0000028C
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                   'h00000290
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                   'h00000294
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                   'h00000298
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                   'h0000029C
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                   'h000002A0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                   'h000002A4
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                   'h000002A8
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                   'h000002AC
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                   'h000002B0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                   'h000002B4
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                   'h000002B8
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                   'h000002BC
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                   'h000002C0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                   'h000002C4
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                   'h000002C8
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                   'h000002CC
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG                                      'h000002D0
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG                                      'h000002D4
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG                                      'h000002D8
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG                                      'h000002DC
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH0_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH0_DQ0_SWI_DQ_TX_RT_M0_R0_CFG                                         'h000002E0
`define CH0_DQ0_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       8:0
`define CH0_DQ0_SWI_DQ_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH0_DQ0_SWI_DQ_TX_RT_M0_R1_CFG                                         'h000002E4
`define CH0_DQ0_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       8:0
`define CH0_DQ0_SWI_DQ_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH0_DQ0_SWI_DQ_TX_RT_M1_R0_CFG                                         'h000002E8
`define CH0_DQ0_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       8:0
`define CH0_DQ0_SWI_DQ_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH0_DQ0_SWI_DQ_TX_RT_M1_R1_CFG                                         'h000002EC
`define CH0_DQ0_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       8:0
`define CH0_DQ0_SWI_DQ_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0                                      'h000002F0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1                                      'h000002F4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2                                      'h000002F8
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3                                      'h000002FC
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4                                      'h00000300
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5                                      'h00000304
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6                                      'h00000308
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7                                      'h0000030C
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8                                      'h00000310
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0                                      'h00000314
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1                                      'h00000318
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2                                      'h0000031C
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3                                      'h00000320
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4                                      'h00000324
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5                                      'h00000328
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6                                      'h0000032C
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7                                      'h00000330
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8                                      'h00000334
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0                                      'h00000338
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1                                      'h0000033C
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2                                      'h00000340
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3                                      'h00000344
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4                                      'h00000348
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5                                      'h0000034C
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6                                      'h00000350
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7                                      'h00000354
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8                                      'h00000358
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0                                      'h0000035C
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1                                      'h00000360
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2                                      'h00000364
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3                                      'h00000368
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4                                      'h0000036C
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5                                      'h00000370
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6                                      'h00000374
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7                                      'h00000378
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8                                      'h0000037C
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000380
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                'h00000384
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                'h00000388
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                'h0000038C
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                'h00000390
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                'h00000394
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                'h00000398
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                'h0000039C
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                'h000003A0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                'h000003A4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                'h000003A8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                'h000003AC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                'h000003B0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                'h000003B4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                'h000003B8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                'h000003BC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                'h000003C0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                'h000003C4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                'h000003C8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                'h000003CC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                'h000003D0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                'h000003D4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                'h000003D8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                'h000003DC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                'h000003E0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                'h000003E4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                'h000003E8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                'h000003EC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                'h000003F0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                'h000003F4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                'h000003F8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                'h000003FC
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                'h00000400
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                'h00000404
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                'h00000408
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                'h0000040C
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000410
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                               'h00000414
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                               'h00000418
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                               'h0000041C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                               'h00000420
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                               'h00000424
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                               'h00000428
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                               'h0000042C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                               'h00000430
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000434
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                               'h00000438
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                               'h0000043C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                               'h00000440
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                               'h00000444
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                               'h00000448
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                               'h0000044C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                               'h00000450
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                               'h00000454
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000458
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                               'h0000045C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                               'h00000460
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                               'h00000464
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                               'h00000468
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                               'h0000046C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                               'h00000470
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                               'h00000474
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                               'h00000478
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h0000047C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                               'h00000480
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                               'h00000484
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                               'h00000488
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                               'h0000048C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                               'h00000490
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                               'h00000494
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                               'h00000498
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                               'h0000049C
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                            29:28
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                            25:24
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                            21:20
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                            17:16
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                            13:12
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                              9:8
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                              5:4
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                              1:0
`define CH0_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0                                      'h000004A0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1                                      'h000004A4
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2                                      'h000004A8
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3                                      'h000004AC
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4                                      'h000004B0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5                                      'h000004B4
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6                                      'h000004B8
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7                                      'h000004BC
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8                                      'h000004C0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0                                      'h000004C4
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1                                      'h000004C8
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2                                      'h000004CC
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3                                      'h000004D0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4                                      'h000004D4
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5                                      'h000004D8
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6                                      'h000004DC
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7                                      'h000004E0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8                                      'h000004E4
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0                                      'h000004E8
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1                                      'h000004EC
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2                                      'h000004F0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3                                      'h000004F4
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4                                      'h000004F8
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5                                      'h000004FC
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6                                      'h00000500
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7                                      'h00000504
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8                                      'h00000508
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0                                      'h0000050C
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1                                      'h00000510
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2                                      'h00000514
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3                                      'h00000518
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4                                      'h0000051C
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5                                      'h00000520
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6                                      'h00000524
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7                                      'h00000528
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8                                      'h0000052C
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000530
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                'h00000534
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                'h00000538
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                'h0000053C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                'h00000540
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                'h00000544
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                'h00000548
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                'h0000054C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                'h00000550
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000554
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                'h00000558
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                'h0000055C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                'h00000560
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                'h00000564
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                'h00000568
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                'h0000056C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                'h00000570
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                'h00000574
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000578
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                'h0000057C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                'h00000580
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                'h00000584
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                'h00000588
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                'h0000058C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                'h00000590
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                'h00000594
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                'h00000598
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                'h0000059C
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                'h000005A0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                'h000005A4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                'h000005A8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                'h000005AC
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                'h000005B0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                'h000005B4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                'h000005B8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                'h000005BC
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0                                      'h000005C0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1                                      'h000005C4
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2                                      'h000005C8
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3                                      'h000005CC
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4                                      'h000005D0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5                                      'h000005D4
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6                                      'h000005D8
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7                                      'h000005DC
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8                                      'h000005E0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0                                      'h000005E4
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1                                      'h000005E8
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2                                      'h000005EC
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3                                      'h000005F0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4                                      'h000005F4
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5                                      'h000005F8
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6                                      'h000005FC
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7                                      'h00000600
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8                                      'h00000604
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0                                      'h00000608
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1                                      'h0000060C
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2                                      'h00000610
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3                                      'h00000614
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4                                      'h00000618
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5                                      'h0000061C
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6                                      'h00000620
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7                                      'h00000624
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8                                      'h00000628
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0                                      'h0000062C
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1                                      'h00000630
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2                                      'h00000634
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3                                      'h00000638
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4                                      'h0000063C
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5                                      'h00000640
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6                                      'h00000644
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7                                      'h00000648
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8                                      'h0000064C
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000650
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                'h00000654
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                'h00000658
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                'h0000065C
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                'h00000660
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                'h00000664
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                'h00000668
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                'h0000066C
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                'h00000670
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000674
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                'h00000678
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                'h0000067C
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                'h00000680
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                'h00000684
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                'h00000688
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                'h0000068C
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                'h00000690
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                'h00000694
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000698
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                'h0000069C
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                'h000006A0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                'h000006A4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                'h000006A8
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                'h000006AC
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                'h000006B0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                'h000006B4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                'h000006B8
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                'h000006BC
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                'h000006C0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                'h000006C4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                'h000006C8
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                'h000006CC
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                'h000006D0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                'h000006D4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                'h000006D8
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                'h000006DC
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                               4
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                               0
`define CH0_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                     'h000006E0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                     'h000006E4
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                     'h000006E8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                     'h000006EC
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                     'h000006F0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                     'h000006F4
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                     'h000006F8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                     'h000006FC
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                     'h00000700
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                     'h00000704
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                     'h00000708
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                     'h0000070C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                     'h00000710
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                     'h00000714
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                     'h00000718
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                     'h0000071C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                     'h00000720
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                     'h00000724
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                     'h00000728
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                     'h0000072C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                     'h00000730
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                     'h00000734
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                     'h00000738
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                     'h0000073C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                     'h00000740
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                     'h00000744
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                     'h00000748
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                     'h0000074C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                     'h00000750
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                     'h00000754
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                     'h00000758
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                     'h0000075C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                     'h00000760
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                     'h00000764
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                     'h00000768
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                     'h0000076C
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                      7:6
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                          8
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                             32'h00000100

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0                                          'h00000770
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_0___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1                                          'h00000774
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_1___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2                                          'h00000778
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_2___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3                                          'h0000077C
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_3___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4                                          'h00000780
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_4___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5                                          'h00000784
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_5___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6                                          'h00000788
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_6___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7                                          'h0000078C
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_7___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8                                          'h00000790
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M0_CFG_8___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0                                          'h00000794
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_0___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1                                          'h00000798
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_1___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2                                          'h0000079C
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_2___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3                                          'h000007A0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_3___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4                                          'h000007A4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_4___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5                                          'h000007A8
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_5___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6                                          'h000007AC
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_6___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7                                          'h000007B0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_7___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8                                          'h000007B4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                        8:6
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                           5
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                       11:9
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                        4
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                         3
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                       2:0
`define CH0_DQ0_SWI_DQ_TX_IO_M1_CFG_8___POR                                  32'h00000040

`define CH0_DQ0_SWI_DQS_RX_M0_CFG                                              'h000007B8
`define CH0_DQ0_SWI_DQS_RX_M0_CFG__WCK_MODE                                             8
`define CH0_DQ0_SWI_DQS_RX_M0_CFG__RGB_MODE                                           2:0
`define CH0_DQ0_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                   13:12
`define CH0_DQ0_SWI_DQS_RX_M0_CFG__FGB_MODE                                           7:4
`define CH0_DQ0_SWI_DQS_RX_M0_CFG___POR                                      32'h00000074

`define CH0_DQ0_SWI_DQS_RX_M1_CFG                                              'h000007BC
`define CH0_DQ0_SWI_DQS_RX_M1_CFG__WCK_MODE                                             8
`define CH0_DQ0_SWI_DQS_RX_M1_CFG__RGB_MODE                                           2:0
`define CH0_DQ0_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                   13:12
`define CH0_DQ0_SWI_DQS_RX_M1_CFG__FGB_MODE                                           7:4
`define CH0_DQ0_SWI_DQS_RX_M1_CFG___POR                                      32'h00000074

`define CH0_DQ0_SWI_DQS_RX_BSCAN_STA                                           'h000007C0
`define CH0_DQ0_SWI_DQS_RX_BSCAN_STA__VAL                                             3:0
`define CH0_DQ0_SWI_DQS_RX_BSCAN_STA___POR                                   32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                  'h000007C4
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                   7:6
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                       8
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                               5:0
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                          32'h00000100

`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                  'h000007C8
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                   7:6
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                       8
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                               5:0
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                          32'h00000100

`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                  'h000007CC
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                   7:6
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                       8
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                               5:0
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                          32'h00000100

`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                  'h000007D0
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                   7:6
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                       8
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                               5:0
`define CH0_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                          32'h00000100

`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG                                    'h000007D4
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG                                    'h000007D8
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG                                    'h000007DC
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG                                    'h000007E0
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                    'h000007E4
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                    'h000007E8
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                    'h000007EC
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                    'h000007F0
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                 'h000007F4
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                 'h000007F8
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                 'h000007FC
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                 'h00000800
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                 'h00000804
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                 'h00000808
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                 'h0000080C
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                 'h00000810
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                13:10
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                  9:6
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                     14
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                  5:0
`define CH0_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                         32'h00000040

`define CH0_DQ0_SWI_DQS_RX_PI_STA                                              'h00000814
`define CH0_DQ0_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                         0
`define CH0_DQ0_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                         1
`define CH0_DQ0_SWI_DQS_RX_PI_STA___POR                                      32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0                                      'h00000818
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1                                      'h0000081C
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0                                      'h00000820
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1                                      'h00000824
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0                                      'h00000828
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1                                      'h0000082C
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0                                      'h00000830
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1                                      'h00000834
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                    'h00000838
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                    23
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                   22
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                  21
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                  18:16
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                        20
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                 19
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                  7:4
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                  3:0
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                15:12
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                 11:8
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                            32'h004A7777

`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                    'h0000083C
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                    23
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                   22
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                  21
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                  18:16
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                        20
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                 19
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                  7:4
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                  3:0
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                15:12
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                 11:8
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                            32'h004A7777

`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                    'h00000840
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                    23
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                   22
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                  21
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                  18:16
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                        20
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                 19
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                  7:4
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                  3:0
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                15:12
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                 11:8
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                            32'h004A7777

`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                    'h00000844
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                    23
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                   22
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                  21
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                  18:16
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                        20
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                 19
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                  7:4
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                  3:0
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                15:12
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                 11:8
`define CH0_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                            32'h004A7777

`define CH0_DQ0_SWI_DQS_RX_IO_STA                                              'h00000848
`define CH0_DQ0_SWI_DQS_RX_IO_STA__CORE_IG                                           31:0
`define CH0_DQ0_SWI_DQS_RX_IO_STA___POR                                      32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0                                      'h0000084C
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1                                      'h00000850
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0                                      'h00000854
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1                                      'h00000858
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0                                      'h0000085C
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1                                      'h00000860
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0                                      'h00000864
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1                                      'h00000868
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG                                          'h0000086C
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                           4
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                    2
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                     0
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                    3
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                     1
`define CH0_DQ0_SWI_DQS_RX_SA_CMN_CFG___POR                                  32'h00000005

`define CH0_DQ0_SWI_DQS_TX_M0_CFG                                              'h00000870
`define CH0_DQ0_SWI_DQS_TX_M0_CFG__WGB_MODE                                           7:4
`define CH0_DQ0_SWI_DQS_TX_M0_CFG__TGB_MODE                                           2:0
`define CH0_DQ0_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                       9:8
`define CH0_DQ0_SWI_DQS_TX_M0_CFG___POR                                      32'h00000087

`define CH0_DQ0_SWI_DQS_TX_M1_CFG                                              'h00000874
`define CH0_DQ0_SWI_DQS_TX_M1_CFG__WGB_MODE                                           7:4
`define CH0_DQ0_SWI_DQS_TX_M1_CFG__TGB_MODE                                           2:0
`define CH0_DQ0_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                       9:8
`define CH0_DQ0_SWI_DQS_TX_M1_CFG___POR                                      32'h00000087

`define CH0_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG                                      'h00000878
`define CH0_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                           1
`define CH0_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                           0
`define CH0_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                              32'h00000000

`define CH0_DQ0_SWI_DQS_TX_BSCAN_CFG                                           'h0000087C
`define CH0_DQ0_SWI_DQS_TX_BSCAN_CFG__VAL                                             3:0
`define CH0_DQ0_SWI_DQS_TX_BSCAN_CFG___POR                                   32'h00000000

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                 'h00000880
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1                                 'h00000884
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2                                 'h00000888
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3                                 'h0000088C
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4                                 'h00000890
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5                                 'h00000894
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6                                 'h00000898
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7                                 'h0000089C
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8                                 'h000008A0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                 'h000008A4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1                                 'h000008A8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2                                 'h000008AC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3                                 'h000008B0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4                                 'h000008B4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5                                 'h000008B8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6                                 'h000008BC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7                                 'h000008C0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8                                 'h000008C4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                           5:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8___POR                         32'h00000001

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                 'h000008C8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1                                 'h000008CC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2                                 'h000008D0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3                                 'h000008D4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4                                 'h000008D8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5                                 'h000008DC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6                                 'h000008E0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7                                 'h000008E4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8                                 'h000008E8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                 'h000008EC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1                                 'h000008F0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2                                 'h000008F4
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3                                 'h000008F8
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4                                 'h000008FC
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5                                 'h00000900
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6                                 'h00000904
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7                                 'h00000908
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8                                 'h0000090C
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                           6:0
`define CH0_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8___POR                         32'h00000002

`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                    'h00000910
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                    'h00000914
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                    'h00000918
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                    'h0000091C
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                  'h00000920
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                  'h00000924
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                  'h00000928
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                  'h0000092C
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                  'h00000930
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                  'h00000934
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                  'h00000938
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                  'h0000093C
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                  'h00000940
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                  'h00000944
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                  'h00000948
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                  'h0000094C
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                  'h00000950
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                  'h00000954
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                  'h00000958
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                  'h0000095C
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                      14
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG                                     'h00000960
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                         14
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG                                     'h00000964
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                         14
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG                                     'h00000968
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                         14
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG                                     'h0000096C
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                    13:10
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                      9:6
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                         14
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                      5:0
`define CH0_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                             32'h00000040

`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                    'h00000970
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                    'h00000974
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                    'h00000978
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                    'h0000097C
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                    'h00000980
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                    'h00000984
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                    'h00000988
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                    'h0000098C
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                     5:0
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ0_SWI_DQS_TX_RT_M0_R0_CFG                                        'h00000990
`define CH0_DQ0_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                      8:0
`define CH0_DQ0_SWI_DQS_TX_RT_M0_R0_CFG___POR                                32'h00000000

`define CH0_DQ0_SWI_DQS_TX_RT_M0_R1_CFG                                        'h00000994
`define CH0_DQ0_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                      8:0
`define CH0_DQ0_SWI_DQS_TX_RT_M0_R1_CFG___POR                                32'h00000000

`define CH0_DQ0_SWI_DQS_TX_RT_M1_R0_CFG                                        'h00000998
`define CH0_DQ0_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                      8:0
`define CH0_DQ0_SWI_DQS_TX_RT_M1_R0_CFG___POR                                32'h00000000

`define CH0_DQ0_SWI_DQS_TX_RT_M1_R1_CFG                                        'h0000099C
`define CH0_DQ0_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                      8:0
`define CH0_DQ0_SWI_DQS_TX_RT_M1_R1_CFG___POR                                32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0                                     'h000009A0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1                                     'h000009A4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2                                     'h000009A8
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3                                     'h000009AC
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4                                     'h000009B0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5                                     'h000009B4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6                                     'h000009B8
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7                                     'h000009BC
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8                                     'h000009C0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0                                     'h000009C4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1                                     'h000009C8
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2                                     'h000009CC
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3                                     'h000009D0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4                                     'h000009D4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5                                     'h000009D8
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6                                     'h000009DC
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7                                     'h000009E0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8                                     'h000009E4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0                                     'h000009E8
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1                                     'h000009EC
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2                                     'h000009F0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3                                     'h000009F4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4                                     'h000009F8
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5                                     'h000009FC
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6                                     'h00000A00
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7                                     'h00000A04
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8                                     'h00000A08
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0                                     'h00000A0C
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1                                     'h00000A10
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2                                     'h00000A14
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3                                     'h00000A18
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4                                     'h00000A1C
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5                                     'h00000A20
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6                                     'h00000A24
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7                                     'h00000A28
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8                                     'h00000A2C
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                               'h00000A30
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1                               'h00000A34
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2                               'h00000A38
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3                               'h00000A3C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4                               'h00000A40
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5                               'h00000A44
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6                               'h00000A48
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7                               'h00000A4C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8                               'h00000A50
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                               'h00000A54
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1                               'h00000A58
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2                               'h00000A5C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3                               'h00000A60
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4                               'h00000A64
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5                               'h00000A68
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6                               'h00000A6C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7                               'h00000A70
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8                               'h00000A74
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                               'h00000A78
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1                               'h00000A7C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2                               'h00000A80
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3                               'h00000A84
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4                               'h00000A88
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5                               'h00000A8C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6                               'h00000A90
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7                               'h00000A94
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8                               'h00000A98
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                               'h00000A9C
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1                               'h00000AA0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2                               'h00000AA4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3                               'h00000AA8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4                               'h00000AAC
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5                               'h00000AB0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6                               'h00000AB4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7                               'h00000AB8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8                               'h00000ABC
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                              'h00000AC0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1                              'h00000AC4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2                              'h00000AC8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3                              'h00000ACC
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4                              'h00000AD0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5                              'h00000AD4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6                              'h00000AD8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7                              'h00000ADC
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8                              'h00000AE0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                              'h00000AE4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1                              'h00000AE8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2                              'h00000AEC
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3                              'h00000AF0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4                              'h00000AF4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5                              'h00000AF8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6                              'h00000AFC
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7                              'h00000B00
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8                              'h00000B04
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                              'h00000B08
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1                              'h00000B0C
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2                              'h00000B10
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3                              'h00000B14
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4                              'h00000B18
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5                              'h00000B1C
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6                              'h00000B20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7                              'h00000B24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8                              'h00000B28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                              'h00000B2C
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1                              'h00000B30
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2                              'h00000B34
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3                              'h00000B38
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4                              'h00000B3C
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5                              'h00000B40
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6                              'h00000B44
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7                              'h00000B48
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8                              'h00000B4C
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                           29:28
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                           25:24
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                           21:20
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                           17:16
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                           13:12
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                             9:8
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                             5:4
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                             1:0
`define CH0_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                      32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0                                     'h00000B50
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1                                     'h00000B54
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2                                     'h00000B58
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3                                     'h00000B5C
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4                                     'h00000B60
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5                                     'h00000B64
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6                                     'h00000B68
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7                                     'h00000B6C
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8                                     'h00000B70
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0                                     'h00000B74
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1                                     'h00000B78
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2                                     'h00000B7C
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3                                     'h00000B80
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4                                     'h00000B84
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5                                     'h00000B88
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6                                     'h00000B8C
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7                                     'h00000B90
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8                                     'h00000B94
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0                                     'h00000B98
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1                                     'h00000B9C
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2                                     'h00000BA0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3                                     'h00000BA4
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4                                     'h00000BA8
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5                                     'h00000BAC
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6                                     'h00000BB0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7                                     'h00000BB4
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8                                     'h00000BB8
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0                                     'h00000BBC
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1                                     'h00000BC0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2                                     'h00000BC4
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3                                     'h00000BC8
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4                                     'h00000BCC
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5                                     'h00000BD0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6                                     'h00000BD4
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7                                     'h00000BD8
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8                                     'h00000BDC
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                               'h00000BE0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1                               'h00000BE4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2                               'h00000BE8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3                               'h00000BEC
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4                               'h00000BF0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5                               'h00000BF4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6                               'h00000BF8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7                               'h00000BFC
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8                               'h00000C00
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                               'h00000C04
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1                               'h00000C08
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2                               'h00000C0C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3                               'h00000C10
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4                               'h00000C14
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5                               'h00000C18
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6                               'h00000C1C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7                               'h00000C20
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8                               'h00000C24
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                               'h00000C28
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1                               'h00000C2C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2                               'h00000C30
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3                               'h00000C34
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4                               'h00000C38
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5                               'h00000C3C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6                               'h00000C40
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7                               'h00000C44
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8                               'h00000C48
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                               'h00000C4C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1                               'h00000C50
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2                               'h00000C54
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3                               'h00000C58
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4                               'h00000C5C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5                               'h00000C60
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6                               'h00000C64
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7                               'h00000C68
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8                               'h00000C6C
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0                                     'h00000C70
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1                                     'h00000C74
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2                                     'h00000C78
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3                                     'h00000C7C
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4                                     'h00000C80
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5                                     'h00000C84
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6                                     'h00000C88
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7                                     'h00000C8C
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8                                     'h00000C90
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0                                     'h00000C94
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1                                     'h00000C98
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2                                     'h00000C9C
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3                                     'h00000CA0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4                                     'h00000CA4
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5                                     'h00000CA8
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6                                     'h00000CAC
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7                                     'h00000CB0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8                                     'h00000CB4
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0                                     'h00000CB8
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1                                     'h00000CBC
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2                                     'h00000CC0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3                                     'h00000CC4
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4                                     'h00000CC8
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5                                     'h00000CCC
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6                                     'h00000CD0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7                                     'h00000CD4
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8                                     'h00000CD8
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0                                     'h00000CDC
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1                                     'h00000CE0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2                                     'h00000CE4
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3                                     'h00000CE8
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4                                     'h00000CEC
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5                                     'h00000CF0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6                                     'h00000CF4
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7                                     'h00000CF8
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8                                     'h00000CFC
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                               'h00000D00
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1                               'h00000D04
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2                               'h00000D08
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3                               'h00000D0C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4                               'h00000D10
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5                               'h00000D14
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6                               'h00000D18
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7                               'h00000D1C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8                               'h00000D20
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                               'h00000D24
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1                               'h00000D28
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2                               'h00000D2C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3                               'h00000D30
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4                               'h00000D34
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5                               'h00000D38
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6                               'h00000D3C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7                               'h00000D40
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8                               'h00000D44
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                               'h00000D48
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1                               'h00000D4C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2                               'h00000D50
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3                               'h00000D54
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4                               'h00000D58
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5                               'h00000D5C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6                               'h00000D60
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7                               'h00000D64
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8                               'h00000D68
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                               'h00000D6C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1                               'h00000D70
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2                               'h00000D74
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3                               'h00000D78
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4                               'h00000D7C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5                               'h00000D80
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6                               'h00000D84
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7                               'h00000D88
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8                               'h00000D8C
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              4
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              0
`define CH0_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                    'h00000D90
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1                                    'h00000D94
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                    'h00000D98
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1                                    'h00000D9C
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                    'h00000DA0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1                                    'h00000DA4
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                    'h00000DA8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1                                    'h00000DAC
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__GEAR                                     7:6
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__EN                                         8
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1___POR                            32'h00000100

`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0                                         'h00000DB0
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                       8:6
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                          5
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                      11:9
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                      4
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                      3
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                      2:0
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_0___POR                                 32'h00000041

`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1                                         'h00000DB4
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__TX_IMPD                                       8:6
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__SW_OVR                                          5
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__RX_IMPD                                      11:9
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_T                                      4
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_C                                      3
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_SEL                                      2:0
`define CH0_DQ0_SWI_DQS_TX_IO_M0_CFG_1___POR                                 32'h00000041

`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0                                         'h00000DB8
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                       8:6
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                          5
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                      11:9
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                      4
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                      3
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                      2:0
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_0___POR                                 32'h00000041

`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1                                         'h00000DBC
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__TX_IMPD                                       8:6
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__SW_OVR                                          5
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__RX_IMPD                                      11:9
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_T                                      4
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_C                                      3
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_SEL                                      2:0
`define CH0_DQ0_SWI_DQS_TX_IO_M1_CFG_1___POR                                 32'h00000041

`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                    'h00000DC0
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                   13
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                    10:5
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                     4:0
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                   12
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                     11
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                            32'h00000001

`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                    'h00000DC4
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                   13
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                    10:5
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                     4:0
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                   12
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                     11
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                            32'h00000001

`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                    'h00000DC8
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                   13
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                    10:5
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                     4:0
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                   12
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                     11
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                            32'h00000001

`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                    'h00000DCC
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                   13
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                    10:5
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                     4:0
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                   12
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                     11
`define CH0_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                            32'h00000001

`define CH0_DQ1_SWI_TOP_CFG                                                    'h00000000
`define CH0_DQ1_SWI_TOP_CFG__WCS_SW_OVR_VAL                                             1
`define CH0_DQ1_SWI_TOP_CFG__WCS_SW_OVR                                                 0
`define CH0_DQ1_SWI_TOP_CFG__TRAINING_MODE                                              9
`define CH0_DQ1_SWI_TOP_CFG__RCS_SW_OVR_VAL                                             3
`define CH0_DQ1_SWI_TOP_CFG__RCS_SW_OVR                                                 2
`define CH0_DQ1_SWI_TOP_CFG__FIFO_CLR                                                   8
`define CH0_DQ1_SWI_TOP_CFG___POR                                            32'h00000000

`define CH0_DQ1_SWI_TOP_STA                                                    'h00000004
`define CH0_DQ1_SWI_TOP_STA__WCS                                                        0
`define CH0_DQ1_SWI_TOP_STA__RCS                                                        1
`define CH0_DQ1_SWI_TOP_STA___POR                                            32'h00000000

`define CH0_DQ1_SWI_DQ_RX_BSCAN_STA                                            'h00000008
`define CH0_DQ1_SWI_DQ_RX_BSCAN_STA__VAL                                              8:0
`define CH0_DQ1_SWI_DQ_RX_BSCAN_STA___POR                                    32'h00000000

`define CH0_DQ1_SWI_DQ_RX_M0_CFG                                               'h0000000C
`define CH0_DQ1_SWI_DQ_RX_M0_CFG__RGB_MODE                                            2:0
`define CH0_DQ1_SWI_DQ_RX_M0_CFG__FGB_MODE                                            7:4
`define CH0_DQ1_SWI_DQ_RX_M0_CFG___POR                                       32'h00000074

`define CH0_DQ1_SWI_DQ_RX_M1_CFG                                               'h00000010
`define CH0_DQ1_SWI_DQ_RX_M1_CFG__RGB_MODE                                            2:0
`define CH0_DQ1_SWI_DQ_RX_M1_CFG__FGB_MODE                                            7:4
`define CH0_DQ1_SWI_DQ_RX_M1_CFG___POR                                       32'h00000074

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0                                       'h00000014
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1                                       'h00000018
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2                                       'h0000001C
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3                                       'h00000020
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4                                       'h00000024
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5                                       'h00000028
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6                                       'h0000002C
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7                                       'h00000030
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8                                       'h00000034
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0                                       'h00000038
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1                                       'h0000003C
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2                                       'h00000040
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3                                       'h00000044
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4                                       'h00000048
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5                                       'h0000004C
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6                                       'h00000050
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7                                       'h00000054
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8                                       'h00000058
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0                                       'h0000005C
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1                                       'h00000060
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2                                       'h00000064
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3                                       'h00000068
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4                                       'h0000006C
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5                                       'h00000070
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6                                       'h00000074
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7                                       'h00000078
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8                                       'h0000007C
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0                                       'h00000080
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1                                       'h00000084
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2                                       'h00000088
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3                                       'h0000008C
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4                                       'h00000090
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5                                       'h00000094
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6                                       'h00000098
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7                                       'h0000009C
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8                                       'h000000A0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                   7:0
`define CH0_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_IO_STA                                               'h000000A4
`define CH0_DQ1_SWI_DQ_RX_IO_STA__CORE_IG                                            31:0
`define CH0_DQ1_SWI_DQ_RX_IO_STA___POR                                       32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0                                       'h000000A8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1                                       'h000000AC
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2                                       'h000000B0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3                                       'h000000B4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4                                       'h000000B8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5                                       'h000000BC
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6                                       'h000000C0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7                                       'h000000C4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8                                       'h000000C8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0                                       'h000000CC
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1                                       'h000000D0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2                                       'h000000D4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3                                       'h000000D8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4                                       'h000000DC
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5                                       'h000000E0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6                                       'h000000E4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7                                       'h000000E8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8                                       'h000000EC
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0                                       'h000000F0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1                                       'h000000F4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2                                       'h000000F8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3                                       'h000000FC
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4                                       'h00000100
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5                                       'h00000104
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6                                       'h00000108
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7                                       'h0000010C
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8                                       'h00000110
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0                                       'h00000114
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1                                       'h00000118
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2                                       'h0000011C
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3                                       'h00000120
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4                                       'h00000124
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5                                       'h00000128
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6                                       'h0000012C
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7                                       'h00000130
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8                                       'h00000134
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                   17
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                  19
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                  18
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                    16
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                              15:12
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                               11:8
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH0_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                   'h00000138
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                   'h0000013C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                   'h00000140
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                   'h00000144
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                   'h00000148
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                   'h0000014C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                   'h00000150
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                   'h00000154
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                   'h00000158
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                   'h0000015C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                   'h00000160
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                   'h00000164
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                   'h00000168
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                   'h0000016C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                   'h00000170
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                   'h00000174
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                   'h00000178
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                   'h0000017C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                   'h00000180
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                   'h00000184
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                   'h00000188
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                   'h0000018C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                   'h00000190
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                   'h00000194
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                   'h00000198
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                   'h0000019C
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                   'h000001A0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                   'h000001A4
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                   'h000001A8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                   'h000001AC
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                   'h000001B0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                   'h000001B4
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                   'h000001B8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                   'h000001BC
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                   'h000001C0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                   'h000001C4
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                 9:8
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                              25:24
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                              17:16
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                  1:0
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                               15:10
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                              31:26
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                              23:18
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                  7:2
`define CH0_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                           32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_0                                             'h000001C8
`define CH0_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_0___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_1                                             'h000001CC
`define CH0_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_1___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_2                                             'h000001D0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_2___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_3                                             'h000001D4
`define CH0_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_3___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_4                                             'h000001D8
`define CH0_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_4___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_5                                             'h000001DC
`define CH0_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_5___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_6                                             'h000001E0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_6___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_7                                             'h000001E4
`define CH0_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_7___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_RX_SA_STA_8                                             'h000001E8
`define CH0_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                           1
`define CH0_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                          3
`define CH0_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                          2
`define CH0_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                            0
`define CH0_DQ1_SWI_DQ_RX_SA_STA_8___POR                                     32'h00000000

`define CH0_DQ1_SWI_DQ_TX_BSCAN_CFG                                            'h000001EC
`define CH0_DQ1_SWI_DQ_TX_BSCAN_CFG__VAL                                              8:0
`define CH0_DQ1_SWI_DQ_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                  'h000001F0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                  'h000001F4
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                  'h000001F8
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                  'h000001FC
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                  'h00000200
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                  'h00000204
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                  'h00000208
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                  'h0000020C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                  'h00000210
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                  'h00000214
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                  'h00000218
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                  'h0000021C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                  'h00000220
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                  'h00000224
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                  'h00000228
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                  'h0000022C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                  'h00000230
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                  'h00000234
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                            5:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                          32'h00000001

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                  'h00000238
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                  'h0000023C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                  'h00000240
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                  'h00000244
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                  'h00000248
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                  'h0000024C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                  'h00000250
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                  'h00000254
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                  'h00000258
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                  'h0000025C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                  'h00000260
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                  'h00000264
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                  'h00000268
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                  'h0000026C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                  'h00000270
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                  'h00000274
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                  'h00000278
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                  'h0000027C
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                            6:0
`define CH0_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                          32'h00000002

`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                     'h00000280
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                     'h00000284
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                     'h00000288
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                     'h0000028C
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                   'h00000290
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                   'h00000294
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                   'h00000298
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                   'h0000029C
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                   'h000002A0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                   'h000002A4
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                   'h000002A8
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                   'h000002AC
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                   'h000002B0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                   'h000002B4
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                   'h000002B8
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                   'h000002BC
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                   'h000002C0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                   'h000002C4
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                   'h000002C8
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                   'h000002CC
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG                                      'h000002D0
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG                                      'h000002D4
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG                                      'h000002D8
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG                                      'h000002DC
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH0_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH0_DQ1_SWI_DQ_TX_RT_M0_R0_CFG                                         'h000002E0
`define CH0_DQ1_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       8:0
`define CH0_DQ1_SWI_DQ_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH0_DQ1_SWI_DQ_TX_RT_M0_R1_CFG                                         'h000002E4
`define CH0_DQ1_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       8:0
`define CH0_DQ1_SWI_DQ_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH0_DQ1_SWI_DQ_TX_RT_M1_R0_CFG                                         'h000002E8
`define CH0_DQ1_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       8:0
`define CH0_DQ1_SWI_DQ_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH0_DQ1_SWI_DQ_TX_RT_M1_R1_CFG                                         'h000002EC
`define CH0_DQ1_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       8:0
`define CH0_DQ1_SWI_DQ_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0                                      'h000002F0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1                                      'h000002F4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2                                      'h000002F8
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3                                      'h000002FC
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4                                      'h00000300
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5                                      'h00000304
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6                                      'h00000308
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7                                      'h0000030C
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8                                      'h00000310
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0                                      'h00000314
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1                                      'h00000318
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2                                      'h0000031C
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3                                      'h00000320
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4                                      'h00000324
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5                                      'h00000328
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6                                      'h0000032C
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7                                      'h00000330
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8                                      'h00000334
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0                                      'h00000338
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1                                      'h0000033C
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2                                      'h00000340
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3                                      'h00000344
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4                                      'h00000348
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5                                      'h0000034C
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6                                      'h00000350
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7                                      'h00000354
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8                                      'h00000358
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0                                      'h0000035C
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1                                      'h00000360
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2                                      'h00000364
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3                                      'h00000368
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4                                      'h0000036C
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5                                      'h00000370
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6                                      'h00000374
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7                                      'h00000378
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8                                      'h0000037C
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                   7
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                   6
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                   5
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                   4
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000380
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                'h00000384
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                'h00000388
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                'h0000038C
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                'h00000390
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                'h00000394
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                'h00000398
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                'h0000039C
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                'h000003A0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                'h000003A4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                'h000003A8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                'h000003AC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                'h000003B0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                'h000003B4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                'h000003B8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                'h000003BC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                'h000003C0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                'h000003C4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                'h000003C8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                'h000003CC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                'h000003D0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                'h000003D4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                'h000003D8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                'h000003DC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                'h000003E0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                'h000003E4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                'h000003E8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                'h000003EC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                'h000003F0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                'h000003F4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                'h000003F8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                'h000003FC
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                'h00000400
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                'h00000404
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                'h00000408
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                'h0000040C
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                           30:28
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                           26:24
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                           22:20
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                           18:16
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           14:12
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            10:8
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             6:4
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             2:0
`define CH0_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000410
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                               'h00000414
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                               'h00000418
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                               'h0000041C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                               'h00000420
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                               'h00000424
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                               'h00000428
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                               'h0000042C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                               'h00000430
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000434
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                               'h00000438
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                               'h0000043C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                               'h00000440
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                               'h00000444
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                               'h00000448
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                               'h0000044C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                               'h00000450
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                               'h00000454
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000458
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                               'h0000045C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                               'h00000460
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                               'h00000464
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                               'h00000468
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                               'h0000046C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                               'h00000470
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                               'h00000474
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                               'h00000478
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h0000047C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                               'h00000480
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                               'h00000484
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                               'h00000488
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                               'h0000048C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                               'h00000490
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                               'h00000494
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                               'h00000498
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                               'h0000049C
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                            29:28
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                            25:24
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                            21:20
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                            17:16
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                            13:12
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                              9:8
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                              5:4
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                              1:0
`define CH0_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0                                      'h000004A0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1                                      'h000004A4
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2                                      'h000004A8
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3                                      'h000004AC
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4                                      'h000004B0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5                                      'h000004B4
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6                                      'h000004B8
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7                                      'h000004BC
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8                                      'h000004C0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0                                      'h000004C4
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1                                      'h000004C8
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2                                      'h000004CC
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3                                      'h000004D0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4                                      'h000004D4
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5                                      'h000004D8
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6                                      'h000004DC
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7                                      'h000004E0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8                                      'h000004E4
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0                                      'h000004E8
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1                                      'h000004EC
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2                                      'h000004F0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3                                      'h000004F4
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4                                      'h000004F8
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5                                      'h000004FC
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6                                      'h00000500
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7                                      'h00000504
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8                                      'h00000508
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0                                      'h0000050C
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1                                      'h00000510
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2                                      'h00000514
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3                                      'h00000518
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4                                      'h0000051C
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5                                      'h00000520
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6                                      'h00000524
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7                                      'h00000528
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8                                      'h0000052C
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000530
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                'h00000534
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                'h00000538
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                'h0000053C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                'h00000540
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                'h00000544
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                'h00000548
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                'h0000054C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                'h00000550
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000554
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                'h00000558
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                'h0000055C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                'h00000560
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                'h00000564
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                'h00000568
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                'h0000056C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                'h00000570
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                'h00000574
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000578
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                'h0000057C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                'h00000580
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                'h00000584
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                'h00000588
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                'h0000058C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                'h00000590
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                'h00000594
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                'h00000598
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                'h0000059C
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                'h000005A0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                'h000005A4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                'h000005A8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                'h000005AC
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                'h000005B0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                'h000005B4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                'h000005B8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                'h000005BC
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           13:12
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             9:8
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             5:4
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             1:0
`define CH0_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0                                      'h000005C0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1                                      'h000005C4
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2                                      'h000005C8
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3                                      'h000005CC
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4                                      'h000005D0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5                                      'h000005D4
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6                                      'h000005D8
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7                                      'h000005DC
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8                                      'h000005E0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0                                      'h000005E4
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1                                      'h000005E8
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2                                      'h000005EC
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3                                      'h000005F0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4                                      'h000005F4
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5                                      'h000005F8
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6                                      'h000005FC
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7                                      'h00000600
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8                                      'h00000604
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0                                      'h00000608
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1                                      'h0000060C
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2                                      'h00000610
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3                                      'h00000614
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4                                      'h00000618
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5                                      'h0000061C
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6                                      'h00000620
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7                                      'h00000624
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8                                      'h00000628
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0                                      'h0000062C
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1                                      'h00000630
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2                                      'h00000634
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3                                      'h00000638
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4                                      'h0000063C
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5                                      'h00000640
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6                                      'h00000644
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7                                      'h00000648
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8                                      'h0000064C
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH0_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000650
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                'h00000654
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                'h00000658
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                'h0000065C
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                'h00000660
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                'h00000664
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                'h00000668
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                'h0000066C
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                'h00000670
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000674
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                'h00000678
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                'h0000067C
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                'h00000680
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                'h00000684
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                'h00000688
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                'h0000068C
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                'h00000690
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                'h00000694
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000698
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                'h0000069C
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                'h000006A0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                'h000006A4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                'h000006A8
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                'h000006AC
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                'h000006B0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                'h000006B4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                'h000006B8
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                'h000006BC
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                'h000006C0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                'h000006C4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                'h000006C8
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                'h000006CC
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                'h000006D0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                'h000006D4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                'h000006D8
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                'h000006DC
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                               4
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                               0
`define CH0_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                     'h000006E0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                     'h000006E4
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                     'h000006E8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                     'h000006EC
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                     'h000006F0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                     'h000006F4
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                     'h000006F8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                     'h000006FC
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                     'h00000700
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                     'h00000704
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                     'h00000708
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                     'h0000070C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                     'h00000710
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                     'h00000714
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                     'h00000718
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                     'h0000071C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                     'h00000720
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                     'h00000724
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                     'h00000728
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                     'h0000072C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                     'h00000730
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                     'h00000734
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                     'h00000738
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                     'h0000073C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                     'h00000740
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                     'h00000744
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                     'h00000748
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                     'h0000074C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                     'h00000750
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                     'h00000754
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                     'h00000758
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                     'h0000075C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                     'h00000760
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                     'h00000764
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                     'h00000768
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                     'h0000076C
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                      7:6
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                          8
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                  5:0
`define CH0_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                             32'h00000100

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0                                          'h00000770
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_0___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1                                          'h00000774
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_1___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2                                          'h00000778
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_2___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3                                          'h0000077C
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_3___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4                                          'h00000780
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_4___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5                                          'h00000784
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_5___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6                                          'h00000788
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_6___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7                                          'h0000078C
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_7___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8                                          'h00000790
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M0_CFG_8___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0                                          'h00000794
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_0___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1                                          'h00000798
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_1___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2                                          'h0000079C
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_2___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3                                          'h000007A0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_3___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4                                          'h000007A4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_4___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5                                          'h000007A8
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_5___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6                                          'h000007AC
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_6___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7                                          'h000007B0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_7___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8                                          'h000007B4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                        8:6
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                           5
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                       11:9
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                        4
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                         3
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                       2:0
`define CH0_DQ1_SWI_DQ_TX_IO_M1_CFG_8___POR                                  32'h00000040

`define CH0_DQ1_SWI_DQS_RX_M0_CFG                                              'h000007B8
`define CH0_DQ1_SWI_DQS_RX_M0_CFG__WCK_MODE                                             8
`define CH0_DQ1_SWI_DQS_RX_M0_CFG__RGB_MODE                                           2:0
`define CH0_DQ1_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                   13:12
`define CH0_DQ1_SWI_DQS_RX_M0_CFG__FGB_MODE                                           7:4
`define CH0_DQ1_SWI_DQS_RX_M0_CFG___POR                                      32'h00000074

`define CH0_DQ1_SWI_DQS_RX_M1_CFG                                              'h000007BC
`define CH0_DQ1_SWI_DQS_RX_M1_CFG__WCK_MODE                                             8
`define CH0_DQ1_SWI_DQS_RX_M1_CFG__RGB_MODE                                           2:0
`define CH0_DQ1_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                   13:12
`define CH0_DQ1_SWI_DQS_RX_M1_CFG__FGB_MODE                                           7:4
`define CH0_DQ1_SWI_DQS_RX_M1_CFG___POR                                      32'h00000074

`define CH0_DQ1_SWI_DQS_RX_BSCAN_STA                                           'h000007C0
`define CH0_DQ1_SWI_DQS_RX_BSCAN_STA__VAL                                             3:0
`define CH0_DQ1_SWI_DQS_RX_BSCAN_STA___POR                                   32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                  'h000007C4
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                   7:6
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                       8
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                               5:0
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                          32'h00000100

`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                  'h000007C8
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                   7:6
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                       8
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                               5:0
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                          32'h00000100

`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                  'h000007CC
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                   7:6
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                       8
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                               5:0
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                          32'h00000100

`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                  'h000007D0
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                   7:6
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                       8
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                               5:0
`define CH0_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                          32'h00000100

`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG                                    'h000007D4
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG                                    'h000007D8
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG                                    'h000007DC
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG                                    'h000007E0
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                    'h000007E4
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                    'h000007E8
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                    'h000007EC
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                    'h000007F0
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                 'h000007F4
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                 'h000007F8
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                 'h000007FC
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                 'h00000800
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                 'h00000804
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                 'h00000808
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                 'h0000080C
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                 'h00000810
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                13:10
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                  9:6
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                     14
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                  5:0
`define CH0_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                         32'h00000040

`define CH0_DQ1_SWI_DQS_RX_PI_STA                                              'h00000814
`define CH0_DQ1_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                         0
`define CH0_DQ1_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                         1
`define CH0_DQ1_SWI_DQS_RX_PI_STA___POR                                      32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0                                      'h00000818
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1                                      'h0000081C
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0                                      'h00000820
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1                                      'h00000824
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0                                      'h00000828
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1                                      'h0000082C
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0                                      'h00000830
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1                                      'h00000834
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH0_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                    'h00000838
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                    23
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                   22
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                  21
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                  18:16
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                        20
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                 19
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                  7:4
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                  3:0
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                15:12
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                 11:8
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                            32'h004A7777

`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                    'h0000083C
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                    23
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                   22
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                  21
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                  18:16
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                        20
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                 19
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                  7:4
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                  3:0
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                15:12
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                 11:8
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                            32'h004A7777

`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                    'h00000840
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                    23
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                   22
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                  21
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                  18:16
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                        20
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                 19
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                  7:4
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                  3:0
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                15:12
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                 11:8
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                            32'h004A7777

`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                    'h00000844
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                    23
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                   22
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                  21
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                  18:16
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                        20
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                 19
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                  7:4
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                  3:0
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                15:12
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                 11:8
`define CH0_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                            32'h004A7777

`define CH0_DQ1_SWI_DQS_RX_IO_STA                                              'h00000848
`define CH0_DQ1_SWI_DQS_RX_IO_STA__CORE_IG                                           31:0
`define CH0_DQ1_SWI_DQS_RX_IO_STA___POR                                      32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0                                      'h0000084C
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1                                      'h00000850
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0                                      'h00000854
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1                                      'h00000858
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0                                      'h0000085C
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1                                      'h00000860
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0                                      'h00000864
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1                                      'h00000868
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                  17
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                 19
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                 18
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                   16
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                7:4
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_270                             15:12
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_180                              11:8
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH0_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG                                          'h0000086C
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                           4
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                    2
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                     0
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                    3
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                     1
`define CH0_DQ1_SWI_DQS_RX_SA_CMN_CFG___POR                                  32'h00000005

`define CH0_DQ1_SWI_DQS_TX_M0_CFG                                              'h00000870
`define CH0_DQ1_SWI_DQS_TX_M0_CFG__WGB_MODE                                           7:4
`define CH0_DQ1_SWI_DQS_TX_M0_CFG__TGB_MODE                                           2:0
`define CH0_DQ1_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                       9:8
`define CH0_DQ1_SWI_DQS_TX_M0_CFG___POR                                      32'h00000087

`define CH0_DQ1_SWI_DQS_TX_M1_CFG                                              'h00000874
`define CH0_DQ1_SWI_DQS_TX_M1_CFG__WGB_MODE                                           7:4
`define CH0_DQ1_SWI_DQS_TX_M1_CFG__TGB_MODE                                           2:0
`define CH0_DQ1_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                       9:8
`define CH0_DQ1_SWI_DQS_TX_M1_CFG___POR                                      32'h00000087

`define CH0_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG                                      'h00000878
`define CH0_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                           1
`define CH0_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                           0
`define CH0_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                              32'h00000000

`define CH0_DQ1_SWI_DQS_TX_BSCAN_CFG                                           'h0000087C
`define CH0_DQ1_SWI_DQS_TX_BSCAN_CFG__VAL                                             3:0
`define CH0_DQ1_SWI_DQS_TX_BSCAN_CFG___POR                                   32'h00000000

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                 'h00000880
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1                                 'h00000884
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2                                 'h00000888
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3                                 'h0000088C
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4                                 'h00000890
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5                                 'h00000894
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6                                 'h00000898
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7                                 'h0000089C
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8                                 'h000008A0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                 'h000008A4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1                                 'h000008A8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2                                 'h000008AC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3                                 'h000008B0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4                                 'h000008B4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5                                 'h000008B8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6                                 'h000008BC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7                                 'h000008C0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8                                 'h000008C4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                           5:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8___POR                         32'h00000001

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                 'h000008C8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1                                 'h000008CC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2                                 'h000008D0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3                                 'h000008D4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4                                 'h000008D8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5                                 'h000008DC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6                                 'h000008E0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7                                 'h000008E4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8                                 'h000008E8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                 'h000008EC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1                                 'h000008F0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2                                 'h000008F4
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3                                 'h000008F8
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4                                 'h000008FC
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5                                 'h00000900
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6                                 'h00000904
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7                                 'h00000908
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8                                 'h0000090C
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                           6:0
`define CH0_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8___POR                         32'h00000002

`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                    'h00000910
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                    'h00000914
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                    'h00000918
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                    'h0000091C
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                     5:0
`define CH0_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                  'h00000920
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                  'h00000924
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                  'h00000928
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                  'h0000092C
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                  'h00000930
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                  'h00000934
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                  'h00000938
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                  'h0000093C
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                  'h00000940
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                  'h00000944
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                  'h00000948
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                  'h0000094C
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                  'h00000950
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                  'h00000954
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                  'h00000958
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                  'h0000095C
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                      14
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH0_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG                                     'h00000960
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                         14
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG                                     'h00000964
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                         14
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG                                     'h00000968
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                         14
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG                                     'h0000096C
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                    13:10
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                      9:6
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                         14
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                      5:0
`define CH0_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                             32'h00000040

`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                    'h00000970
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                    'h00000974
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                    'h00000978
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                    'h0000097C
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                    'h00000980
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                    'h00000984
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                    'h00000988
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                    'h0000098C
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                   13:10
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                     5:0
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                     9:6
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                        14
`define CH0_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                            32'h00000040

`define CH0_DQ1_SWI_DQS_TX_RT_M0_R0_CFG                                        'h00000990
`define CH0_DQ1_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                      8:0
`define CH0_DQ1_SWI_DQS_TX_RT_M0_R0_CFG___POR                                32'h00000000

`define CH0_DQ1_SWI_DQS_TX_RT_M0_R1_CFG                                        'h00000994
`define CH0_DQ1_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                      8:0
`define CH0_DQ1_SWI_DQS_TX_RT_M0_R1_CFG___POR                                32'h00000000

`define CH0_DQ1_SWI_DQS_TX_RT_M1_R0_CFG                                        'h00000998
`define CH0_DQ1_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                      8:0
`define CH0_DQ1_SWI_DQS_TX_RT_M1_R0_CFG___POR                                32'h00000000

`define CH0_DQ1_SWI_DQS_TX_RT_M1_R1_CFG                                        'h0000099C
`define CH0_DQ1_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                      8:0
`define CH0_DQ1_SWI_DQS_TX_RT_M1_R1_CFG___POR                                32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0                                     'h000009A0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1                                     'h000009A4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2                                     'h000009A8
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3                                     'h000009AC
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4                                     'h000009B0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5                                     'h000009B4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6                                     'h000009B8
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7                                     'h000009BC
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8                                     'h000009C0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0                                     'h000009C4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1                                     'h000009C8
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2                                     'h000009CC
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3                                     'h000009D0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4                                     'h000009D4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5                                     'h000009D8
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6                                     'h000009DC
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7                                     'h000009E0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8                                     'h000009E4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0                                     'h000009E8
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1                                     'h000009EC
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2                                     'h000009F0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3                                     'h000009F4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4                                     'h000009F8
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5                                     'h000009FC
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6                                     'h00000A00
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7                                     'h00000A04
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8                                     'h00000A08
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0                                     'h00000A0C
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1                                     'h00000A10
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2                                     'h00000A14
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3                                     'h00000A18
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4                                     'h00000A1C
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5                                     'h00000A20
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6                                     'h00000A24
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7                                     'h00000A28
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8                                     'h00000A2C
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                  7
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                  6
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                  5
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                  4
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                               'h00000A30
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1                               'h00000A34
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2                               'h00000A38
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3                               'h00000A3C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4                               'h00000A40
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5                               'h00000A44
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6                               'h00000A48
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7                               'h00000A4C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8                               'h00000A50
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                               'h00000A54
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1                               'h00000A58
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2                               'h00000A5C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3                               'h00000A60
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4                               'h00000A64
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5                               'h00000A68
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6                               'h00000A6C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7                               'h00000A70
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8                               'h00000A74
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                               'h00000A78
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1                               'h00000A7C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2                               'h00000A80
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3                               'h00000A84
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4                               'h00000A88
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5                               'h00000A8C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6                               'h00000A90
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7                               'h00000A94
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8                               'h00000A98
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                               'h00000A9C
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1                               'h00000AA0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2                               'h00000AA4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3                               'h00000AA8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4                               'h00000AAC
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5                               'h00000AB0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6                               'h00000AB4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7                               'h00000AB8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8                               'h00000ABC
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                          30:28
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                          26:24
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                          22:20
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                          18:16
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          14:12
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                           10:8
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            6:4
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            2:0
`define CH0_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                              'h00000AC0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1                              'h00000AC4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2                              'h00000AC8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3                              'h00000ACC
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4                              'h00000AD0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5                              'h00000AD4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6                              'h00000AD8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7                              'h00000ADC
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8                              'h00000AE0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                              'h00000AE4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1                              'h00000AE8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2                              'h00000AEC
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3                              'h00000AF0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4                              'h00000AF4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5                              'h00000AF8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6                              'h00000AFC
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7                              'h00000B00
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8                              'h00000B04
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                              'h00000B08
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1                              'h00000B0C
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2                              'h00000B10
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3                              'h00000B14
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4                              'h00000B18
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5                              'h00000B1C
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6                              'h00000B20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7                              'h00000B24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8                              'h00000B28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                              'h00000B2C
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1                              'h00000B30
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2                              'h00000B34
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3                              'h00000B38
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4                              'h00000B3C
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5                              'h00000B40
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6                              'h00000B44
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7                              'h00000B48
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8                              'h00000B4C
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                           29:28
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                           25:24
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                           21:20
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                           17:16
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                           13:12
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                             9:8
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                             5:4
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                             1:0
`define CH0_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                      32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0                                     'h00000B50
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1                                     'h00000B54
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2                                     'h00000B58
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3                                     'h00000B5C
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4                                     'h00000B60
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5                                     'h00000B64
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6                                     'h00000B68
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7                                     'h00000B6C
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8                                     'h00000B70
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0                                     'h00000B74
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1                                     'h00000B78
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2                                     'h00000B7C
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3                                     'h00000B80
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4                                     'h00000B84
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5                                     'h00000B88
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6                                     'h00000B8C
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7                                     'h00000B90
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8                                     'h00000B94
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0                                     'h00000B98
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1                                     'h00000B9C
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2                                     'h00000BA0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3                                     'h00000BA4
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4                                     'h00000BA8
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5                                     'h00000BAC
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6                                     'h00000BB0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7                                     'h00000BB4
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8                                     'h00000BB8
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0                                     'h00000BBC
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1                                     'h00000BC0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2                                     'h00000BC4
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3                                     'h00000BC8
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4                                     'h00000BCC
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5                                     'h00000BD0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6                                     'h00000BD4
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7                                     'h00000BD8
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8                                     'h00000BDC
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                               'h00000BE0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1                               'h00000BE4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2                               'h00000BE8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3                               'h00000BEC
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4                               'h00000BF0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5                               'h00000BF4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6                               'h00000BF8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7                               'h00000BFC
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8                               'h00000C00
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                               'h00000C04
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1                               'h00000C08
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2                               'h00000C0C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3                               'h00000C10
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4                               'h00000C14
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5                               'h00000C18
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6                               'h00000C1C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7                               'h00000C20
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8                               'h00000C24
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                               'h00000C28
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1                               'h00000C2C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2                               'h00000C30
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3                               'h00000C34
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4                               'h00000C38
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5                               'h00000C3C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6                               'h00000C40
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7                               'h00000C44
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8                               'h00000C48
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                               'h00000C4C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1                               'h00000C50
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2                               'h00000C54
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3                               'h00000C58
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4                               'h00000C5C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5                               'h00000C60
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6                               'h00000C64
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7                               'h00000C68
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8                               'h00000C6C
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          13:12
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            9:8
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            5:4
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            1:0
`define CH0_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0                                     'h00000C70
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1                                     'h00000C74
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2                                     'h00000C78
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3                                     'h00000C7C
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4                                     'h00000C80
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5                                     'h00000C84
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6                                     'h00000C88
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7                                     'h00000C8C
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8                                     'h00000C90
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0                                     'h00000C94
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1                                     'h00000C98
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2                                     'h00000C9C
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3                                     'h00000CA0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4                                     'h00000CA4
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5                                     'h00000CA8
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6                                     'h00000CAC
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7                                     'h00000CB0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8                                     'h00000CB4
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0                                     'h00000CB8
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1                                     'h00000CBC
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2                                     'h00000CC0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3                                     'h00000CC4
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4                                     'h00000CC8
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5                                     'h00000CCC
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6                                     'h00000CD0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7                                     'h00000CD4
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8                                     'h00000CD8
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0                                     'h00000CDC
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1                                     'h00000CE0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2                                     'h00000CE4
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3                                     'h00000CE8
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4                                     'h00000CEC
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5                                     'h00000CF0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6                                     'h00000CF4
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7                                     'h00000CF8
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8                                     'h00000CFC
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH0_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                               'h00000D00
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1                               'h00000D04
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2                               'h00000D08
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3                               'h00000D0C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4                               'h00000D10
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5                               'h00000D14
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6                               'h00000D18
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7                               'h00000D1C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8                               'h00000D20
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                               'h00000D24
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1                               'h00000D28
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2                               'h00000D2C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3                               'h00000D30
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4                               'h00000D34
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5                               'h00000D38
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6                               'h00000D3C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7                               'h00000D40
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8                               'h00000D44
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                               'h00000D48
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1                               'h00000D4C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2                               'h00000D50
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3                               'h00000D54
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4                               'h00000D58
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5                               'h00000D5C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6                               'h00000D60
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7                               'h00000D64
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8                               'h00000D68
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                               'h00000D6C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1                               'h00000D70
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2                               'h00000D74
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3                               'h00000D78
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4                               'h00000D7C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5                               'h00000D80
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6                               'h00000D84
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7                               'h00000D88
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8                               'h00000D8C
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              4
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              0
`define CH0_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                    'h00000D90
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1                                    'h00000D94
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                    'h00000D98
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1                                    'h00000D9C
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                    'h00000DA0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1                                    'h00000DA4
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                    'h00000DA8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1                                    'h00000DAC
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__GEAR                                     7:6
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__EN                                         8
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                 5:0
`define CH0_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1___POR                            32'h00000100

`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0                                         'h00000DB0
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                       8:6
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                          5
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                      11:9
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                      4
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                      3
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                      2:0
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_0___POR                                 32'h00000041

`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1                                         'h00000DB4
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__TX_IMPD                                       8:6
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__SW_OVR                                          5
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__RX_IMPD                                      11:9
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_T                                      4
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_C                                      3
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_SEL                                      2:0
`define CH0_DQ1_SWI_DQS_TX_IO_M0_CFG_1___POR                                 32'h00000041

`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0                                         'h00000DB8
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                       8:6
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                          5
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                      11:9
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                      4
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                      3
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                      2:0
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_0___POR                                 32'h00000041

`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1                                         'h00000DBC
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__TX_IMPD                                       8:6
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__SW_OVR                                          5
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__RX_IMPD                                      11:9
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_T                                      4
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_C                                      3
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_SEL                                      2:0
`define CH0_DQ1_SWI_DQS_TX_IO_M1_CFG_1___POR                                 32'h00000041

`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                    'h00000DC0
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                   13
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                    10:5
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                     4:0
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                   12
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                     11
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                            32'h00000001

`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                    'h00000DC4
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                   13
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                    10:5
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                     4:0
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                   12
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                     11
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                            32'h00000001

`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                    'h00000DC8
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                   13
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                    10:5
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                     4:0
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                   12
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                     11
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                            32'h00000001

`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                    'h00000DCC
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                   13
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                    10:5
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                     4:0
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                   12
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                     11
`define CH0_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                            32'h00000001

`define CH0_CA_SWI_TOP_CFG                                                     'h00000000
`define CH0_CA_SWI_TOP_CFG__WCS_SW_OVR_VAL                                              1
`define CH0_CA_SWI_TOP_CFG__WCS_SW_OVR                                                  0
`define CH0_CA_SWI_TOP_CFG__TRAINING_MODE                                               9
`define CH0_CA_SWI_TOP_CFG__RCS_SW_OVR_VAL                                              3
`define CH0_CA_SWI_TOP_CFG__RCS_SW_OVR                                                  2
`define CH0_CA_SWI_TOP_CFG__FIFO_CLR                                                    8
`define CH0_CA_SWI_TOP_CFG___POR                                             32'h00000000

`define CH0_CA_SWI_TOP_STA                                                     'h00000004
`define CH0_CA_SWI_TOP_STA__WCS                                                         0
`define CH0_CA_SWI_TOP_STA__RCS                                                         1
`define CH0_CA_SWI_TOP_STA___POR                                             32'h00000000

`define CH0_CA_SWI_DQ_RX_BSCAN_STA                                             'h00000008
`define CH0_CA_SWI_DQ_RX_BSCAN_STA__VAL                                              10:0
`define CH0_CA_SWI_DQ_RX_BSCAN_STA___POR                                     32'h00000000

`define CH0_CA_SWI_DQ_RX_M0_CFG                                                'h0000000C
`define CH0_CA_SWI_DQ_RX_M0_CFG__RGB_MODE                                             2:0
`define CH0_CA_SWI_DQ_RX_M0_CFG__FGB_MODE                                             7:4
`define CH0_CA_SWI_DQ_RX_M0_CFG___POR                                        32'h00000074

`define CH0_CA_SWI_DQ_RX_M1_CFG                                                'h00000010
`define CH0_CA_SWI_DQ_RX_M1_CFG__RGB_MODE                                             2:0
`define CH0_CA_SWI_DQ_RX_M1_CFG__FGB_MODE                                             7:4
`define CH0_CA_SWI_DQ_RX_M1_CFG___POR                                        32'h00000074

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_0                                        'h00000014
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_1                                        'h00000018
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_2                                        'h0000001C
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_3                                        'h00000020
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_4                                        'h00000024
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_5                                        'h00000028
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_6                                        'h0000002C
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_7                                        'h00000030
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_8                                        'h00000034
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_9                                        'h00000038
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_9__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_10                                       'h0000003C
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_10__RESERVED0                                   7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R0_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_0                                        'h00000040
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_1                                        'h00000044
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_2                                        'h00000048
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_3                                        'h0000004C
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_4                                        'h00000050
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_5                                        'h00000054
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_6                                        'h00000058
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_7                                        'h0000005C
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_8                                        'h00000060
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_9                                        'h00000064
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_9__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_10                                       'h00000068
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_10__RESERVED0                                   7:0
`define CH0_CA_SWI_DQ_RX_IO_M0_R1_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_0                                        'h0000006C
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_1                                        'h00000070
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_2                                        'h00000074
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_3                                        'h00000078
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_4                                        'h0000007C
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_5                                        'h00000080
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_6                                        'h00000084
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_7                                        'h00000088
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_8                                        'h0000008C
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_9                                        'h00000090
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_9__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_10                                       'h00000094
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_10__RESERVED0                                   7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R0_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_0                                        'h00000098
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_1                                        'h0000009C
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_2                                        'h000000A0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_3                                        'h000000A4
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_4                                        'h000000A8
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_5                                        'h000000AC
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_6                                        'h000000B0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_7                                        'h000000B4
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_8                                        'h000000B8
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_9                                        'h000000BC
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_9__RESERVED0                                    7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_10                                       'h000000C0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_10__RESERVED0                                   7:0
`define CH0_CA_SWI_DQ_RX_IO_M1_R1_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_IO_STA                                                'h000000C4
`define CH0_CA_SWI_DQ_RX_IO_STA__CORE_IG                                             31:0
`define CH0_CA_SWI_DQ_RX_IO_STA___POR                                        32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0                                        'h000000C8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1                                        'h000000CC
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2                                        'h000000D0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3                                        'h000000D4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4                                        'h000000D8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5                                        'h000000DC
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6                                        'h000000E0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7                                        'h000000E4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8                                        'h000000E8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9                                        'h000000EC
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10                                       'h000000F0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R0_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0                                        'h000000F4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1                                        'h000000F8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2                                        'h000000FC
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3                                        'h00000100
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4                                        'h00000104
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5                                        'h00000108
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6                                        'h0000010C
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7                                        'h00000110
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8                                        'h00000114
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9                                        'h00000118
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10                                       'h0000011C
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQ_RX_SA_M0_R1_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0                                        'h00000120
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1                                        'h00000124
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2                                        'h00000128
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3                                        'h0000012C
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4                                        'h00000130
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5                                        'h00000134
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6                                        'h00000138
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7                                        'h0000013C
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8                                        'h00000140
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9                                        'h00000144
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10                                       'h00000148
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R0_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0                                        'h0000014C
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1                                        'h00000150
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2                                        'h00000154
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3                                        'h00000158
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4                                        'h0000015C
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5                                        'h00000160
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6                                        'h00000164
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7                                        'h00000168
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8                                        'h0000016C
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9                                        'h00000170
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_90                                    17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_270                                   19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_180                                   18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_0                                     16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_90                                  7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_270                               15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_180                                11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_0                                   3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_9___POR                                32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10                                       'h00000174
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQ_RX_SA_M1_R1_CFG_10___POR                               32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                    'h00000178
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                    'h0000017C
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                    'h00000180
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                    'h00000184
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                    'h00000188
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                    'h0000018C
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                    'h00000190
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                    'h00000194
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                    'h00000198
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9                                    'h0000019C
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10                                   'h000001A0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_90                                 9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_270                              25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_180                              17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_0                                  1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_90                               15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_270                              31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_180                              23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_0                                  7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10___POR                           32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                    'h000001A4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                    'h000001A8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                    'h000001AC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                    'h000001B0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                    'h000001B4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                    'h000001B8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                    'h000001BC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                    'h000001C0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                    'h000001C4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9                                    'h000001C8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10                                   'h000001CC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_90                                 9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_270                              25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_180                              17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_0                                  1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_90                               15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_270                              31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_180                              23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_0                                  7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10___POR                           32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                    'h000001D0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                    'h000001D4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                    'h000001D8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                    'h000001DC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                    'h000001E0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                    'h000001E4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                    'h000001E8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                    'h000001EC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                    'h000001F0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9                                    'h000001F4
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10                                   'h000001F8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_90                                 9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_270                              25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_180                              17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_0                                  1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_90                               15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_270                              31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_180                              23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_0                                  7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10___POR                           32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                    'h000001FC
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                    'h00000200
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                    'h00000204
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                    'h00000208
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                    'h0000020C
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                    'h00000210
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                    'h00000214
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                    'h00000218
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                    'h0000021C
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9                                    'h00000220
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_90                                  9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_270                               25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_180                               17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_0                                   1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_90                                15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_270                               31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_180                               23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_0                                   7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9___POR                            32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10                                   'h00000224
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_90                                 9:8
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_270                              25:24
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_180                              17:16
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_0                                  1:0
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_90                               15:10
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_270                              31:26
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_180                              23:18
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_0                                  7:2
`define CH0_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10___POR                           32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_0                                              'h00000228
`define CH0_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_0___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_1                                              'h0000022C
`define CH0_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_1___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_2                                              'h00000230
`define CH0_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_2___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_3                                              'h00000234
`define CH0_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_3___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_4                                              'h00000238
`define CH0_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_4___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_5                                              'h0000023C
`define CH0_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_5___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_6                                              'h00000240
`define CH0_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_6___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_7                                              'h00000244
`define CH0_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_7___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_8                                              'h00000248
`define CH0_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_8___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_9                                              'h0000024C
`define CH0_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_90                                            1
`define CH0_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_270                                           3
`define CH0_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_180                                           2
`define CH0_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_0                                             0
`define CH0_CA_SWI_DQ_RX_SA_STA_9___POR                                      32'h00000000

`define CH0_CA_SWI_DQ_RX_SA_STA_10                                             'h00000250
`define CH0_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_90                                           1
`define CH0_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_270                                          3
`define CH0_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_180                                          2
`define CH0_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_0                                            0
`define CH0_CA_SWI_DQ_RX_SA_STA_10___POR                                     32'h00000000

`define CH0_CA_SWI_DQ_TX_BSCAN_CFG                                             'h00000254
`define CH0_CA_SWI_DQ_TX_BSCAN_CFG__VAL                                              10:0
`define CH0_CA_SWI_DQ_TX_BSCAN_CFG___POR                                     32'h00000000

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                   'h00000258
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                   'h0000025C
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                   'h00000260
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                   'h00000264
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                   'h00000268
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                   'h0000026C
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                   'h00000270
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                   'h00000274
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                   'h00000278
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9                                   'h0000027C
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10                                  'h00000280
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10__EGRESS_MODE                            5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10___POR                          32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                   'h00000284
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                   'h00000288
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                   'h0000028C
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                   'h00000290
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                   'h00000294
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                   'h00000298
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                   'h0000029C
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                   'h000002A0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                   'h000002A4
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9                                   'h000002A8
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9__EGRESS_MODE                             5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9___POR                           32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10                                  'h000002AC
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10__EGRESS_MODE                            5:0
`define CH0_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10___POR                          32'h00000001

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                   'h000002B0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                   'h000002B4
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                   'h000002B8
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                   'h000002BC
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                   'h000002C0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                   'h000002C4
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                   'h000002C8
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                   'h000002CC
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                   'h000002D0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9                                   'h000002D4
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10                                  'h000002D8
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10__EGRESS_MODE                            6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10___POR                          32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                   'h000002DC
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                   'h000002E0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                   'h000002E4
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                   'h000002E8
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                   'h000002EC
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                   'h000002F0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                   'h000002F4
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                   'h000002F8
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                   'h000002FC
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9                                   'h00000300
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9__EGRESS_MODE                             6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9___POR                           32'h00000002

`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10                                  'h00000304
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10__EGRESS_MODE                            6:0
`define CH0_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10___POR                          32'h00000002

`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                      'h00000308
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                          14
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                      'h0000030C
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                          14
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                      'h00000310
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                          14
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                      'h00000314
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                          14
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                    'h00000318
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                    'h0000031C
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                    'h00000320
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                    'h00000324
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                    'h00000328
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                    'h0000032C
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                    'h00000330
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                    'h00000334
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                    'h00000338
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                    'h0000033C
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                    'h00000340
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                    'h00000344
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                    'h00000348
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                    'h0000034C
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                    'h00000350
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                    'h00000354
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                   13:10
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                     9:6
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                        14
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                     5:0
`define CH0_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                            32'h00000040

`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG                                       'h00000358
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                      13:10
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                        9:6
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                           14
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                        5:0
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                               32'h00000040

`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG                                       'h0000035C
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                      13:10
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                        9:6
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                           14
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                        5:0
`define CH0_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                               32'h00000040

`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG                                       'h00000360
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                      13:10
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                        9:6
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                           14
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                        5:0
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                               32'h00000040

`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG                                       'h00000364
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                      13:10
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                        9:6
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                           14
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                        5:0
`define CH0_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                               32'h00000040

`define CH0_CA_SWI_DQ_TX_RT_M0_R0_CFG                                          'h00000368
`define CH0_CA_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       10:0
`define CH0_CA_SWI_DQ_TX_RT_M0_R0_CFG___POR                                  32'h00000000

`define CH0_CA_SWI_DQ_TX_RT_M0_R1_CFG                                          'h0000036C
`define CH0_CA_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       10:0
`define CH0_CA_SWI_DQ_TX_RT_M0_R1_CFG___POR                                  32'h00000000

`define CH0_CA_SWI_DQ_TX_RT_M1_R0_CFG                                          'h00000370
`define CH0_CA_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       10:0
`define CH0_CA_SWI_DQ_TX_RT_M1_R0_CFG___POR                                  32'h00000000

`define CH0_CA_SWI_DQ_TX_RT_M1_R1_CFG                                          'h00000374
`define CH0_CA_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       10:0
`define CH0_CA_SWI_DQ_TX_RT_M1_R1_CFG___POR                                  32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0                                       'h00000378
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1                                       'h0000037C
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2                                       'h00000380
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3                                       'h00000384
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4                                       'h00000388
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5                                       'h0000038C
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6                                       'h00000390
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7                                       'h00000394
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8                                       'h00000398
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9                                       'h0000039C
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10                                      'h000003A0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0                                       'h000003A4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1                                       'h000003A8
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2                                       'h000003AC
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3                                       'h000003B0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4                                       'h000003B4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5                                       'h000003B8
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6                                       'h000003BC
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7                                       'h000003C0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8                                       'h000003C4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9                                       'h000003C8
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10                                      'h000003CC
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0                                       'h000003D0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1                                       'h000003D4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2                                       'h000003D8
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3                                       'h000003DC
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4                                       'h000003E0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5                                       'h000003E4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6                                       'h000003E8
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7                                       'h000003EC
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8                                       'h000003F0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9                                       'h000003F4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10                                      'h000003F8
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0                                       'h000003FC
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1                                       'h00000400
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2                                       'h00000404
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3                                       'h00000408
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4                                       'h0000040C
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5                                       'h00000410
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6                                       'h00000414
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7                                       'h00000418
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8                                       'h0000041C
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9                                       'h00000420
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P7                                    7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P6                                    6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P5                                    5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P4                                    4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10                                      'h00000424
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                 'h00000428
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                 'h0000042C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                 'h00000430
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                 'h00000434
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                 'h00000438
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                 'h0000043C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                 'h00000440
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                 'h00000444
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                 'h00000448
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9                                 'h0000044C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10                                'h00000450
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                 'h00000454
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                 'h00000458
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                 'h0000045C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                 'h00000460
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                 'h00000464
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                 'h00000468
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                 'h0000046C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                 'h00000470
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                 'h00000474
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9                                 'h00000478
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10                                'h0000047C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                 'h00000480
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                 'h00000484
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                 'h00000488
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                 'h0000048C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                 'h00000490
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                 'h00000494
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                 'h00000498
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                 'h0000049C
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                 'h000004A0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9                                 'h000004A4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10                                'h000004A8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                 'h000004AC
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                 'h000004B0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                 'h000004B4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                 'h000004B8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                 'h000004BC
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                 'h000004C0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                 'h000004C4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                 'h000004C8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                 'h000004CC
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9                                 'h000004D0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P7                            30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P6                            26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P5                            22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P4                            18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P3                            14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P2                             10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                              6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                              2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10                                'h000004D4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                                'h000004D8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                                'h000004DC
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                                'h000004E0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                                'h000004E4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                                'h000004E8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                                'h000004EC
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                                'h000004F0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                                'h000004F4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                                'h000004F8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9                                'h000004FC
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10                               'h00000500
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P7                            29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P6                            25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P5                            21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P4                            17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P3                            13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P2                              9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P1                              5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P0                              1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10___POR                       32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                                'h00000504
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                                'h00000508
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                                'h0000050C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                                'h00000510
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                                'h00000514
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                                'h00000518
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                                'h0000051C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                                'h00000520
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                                'h00000524
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9                                'h00000528
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10                               'h0000052C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P7                            29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P6                            25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P5                            21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P4                            17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P3                            13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P2                              9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P1                              5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P0                              1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10___POR                       32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                                'h00000530
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                                'h00000534
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                                'h00000538
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                                'h0000053C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                                'h00000540
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                                'h00000544
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                                'h00000548
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                                'h0000054C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                                'h00000550
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9                                'h00000554
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10                               'h00000558
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P7                            29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P6                            25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P5                            21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P4                            17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P3                            13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P2                              9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P1                              5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P0                              1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10___POR                       32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                                'h0000055C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                                'h00000560
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                                'h00000564
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                                'h00000568
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                                'h0000056C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                                'h00000570
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                                'h00000574
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                                'h00000578
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                                'h0000057C
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9                                'h00000580
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P7                             29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P6                             25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P5                             21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P4                             17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P3                             13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P2                               9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P1                               5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P0                               1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10                               'h00000584
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P7                            29:28
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P6                            25:24
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P5                            21:20
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P4                            17:16
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P3                            13:12
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P2                              9:8
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P1                              5:4
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P0                              1:0
`define CH0_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10___POR                       32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0                                       'h00000588
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1                                       'h0000058C
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2                                       'h00000590
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3                                       'h00000594
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4                                       'h00000598
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5                                       'h0000059C
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6                                       'h000005A0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7                                       'h000005A4
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8                                       'h000005A8
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9                                       'h000005AC
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10                                      'h000005B0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0                                       'h000005B4
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1                                       'h000005B8
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2                                       'h000005BC
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3                                       'h000005C0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4                                       'h000005C4
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5                                       'h000005C8
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6                                       'h000005CC
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7                                       'h000005D0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8                                       'h000005D4
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9                                       'h000005D8
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10                                      'h000005DC
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0                                       'h000005E0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1                                       'h000005E4
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2                                       'h000005E8
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3                                       'h000005EC
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4                                       'h000005F0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5                                       'h000005F4
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6                                       'h000005F8
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7                                       'h000005FC
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8                                       'h00000600
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9                                       'h00000604
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10                                      'h00000608
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0                                       'h0000060C
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1                                       'h00000610
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2                                       'h00000614
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3                                       'h00000618
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4                                       'h0000061C
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5                                       'h00000620
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6                                       'h00000624
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7                                       'h00000628
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8                                       'h0000062C
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9                                       'h00000630
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P3                                    3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P2                                    2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10                                      'h00000634
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                 'h00000638
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                 'h0000063C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                 'h00000640
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                 'h00000644
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                 'h00000648
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                 'h0000064C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                 'h00000650
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                 'h00000654
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                 'h00000658
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9                                 'h0000065C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10                                'h00000660
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                 'h00000664
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                 'h00000668
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                 'h0000066C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                 'h00000670
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                 'h00000674
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                 'h00000678
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                 'h0000067C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                 'h00000680
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                 'h00000684
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9                                 'h00000688
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10                                'h0000068C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                 'h00000690
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                 'h00000694
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                 'h00000698
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                 'h0000069C
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                 'h000006A0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                 'h000006A4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                 'h000006A8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                 'h000006AC
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                 'h000006B0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9                                 'h000006B4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10                                'h000006B8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                 'h000006BC
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                 'h000006C0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                 'h000006C4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                 'h000006C8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                 'h000006CC
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                 'h000006D0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                 'h000006D4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                 'h000006D8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                 'h000006DC
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9                                 'h000006E0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P3                            13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P2                              9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                              5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                              1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10                                'h000006E4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0                                       'h000006E8
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1                                       'h000006EC
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2                                       'h000006F0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3                                       'h000006F4
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4                                       'h000006F8
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5                                       'h000006FC
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6                                       'h00000700
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7                                       'h00000704
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8                                       'h00000708
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9                                       'h0000070C
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10                                      'h00000710
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0                                       'h00000714
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1                                       'h00000718
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2                                       'h0000071C
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3                                       'h00000720
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4                                       'h00000724
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5                                       'h00000728
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6                                       'h0000072C
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7                                       'h00000730
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8                                       'h00000734
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9                                       'h00000738
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10                                      'h0000073C
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0                                       'h00000740
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1                                       'h00000744
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2                                       'h00000748
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3                                       'h0000074C
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4                                       'h00000750
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5                                       'h00000754
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6                                       'h00000758
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7                                       'h0000075C
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8                                       'h00000760
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9                                       'h00000764
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10                                      'h00000768
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0                                       'h0000076C
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1                                       'h00000770
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2                                       'h00000774
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3                                       'h00000778
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4                                       'h0000077C
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5                                       'h00000780
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6                                       'h00000784
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7                                       'h00000788
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8                                       'h0000078C
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9                                       'h00000790
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10                                      'h00000794
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                 'h00000798
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                 'h0000079C
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                 'h000007A0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                 'h000007A4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                 'h000007A8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                 'h000007AC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                 'h000007B0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                 'h000007B4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                 'h000007B8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9                                 'h000007BC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10                                'h000007C0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                               4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                               0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                 'h000007C4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                 'h000007C8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                 'h000007CC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                 'h000007D0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                 'h000007D4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                 'h000007D8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                 'h000007DC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                 'h000007E0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                 'h000007E4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9                                 'h000007E8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10                                'h000007EC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                               4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                               0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                 'h000007F0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                 'h000007F4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                 'h000007F8
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                 'h000007FC
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                 'h00000800
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                 'h00000804
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                 'h00000808
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                 'h0000080C
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                 'h00000810
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9                                 'h00000814
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10                                'h00000818
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                               4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                               0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                 'h0000081C
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                 'h00000820
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                 'h00000824
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                 'h00000828
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                 'h0000082C
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                 'h00000830
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                 'h00000834
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                 'h00000838
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                 'h0000083C
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9                                 'h00000840
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                                4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                                0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10                                'h00000844
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                               4
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                               0
`define CH0_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                      'h00000848
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                      'h0000084C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                      'h00000850
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                      'h00000854
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                      'h00000858
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                      'h0000085C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                      'h00000860
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                      'h00000864
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                      'h00000868
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9                                      'h0000086C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10                                     'h00000870
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__GEAR                                      7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__EN                                          8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10___POR                             32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                      'h00000874
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                      'h00000878
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                      'h0000087C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                      'h00000880
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                      'h00000884
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                      'h00000888
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                      'h0000088C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                      'h00000890
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                      'h00000894
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9                                      'h00000898
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10                                     'h0000089C
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__GEAR                                      7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__EN                                          8
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10___POR                             32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                      'h000008A0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                      'h000008A4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                      'h000008A8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                      'h000008AC
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                      'h000008B0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                      'h000008B4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                      'h000008B8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                      'h000008BC
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                      'h000008C0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9                                      'h000008C4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10                                     'h000008C8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__GEAR                                      7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__EN                                          8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10___POR                             32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                      'h000008CC
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                      'h000008D0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                      'h000008D4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                      'h000008D8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                      'h000008DC
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                      'h000008E0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                      'h000008E4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                      'h000008E8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                      'h000008EC
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9                                      'h000008F0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__GEAR                                       7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__EN                                           8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__CTRL_BIN                                   5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9___POR                              32'h00000100

`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10                                     'h000008F4
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__GEAR                                      7:6
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__EN                                          8
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10___POR                             32'h00000100

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0                                           'h000008F8
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_0___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1                                           'h000008FC
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_1___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2                                           'h00000900
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_2___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3                                           'h00000904
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_3___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4                                           'h00000908
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_4___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5                                           'h0000090C
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_5___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6                                           'h00000910
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_6___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7                                           'h00000914
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_7___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8                                           'h00000918
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_8___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9                                           'h0000091C
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_9___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10                                          'h00000920
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__TX_IMPD                                        8:6
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__SW_OVR                                           5
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__RX_IMPD                                       11:9
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__RESERVED0                                        4
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__OVRD_VAL                                         3
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10__OVRD_SEL                                       2:0
`define CH0_CA_SWI_DQ_TX_IO_M0_CFG_10___POR                                  32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0                                           'h00000924
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_0___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1                                           'h00000928
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_1___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2                                           'h0000092C
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_2___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3                                           'h00000930
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_3___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4                                           'h00000934
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_4___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5                                           'h00000938
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_5___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6                                           'h0000093C
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_6___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7                                           'h00000940
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_7___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8                                           'h00000944
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_8___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9                                           'h00000948
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__TX_IMPD                                         8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__SW_OVR                                            5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__RX_IMPD                                        11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__RESERVED0                                         4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__OVRD_VAL                                          3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9__OVRD_SEL                                        2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_9___POR                                   32'h00000040

`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10                                          'h0000094C
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__TX_IMPD                                        8:6
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__SW_OVR                                           5
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__RX_IMPD                                       11:9
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__RESERVED0                                        4
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__OVRD_VAL                                         3
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10__OVRD_SEL                                       2:0
`define CH0_CA_SWI_DQ_TX_IO_M1_CFG_10___POR                                  32'h00000040

`define CH0_CA_SWI_DQS_RX_M0_CFG                                               'h00000950
`define CH0_CA_SWI_DQS_RX_M0_CFG__WCK_MODE                                              8
`define CH0_CA_SWI_DQS_RX_M0_CFG__RGB_MODE                                            2:0
`define CH0_CA_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                    13:12
`define CH0_CA_SWI_DQS_RX_M0_CFG__FGB_MODE                                            7:4
`define CH0_CA_SWI_DQS_RX_M0_CFG___POR                                       32'h00000074

`define CH0_CA_SWI_DQS_RX_M1_CFG                                               'h00000954
`define CH0_CA_SWI_DQS_RX_M1_CFG__WCK_MODE                                              8
`define CH0_CA_SWI_DQS_RX_M1_CFG__RGB_MODE                                            2:0
`define CH0_CA_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                    13:12
`define CH0_CA_SWI_DQS_RX_M1_CFG__FGB_MODE                                            7:4
`define CH0_CA_SWI_DQS_RX_M1_CFG___POR                                       32'h00000074

`define CH0_CA_SWI_DQS_RX_BSCAN_STA                                            'h00000958
`define CH0_CA_SWI_DQS_RX_BSCAN_STA__VAL                                              1:0
`define CH0_CA_SWI_DQS_RX_BSCAN_STA___POR                                    32'h00000000

`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                   'h0000095C
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                    7:6
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                        8
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                                5:0
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                           32'h00000100

`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                   'h00000960
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                    7:6
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                        8
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                                5:0
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                           32'h00000100

`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                   'h00000964
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                    7:6
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                        8
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                                5:0
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                           32'h00000100

`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                   'h00000968
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                    7:6
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                        8
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                                5:0
`define CH0_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                           32'h00000100

`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG                                     'h0000096C
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG                                     'h00000970
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG                                     'h00000974
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG                                     'h00000978
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                     'h0000097C
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                     'h00000980
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                     'h00000984
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                     'h00000988
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                  'h0000098C
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                  'h00000990
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                  'h00000994
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                  'h00000998
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                  'h0000099C
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                  'h000009A0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                  'h000009A4
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                  'h000009A8
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                      14
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH0_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH0_CA_SWI_DQS_RX_PI_STA                                               'h000009AC
`define CH0_CA_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                          0
`define CH0_CA_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                          1
`define CH0_CA_SWI_DQS_RX_PI_STA___POR                                       32'h00000000

`define CH0_CA_SWI_DQS_RX_IO_M0_R0_CFG_0                                       'h000009B0
`define CH0_CA_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                 15:8
`define CH0_CA_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                  7:0
`define CH0_CA_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_IO_M0_R1_CFG_0                                       'h000009B4
`define CH0_CA_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                 15:8
`define CH0_CA_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                  7:0
`define CH0_CA_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_IO_M1_R0_CFG_0                                       'h000009B8
`define CH0_CA_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                 15:8
`define CH0_CA_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                  7:0
`define CH0_CA_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_IO_M1_R1_CFG_0                                       'h000009BC
`define CH0_CA_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                 15:8
`define CH0_CA_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                  7:0
`define CH0_CA_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                     'h000009C0
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                     23
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                    22
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                   21
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                   18:16
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                         20
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                  19
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                   7:4
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                   3:0
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                 15:12
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                  11:8
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                             32'h004A7777

`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                     'h000009C4
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                     23
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                    22
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                   21
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                   18:16
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                         20
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                  19
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                   7:4
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                   3:0
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                 15:12
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                  11:8
`define CH0_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                             32'h004A7777

`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                     'h000009C8
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                     23
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                    22
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                   21
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                   18:16
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                         20
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                  19
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                   7:4
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                   3:0
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                 15:12
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                  11:8
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                             32'h004A7777

`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                     'h000009CC
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                     23
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                    22
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                   21
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                   18:16
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                         20
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                  19
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                   7:4
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                   3:0
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                 15:12
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                  11:8
`define CH0_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                             32'h004A7777

`define CH0_CA_SWI_DQS_RX_IO_STA                                               'h000009D0
`define CH0_CA_SWI_DQS_RX_IO_STA__CORE_IG                                            31:0
`define CH0_CA_SWI_DQS_RX_IO_STA___POR                                       32'h00000000

`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0                                       'h000009D4
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0                                       'h000009D8
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0                                       'h000009DC
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0                                       'h000009E0
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH0_CA_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG                                           'h000009E4
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                            4
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                     2
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                      0
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                     3
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                      1
`define CH0_CA_SWI_DQS_RX_SA_CMN_CFG___POR                                   32'h00000005

`define CH0_CA_SWI_DQS_TX_M0_CFG                                               'h000009E8
`define CH0_CA_SWI_DQS_TX_M0_CFG__WGB_MODE                                            7:4
`define CH0_CA_SWI_DQS_TX_M0_CFG__TGB_MODE                                            2:0
`define CH0_CA_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                        9:8
`define CH0_CA_SWI_DQS_TX_M0_CFG___POR                                       32'h00000087

`define CH0_CA_SWI_DQS_TX_M1_CFG                                               'h000009EC
`define CH0_CA_SWI_DQS_TX_M1_CFG__WGB_MODE                                            7:4
`define CH0_CA_SWI_DQS_TX_M1_CFG__TGB_MODE                                            2:0
`define CH0_CA_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                        9:8
`define CH0_CA_SWI_DQS_TX_M1_CFG___POR                                       32'h00000087

`define CH0_CA_SWI_DQS_TX_BSCAN_CTRL_CFG                                       'h000009F0
`define CH0_CA_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                            1
`define CH0_CA_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                            0
`define CH0_CA_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                               32'h00000000

`define CH0_CA_SWI_DQS_TX_BSCAN_CFG                                            'h000009F4
`define CH0_CA_SWI_DQS_TX_BSCAN_CFG__VAL                                              1:0
`define CH0_CA_SWI_DQS_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                  'h000009F8
`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                  'h000009FC
`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH0_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                  'h00000A00
`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                  'h00000A04
`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH0_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                     'h00000A08
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                     'h00000A0C
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                     'h00000A10
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                     'h00000A14
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH0_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                   'h00000A18
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                   'h00000A1C
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                   'h00000A20
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                   'h00000A24
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                   'h00000A28
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                   'h00000A2C
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                   'h00000A30
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                   'h00000A34
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                   'h00000A38
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                   'h00000A3C
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                   'h00000A40
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                   'h00000A44
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                   'h00000A48
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                   'h00000A4C
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                   'h00000A50
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                   'h00000A54
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH0_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG                                      'h00000A58
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG                                      'h00000A5C
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG                                      'h00000A60
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG                                      'h00000A64
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH0_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                     'h00000A68
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                     'h00000A6C
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                     'h00000A70
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                     'h00000A74
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                     'h00000A78
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                     'h00000A7C
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                     'h00000A80
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                     'h00000A84
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                    13:10
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                      5:0
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                      9:6
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                         14
`define CH0_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                             32'h00000040

`define CH0_CA_SWI_DQS_TX_RT_M0_R0_CFG                                         'h00000A88
`define CH0_CA_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                         0
`define CH0_CA_SWI_DQS_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH0_CA_SWI_DQS_TX_RT_M0_R1_CFG                                         'h00000A8C
`define CH0_CA_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                         0
`define CH0_CA_SWI_DQS_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH0_CA_SWI_DQS_TX_RT_M1_R0_CFG                                         'h00000A90
`define CH0_CA_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                         0
`define CH0_CA_SWI_DQS_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH0_CA_SWI_DQS_TX_RT_M1_R1_CFG                                         'h00000A94
`define CH0_CA_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                         0
`define CH0_CA_SWI_DQS_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0                                      'h00000A98
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0                                      'h00000A9C
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0                                      'h00000AA0
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0                                      'h00000AA4
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000AA8
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                                'h00000AAC
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                                'h00000AB0
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                                'h00000AB4
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH0_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000AB8
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000ABC
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000AC0
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h00000AC4
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH0_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0                                      'h00000AC8
`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0                                      'h00000ACC
`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0                                      'h00000AD0
`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0                                      'h00000AD4
`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000AD8
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000ADC
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000AE0
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                                'h00000AE4
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH0_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0                                      'h00000AE8
`define CH0_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0                                      'h00000AEC
`define CH0_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0                                      'h00000AF0
`define CH0_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0                                      'h00000AF4
`define CH0_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH0_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH0_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000AF8
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000AFC
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000B00
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                                'h00000B04
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH0_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH0_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                     'h00000B08
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH0_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                     'h00000B0C
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH0_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                     'h00000B10
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH0_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                     'h00000B14
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH0_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0                                          'h00000B18
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                       4
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                       3
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH0_CA_SWI_DQS_TX_IO_M0_CFG_0___POR                                  32'h00000041

`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0                                          'h00000B1C
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                       4
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                       3
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH0_CA_SWI_DQS_TX_IO_M1_CFG_0___POR                                  32'h00000041

`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                     'h00000B20
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                    13
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                     10:5
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                      4:0
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                    12
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                      11
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                             32'h00000001

`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                     'h00000B24
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                    13
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                     10:5
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                      4:0
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                    12
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                      11
`define CH0_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                             32'h00000001

`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                     'h00000B28
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                    13
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                     10:5
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                      4:0
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                    12
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                      11
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                             32'h00000001

`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                     'h00000B2C
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                    13
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                     10:5
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                      4:0
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                    12
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                      11
`define CH0_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                             32'h00000001

`define CH1_DQ0_SWI_TOP_CFG                                                    'h00000000
`define CH1_DQ0_SWI_TOP_CFG__WCS_SW_OVR_VAL                                             1
`define CH1_DQ0_SWI_TOP_CFG__WCS_SW_OVR                                                 0
`define CH1_DQ0_SWI_TOP_CFG__TRAINING_MODE                                              9
`define CH1_DQ0_SWI_TOP_CFG__RCS_SW_OVR_VAL                                             3
`define CH1_DQ0_SWI_TOP_CFG__RCS_SW_OVR                                                 2
`define CH1_DQ0_SWI_TOP_CFG__FIFO_CLR                                                   8
`define CH1_DQ0_SWI_TOP_CFG___POR                                            32'h00000000

`define CH1_DQ0_SWI_TOP_STA                                                    'h00000004
`define CH1_DQ0_SWI_TOP_STA__WCS                                                        0
`define CH1_DQ0_SWI_TOP_STA__RCS                                                        1
`define CH1_DQ0_SWI_TOP_STA___POR                                            32'h00000000

`define CH1_DQ0_SWI_DQ_RX_BSCAN_STA                                            'h00000008
`define CH1_DQ0_SWI_DQ_RX_BSCAN_STA__VAL                                              8:0
`define CH1_DQ0_SWI_DQ_RX_BSCAN_STA___POR                                    32'h00000000

`define CH1_DQ0_SWI_DQ_RX_M0_CFG                                               'h0000000C
`define CH1_DQ0_SWI_DQ_RX_M0_CFG__RGB_MODE                                            2:0
`define CH1_DQ0_SWI_DQ_RX_M0_CFG__FGB_MODE                                            7:4
`define CH1_DQ0_SWI_DQ_RX_M0_CFG___POR                                       32'h00000074

`define CH1_DQ0_SWI_DQ_RX_M1_CFG                                               'h00000010
`define CH1_DQ0_SWI_DQ_RX_M1_CFG__RGB_MODE                                            2:0
`define CH1_DQ0_SWI_DQ_RX_M1_CFG__FGB_MODE                                            7:4
`define CH1_DQ0_SWI_DQ_RX_M1_CFG___POR                                       32'h00000074

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0                                       'h00000014
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1                                       'h00000018
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2                                       'h0000001C
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3                                       'h00000020
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4                                       'h00000024
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5                                       'h00000028
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6                                       'h0000002C
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7                                       'h00000030
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8                                       'h00000034
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0                                       'h00000038
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1                                       'h0000003C
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2                                       'h00000040
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3                                       'h00000044
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4                                       'h00000048
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5                                       'h0000004C
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6                                       'h00000050
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7                                       'h00000054
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8                                       'h00000058
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0                                       'h0000005C
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1                                       'h00000060
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2                                       'h00000064
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3                                       'h00000068
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4                                       'h0000006C
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5                                       'h00000070
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6                                       'h00000074
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7                                       'h00000078
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8                                       'h0000007C
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0                                       'h00000080
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1                                       'h00000084
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2                                       'h00000088
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3                                       'h0000008C
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4                                       'h00000090
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5                                       'h00000094
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6                                       'h00000098
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7                                       'h0000009C
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8                                       'h000000A0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                   7:0
`define CH1_DQ0_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_IO_STA                                               'h000000A4
`define CH1_DQ0_SWI_DQ_RX_IO_STA__CORE_IG                                            31:0
`define CH1_DQ0_SWI_DQ_RX_IO_STA___POR                                       32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0                                       'h000000A8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1                                       'h000000AC
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2                                       'h000000B0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3                                       'h000000B4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4                                       'h000000B8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5                                       'h000000BC
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6                                       'h000000C0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7                                       'h000000C4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8                                       'h000000C8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0                                       'h000000CC
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1                                       'h000000D0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2                                       'h000000D4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3                                       'h000000D8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4                                       'h000000DC
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5                                       'h000000E0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6                                       'h000000E4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7                                       'h000000E8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8                                       'h000000EC
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0                                       'h000000F0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1                                       'h000000F4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2                                       'h000000F8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3                                       'h000000FC
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4                                       'h00000100
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5                                       'h00000104
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6                                       'h00000108
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7                                       'h0000010C
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8                                       'h00000110
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0                                       'h00000114
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1                                       'h00000118
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2                                       'h0000011C
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3                                       'h00000120
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4                                       'h00000124
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5                                       'h00000128
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6                                       'h0000012C
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7                                       'h00000130
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8                                       'h00000134
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ0_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                   'h00000138
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                   'h0000013C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                   'h00000140
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                   'h00000144
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                   'h00000148
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                   'h0000014C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                   'h00000150
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                   'h00000154
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                   'h00000158
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                   'h0000015C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                   'h00000160
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                   'h00000164
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                   'h00000168
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                   'h0000016C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                   'h00000170
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                   'h00000174
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                   'h00000178
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                   'h0000017C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                   'h00000180
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                   'h00000184
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                   'h00000188
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                   'h0000018C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                   'h00000190
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                   'h00000194
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                   'h00000198
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                   'h0000019C
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                   'h000001A0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                   'h000001A4
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                   'h000001A8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                   'h000001AC
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                   'h000001B0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                   'h000001B4
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                   'h000001B8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                   'h000001BC
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                   'h000001C0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                   'h000001C4
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                 9:8
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                              25:24
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                              17:16
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                  1:0
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                               15:10
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                              31:26
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                              23:18
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                  7:2
`define CH1_DQ0_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                           32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_0                                             'h000001C8
`define CH1_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_0___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_1                                             'h000001CC
`define CH1_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_1___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_2                                             'h000001D0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_2___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_3                                             'h000001D4
`define CH1_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_3___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_4                                             'h000001D8
`define CH1_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_4___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_5                                             'h000001DC
`define CH1_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_5___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_6                                             'h000001E0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_6___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_7                                             'h000001E4
`define CH1_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_7___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_RX_SA_STA_8                                             'h000001E8
`define CH1_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                           1
`define CH1_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                          3
`define CH1_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                          2
`define CH1_DQ0_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                            0
`define CH1_DQ0_SWI_DQ_RX_SA_STA_8___POR                                     32'h00000000

`define CH1_DQ0_SWI_DQ_TX_BSCAN_CFG                                            'h000001EC
`define CH1_DQ0_SWI_DQ_TX_BSCAN_CFG__VAL                                              8:0
`define CH1_DQ0_SWI_DQ_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                  'h000001F0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                  'h000001F4
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                  'h000001F8
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                  'h000001FC
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                  'h00000200
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                  'h00000204
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                  'h00000208
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                  'h0000020C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                  'h00000210
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                  'h00000214
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                  'h00000218
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                  'h0000021C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                  'h00000220
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                  'h00000224
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                  'h00000228
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                  'h0000022C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                  'h00000230
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                  'h00000234
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                            5:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                          32'h00000001

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                  'h00000238
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                  'h0000023C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                  'h00000240
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                  'h00000244
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                  'h00000248
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                  'h0000024C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                  'h00000250
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                  'h00000254
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                  'h00000258
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                  'h0000025C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                  'h00000260
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                  'h00000264
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                  'h00000268
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                  'h0000026C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                  'h00000270
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                  'h00000274
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                  'h00000278
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                  'h0000027C
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                            6:0
`define CH1_DQ0_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                          32'h00000002

`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                     'h00000280
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                     'h00000284
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                     'h00000288
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                     'h0000028C
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                   'h00000290
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                   'h00000294
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                   'h00000298
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                   'h0000029C
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                   'h000002A0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                   'h000002A4
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                   'h000002A8
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                   'h000002AC
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                   'h000002B0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                   'h000002B4
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                   'h000002B8
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                   'h000002BC
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                   'h000002C0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                   'h000002C4
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                   'h000002C8
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                   'h000002CC
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ0_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG                                      'h000002D0
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG                                      'h000002D4
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG                                      'h000002D8
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG                                      'h000002DC
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH1_DQ0_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH1_DQ0_SWI_DQ_TX_RT_M0_R0_CFG                                         'h000002E0
`define CH1_DQ0_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       8:0
`define CH1_DQ0_SWI_DQ_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH1_DQ0_SWI_DQ_TX_RT_M0_R1_CFG                                         'h000002E4
`define CH1_DQ0_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       8:0
`define CH1_DQ0_SWI_DQ_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH1_DQ0_SWI_DQ_TX_RT_M1_R0_CFG                                         'h000002E8
`define CH1_DQ0_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       8:0
`define CH1_DQ0_SWI_DQ_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH1_DQ0_SWI_DQ_TX_RT_M1_R1_CFG                                         'h000002EC
`define CH1_DQ0_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       8:0
`define CH1_DQ0_SWI_DQ_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0                                      'h000002F0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1                                      'h000002F4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2                                      'h000002F8
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3                                      'h000002FC
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4                                      'h00000300
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5                                      'h00000304
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6                                      'h00000308
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7                                      'h0000030C
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8                                      'h00000310
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0                                      'h00000314
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1                                      'h00000318
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2                                      'h0000031C
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3                                      'h00000320
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4                                      'h00000324
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5                                      'h00000328
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6                                      'h0000032C
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7                                      'h00000330
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8                                      'h00000334
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0                                      'h00000338
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1                                      'h0000033C
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2                                      'h00000340
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3                                      'h00000344
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4                                      'h00000348
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5                                      'h0000034C
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6                                      'h00000350
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7                                      'h00000354
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8                                      'h00000358
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0                                      'h0000035C
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1                                      'h00000360
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2                                      'h00000364
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3                                      'h00000368
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4                                      'h0000036C
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5                                      'h00000370
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6                                      'h00000374
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7                                      'h00000378
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8                                      'h0000037C
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000380
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                'h00000384
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                'h00000388
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                'h0000038C
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                'h00000390
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                'h00000394
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                'h00000398
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                'h0000039C
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                'h000003A0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                'h000003A4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                'h000003A8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                'h000003AC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                'h000003B0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                'h000003B4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                'h000003B8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                'h000003BC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                'h000003C0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                'h000003C4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                'h000003C8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                'h000003CC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                'h000003D0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                'h000003D4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                'h000003D8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                'h000003DC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                'h000003E0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                'h000003E4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                'h000003E8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                'h000003EC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                'h000003F0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                'h000003F4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                'h000003F8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                'h000003FC
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                'h00000400
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                'h00000404
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                'h00000408
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                'h0000040C
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ0_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000410
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                               'h00000414
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                               'h00000418
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                               'h0000041C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                               'h00000420
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                               'h00000424
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                               'h00000428
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                               'h0000042C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                               'h00000430
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000434
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                               'h00000438
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                               'h0000043C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                               'h00000440
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                               'h00000444
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                               'h00000448
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                               'h0000044C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                               'h00000450
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                               'h00000454
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000458
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                               'h0000045C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                               'h00000460
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                               'h00000464
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                               'h00000468
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                               'h0000046C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                               'h00000470
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                               'h00000474
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                               'h00000478
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h0000047C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                               'h00000480
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                               'h00000484
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                               'h00000488
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                               'h0000048C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                               'h00000490
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                               'h00000494
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                               'h00000498
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                               'h0000049C
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                            29:28
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                            25:24
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                            21:20
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                            17:16
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                            13:12
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                              9:8
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                              5:4
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                              1:0
`define CH1_DQ0_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0                                      'h000004A0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1                                      'h000004A4
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2                                      'h000004A8
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3                                      'h000004AC
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4                                      'h000004B0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5                                      'h000004B4
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6                                      'h000004B8
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7                                      'h000004BC
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8                                      'h000004C0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0                                      'h000004C4
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1                                      'h000004C8
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2                                      'h000004CC
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3                                      'h000004D0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4                                      'h000004D4
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5                                      'h000004D8
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6                                      'h000004DC
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7                                      'h000004E0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8                                      'h000004E4
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0                                      'h000004E8
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1                                      'h000004EC
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2                                      'h000004F0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3                                      'h000004F4
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4                                      'h000004F8
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5                                      'h000004FC
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6                                      'h00000500
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7                                      'h00000504
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8                                      'h00000508
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0                                      'h0000050C
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1                                      'h00000510
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2                                      'h00000514
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3                                      'h00000518
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4                                      'h0000051C
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5                                      'h00000520
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6                                      'h00000524
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7                                      'h00000528
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8                                      'h0000052C
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000530
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                'h00000534
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                'h00000538
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                'h0000053C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                'h00000540
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                'h00000544
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                'h00000548
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                'h0000054C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                'h00000550
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000554
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                'h00000558
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                'h0000055C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                'h00000560
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                'h00000564
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                'h00000568
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                'h0000056C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                'h00000570
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                'h00000574
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000578
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                'h0000057C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                'h00000580
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                'h00000584
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                'h00000588
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                'h0000058C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                'h00000590
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                'h00000594
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                'h00000598
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                'h0000059C
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                'h000005A0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                'h000005A4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                'h000005A8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                'h000005AC
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                'h000005B0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                'h000005B4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                'h000005B8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                'h000005BC
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ0_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0                                      'h000005C0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1                                      'h000005C4
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2                                      'h000005C8
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3                                      'h000005CC
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4                                      'h000005D0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5                                      'h000005D4
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6                                      'h000005D8
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7                                      'h000005DC
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8                                      'h000005E0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0                                      'h000005E4
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1                                      'h000005E8
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2                                      'h000005EC
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3                                      'h000005F0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4                                      'h000005F4
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5                                      'h000005F8
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6                                      'h000005FC
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7                                      'h00000600
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8                                      'h00000604
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0                                      'h00000608
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1                                      'h0000060C
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2                                      'h00000610
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3                                      'h00000614
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4                                      'h00000618
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5                                      'h0000061C
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6                                      'h00000620
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7                                      'h00000624
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8                                      'h00000628
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0                                      'h0000062C
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1                                      'h00000630
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2                                      'h00000634
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3                                      'h00000638
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4                                      'h0000063C
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5                                      'h00000640
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6                                      'h00000644
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7                                      'h00000648
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8                                      'h0000064C
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ0_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000650
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                'h00000654
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                'h00000658
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                'h0000065C
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                'h00000660
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                'h00000664
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                'h00000668
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                'h0000066C
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                'h00000670
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000674
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                'h00000678
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                'h0000067C
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                'h00000680
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                'h00000684
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                'h00000688
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                'h0000068C
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                'h00000690
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                'h00000694
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000698
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                'h0000069C
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                'h000006A0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                'h000006A4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                'h000006A8
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                'h000006AC
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                'h000006B0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                'h000006B4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                'h000006B8
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                'h000006BC
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                'h000006C0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                'h000006C4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                'h000006C8
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                'h000006CC
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                'h000006D0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                'h000006D4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                'h000006D8
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                'h000006DC
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                               4
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                               0
`define CH1_DQ0_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                     'h000006E0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                     'h000006E4
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                     'h000006E8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                     'h000006EC
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                     'h000006F0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                     'h000006F4
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                     'h000006F8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                     'h000006FC
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                     'h00000700
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                     'h00000704
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                     'h00000708
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                     'h0000070C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                     'h00000710
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                     'h00000714
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                     'h00000718
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                     'h0000071C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                     'h00000720
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                     'h00000724
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                     'h00000728
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                     'h0000072C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                     'h00000730
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                     'h00000734
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                     'h00000738
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                     'h0000073C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                     'h00000740
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                     'h00000744
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                     'h00000748
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                     'h0000074C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                     'h00000750
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                     'h00000754
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                     'h00000758
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                     'h0000075C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                     'h00000760
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                     'h00000764
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                     'h00000768
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                     'h0000076C
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                      7:6
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                          8
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ0_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                             32'h00000100

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0                                          'h00000770
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_0___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1                                          'h00000774
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_1___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2                                          'h00000778
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_2___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3                                          'h0000077C
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_3___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4                                          'h00000780
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_4___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5                                          'h00000784
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_5___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6                                          'h00000788
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_6___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7                                          'h0000078C
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_7___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8                                          'h00000790
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M0_CFG_8___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0                                          'h00000794
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_0___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1                                          'h00000798
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_1___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2                                          'h0000079C
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_2___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3                                          'h000007A0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_3___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4                                          'h000007A4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_4___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5                                          'h000007A8
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_5___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6                                          'h000007AC
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_6___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7                                          'h000007B0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_7___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8                                          'h000007B4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                        8:6
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                           5
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                       11:9
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                        4
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                         3
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                       2:0
`define CH1_DQ0_SWI_DQ_TX_IO_M1_CFG_8___POR                                  32'h00000040

`define CH1_DQ0_SWI_DQS_RX_M0_CFG                                              'h000007B8
`define CH1_DQ0_SWI_DQS_RX_M0_CFG__WCK_MODE                                             8
`define CH1_DQ0_SWI_DQS_RX_M0_CFG__RGB_MODE                                           2:0
`define CH1_DQ0_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                   13:12
`define CH1_DQ0_SWI_DQS_RX_M0_CFG__FGB_MODE                                           7:4
`define CH1_DQ0_SWI_DQS_RX_M0_CFG___POR                                      32'h00000074

`define CH1_DQ0_SWI_DQS_RX_M1_CFG                                              'h000007BC
`define CH1_DQ0_SWI_DQS_RX_M1_CFG__WCK_MODE                                             8
`define CH1_DQ0_SWI_DQS_RX_M1_CFG__RGB_MODE                                           2:0
`define CH1_DQ0_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                   13:12
`define CH1_DQ0_SWI_DQS_RX_M1_CFG__FGB_MODE                                           7:4
`define CH1_DQ0_SWI_DQS_RX_M1_CFG___POR                                      32'h00000074

`define CH1_DQ0_SWI_DQS_RX_BSCAN_STA                                           'h000007C0
`define CH1_DQ0_SWI_DQS_RX_BSCAN_STA__VAL                                             3:0
`define CH1_DQ0_SWI_DQS_RX_BSCAN_STA___POR                                   32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                  'h000007C4
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                   7:6
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                       8
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                               5:0
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                          32'h00000100

`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                  'h000007C8
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                   7:6
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                       8
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                               5:0
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                          32'h00000100

`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                  'h000007CC
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                   7:6
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                       8
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                               5:0
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                          32'h00000100

`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                  'h000007D0
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                   7:6
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                       8
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                               5:0
`define CH1_DQ0_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                          32'h00000100

`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG                                    'h000007D4
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG                                    'h000007D8
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG                                    'h000007DC
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG                                    'h000007E0
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                    'h000007E4
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                    'h000007E8
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                    'h000007EC
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                    'h000007F0
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                 'h000007F4
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                 'h000007F8
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                 'h000007FC
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                 'h00000800
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                 'h00000804
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                 'h00000808
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                 'h0000080C
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                 'h00000810
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                13:10
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                  9:6
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                     14
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                  5:0
`define CH1_DQ0_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                         32'h00000040

`define CH1_DQ0_SWI_DQS_RX_PI_STA                                              'h00000814
`define CH1_DQ0_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                         0
`define CH1_DQ0_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                         1
`define CH1_DQ0_SWI_DQS_RX_PI_STA___POR                                      32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0                                      'h00000818
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1                                      'h0000081C
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0                                      'h00000820
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1                                      'h00000824
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0                                      'h00000828
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1                                      'h0000082C
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0                                      'h00000830
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1                                      'h00000834
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ0_SWI_DQS_RX_IO_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                    'h00000838
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                    23
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                   22
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                  21
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                  18:16
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                        20
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                 19
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                  7:4
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                  3:0
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                15:12
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                 11:8
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                            32'h004A7777

`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                    'h0000083C
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                    23
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                   22
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                  21
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                  18:16
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                        20
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                 19
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                  7:4
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                  3:0
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                15:12
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                 11:8
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                            32'h004A7777

`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                    'h00000840
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                    23
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                   22
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                  21
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                  18:16
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                        20
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                 19
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                  7:4
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                  3:0
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                15:12
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                 11:8
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                            32'h004A7777

`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                    'h00000844
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                    23
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                   22
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                  21
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                  18:16
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                        20
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                 19
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                  7:4
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                  3:0
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                15:12
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                 11:8
`define CH1_DQ0_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                            32'h004A7777

`define CH1_DQ0_SWI_DQS_RX_IO_STA                                              'h00000848
`define CH1_DQ0_SWI_DQS_RX_IO_STA__CORE_IG                                           31:0
`define CH1_DQ0_SWI_DQS_RX_IO_STA___POR                                      32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0                                      'h0000084C
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1                                      'h00000850
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0                                      'h00000854
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1                                      'h00000858
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0                                      'h0000085C
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1                                      'h00000860
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0                                      'h00000864
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1                                      'h00000868
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ0_SWI_DQS_RX_SA_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG                                          'h0000086C
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                           4
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                    2
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                     0
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                    3
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                     1
`define CH1_DQ0_SWI_DQS_RX_SA_CMN_CFG___POR                                  32'h00000005

`define CH1_DQ0_SWI_DQS_TX_M0_CFG                                              'h00000870
`define CH1_DQ0_SWI_DQS_TX_M0_CFG__WGB_MODE                                           7:4
`define CH1_DQ0_SWI_DQS_TX_M0_CFG__TGB_MODE                                           2:0
`define CH1_DQ0_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                       9:8
`define CH1_DQ0_SWI_DQS_TX_M0_CFG___POR                                      32'h00000087

`define CH1_DQ0_SWI_DQS_TX_M1_CFG                                              'h00000874
`define CH1_DQ0_SWI_DQS_TX_M1_CFG__WGB_MODE                                           7:4
`define CH1_DQ0_SWI_DQS_TX_M1_CFG__TGB_MODE                                           2:0
`define CH1_DQ0_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                       9:8
`define CH1_DQ0_SWI_DQS_TX_M1_CFG___POR                                      32'h00000087

`define CH1_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG                                      'h00000878
`define CH1_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                           1
`define CH1_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                           0
`define CH1_DQ0_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                              32'h00000000

`define CH1_DQ0_SWI_DQS_TX_BSCAN_CFG                                           'h0000087C
`define CH1_DQ0_SWI_DQS_TX_BSCAN_CFG__VAL                                             3:0
`define CH1_DQ0_SWI_DQS_TX_BSCAN_CFG___POR                                   32'h00000000

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                 'h00000880
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1                                 'h00000884
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2                                 'h00000888
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3                                 'h0000088C
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4                                 'h00000890
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5                                 'h00000894
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6                                 'h00000898
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7                                 'h0000089C
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8                                 'h000008A0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                 'h000008A4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1                                 'h000008A8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2                                 'h000008AC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3                                 'h000008B0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4                                 'h000008B4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5                                 'h000008B8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6                                 'h000008BC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7                                 'h000008C0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8                                 'h000008C4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                           5:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8___POR                         32'h00000001

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                 'h000008C8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1                                 'h000008CC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2                                 'h000008D0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3                                 'h000008D4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4                                 'h000008D8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5                                 'h000008DC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6                                 'h000008E0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7                                 'h000008E4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8                                 'h000008E8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                 'h000008EC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1                                 'h000008F0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2                                 'h000008F4
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3                                 'h000008F8
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4                                 'h000008FC
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5                                 'h00000900
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6                                 'h00000904
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7                                 'h00000908
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8                                 'h0000090C
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                           6:0
`define CH1_DQ0_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8___POR                         32'h00000002

`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                    'h00000910
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                    'h00000914
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                    'h00000918
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                    'h0000091C
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ0_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                  'h00000920
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                  'h00000924
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                  'h00000928
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                  'h0000092C
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                  'h00000930
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                  'h00000934
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                  'h00000938
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                  'h0000093C
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                  'h00000940
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                  'h00000944
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                  'h00000948
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                  'h0000094C
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                  'h00000950
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                  'h00000954
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                  'h00000958
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                  'h0000095C
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                      14
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ0_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG                                     'h00000960
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                         14
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG                                     'h00000964
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                         14
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG                                     'h00000968
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                         14
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG                                     'h0000096C
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                    13:10
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                      9:6
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                         14
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                      5:0
`define CH1_DQ0_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                             32'h00000040

`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                    'h00000970
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                    'h00000974
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                    'h00000978
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                    'h0000097C
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                    'h00000980
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                    'h00000984
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                    'h00000988
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                    'h0000098C
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                     5:0
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ0_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ0_SWI_DQS_TX_RT_M0_R0_CFG                                        'h00000990
`define CH1_DQ0_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                      8:0
`define CH1_DQ0_SWI_DQS_TX_RT_M0_R0_CFG___POR                                32'h00000000

`define CH1_DQ0_SWI_DQS_TX_RT_M0_R1_CFG                                        'h00000994
`define CH1_DQ0_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                      8:0
`define CH1_DQ0_SWI_DQS_TX_RT_M0_R1_CFG___POR                                32'h00000000

`define CH1_DQ0_SWI_DQS_TX_RT_M1_R0_CFG                                        'h00000998
`define CH1_DQ0_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                      8:0
`define CH1_DQ0_SWI_DQS_TX_RT_M1_R0_CFG___POR                                32'h00000000

`define CH1_DQ0_SWI_DQS_TX_RT_M1_R1_CFG                                        'h0000099C
`define CH1_DQ0_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                      8:0
`define CH1_DQ0_SWI_DQS_TX_RT_M1_R1_CFG___POR                                32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0                                     'h000009A0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1                                     'h000009A4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2                                     'h000009A8
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3                                     'h000009AC
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4                                     'h000009B0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5                                     'h000009B4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6                                     'h000009B8
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7                                     'h000009BC
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8                                     'h000009C0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0                                     'h000009C4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1                                     'h000009C8
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2                                     'h000009CC
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3                                     'h000009D0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4                                     'h000009D4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5                                     'h000009D8
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6                                     'h000009DC
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7                                     'h000009E0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8                                     'h000009E4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0                                     'h000009E8
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1                                     'h000009EC
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2                                     'h000009F0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3                                     'h000009F4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4                                     'h000009F8
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5                                     'h000009FC
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6                                     'h00000A00
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7                                     'h00000A04
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8                                     'h00000A08
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0                                     'h00000A0C
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1                                     'h00000A10
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2                                     'h00000A14
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3                                     'h00000A18
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4                                     'h00000A1C
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5                                     'h00000A20
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6                                     'h00000A24
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7                                     'h00000A28
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8                                     'h00000A2C
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_SDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                               'h00000A30
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1                               'h00000A34
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2                               'h00000A38
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3                               'h00000A3C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4                               'h00000A40
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5                               'h00000A44
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6                               'h00000A48
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7                               'h00000A4C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8                               'h00000A50
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                               'h00000A54
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1                               'h00000A58
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2                               'h00000A5C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3                               'h00000A60
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4                               'h00000A64
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5                               'h00000A68
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6                               'h00000A6C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7                               'h00000A70
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8                               'h00000A74
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                               'h00000A78
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1                               'h00000A7C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2                               'h00000A80
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3                               'h00000A84
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4                               'h00000A88
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5                               'h00000A8C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6                               'h00000A90
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7                               'h00000A94
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8                               'h00000A98
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                               'h00000A9C
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1                               'h00000AA0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2                               'h00000AA4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3                               'h00000AA8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4                               'h00000AAC
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5                               'h00000AB0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6                               'h00000AB4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7                               'h00000AB8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8                               'h00000ABC
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ0_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                              'h00000AC0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1                              'h00000AC4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2                              'h00000AC8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3                              'h00000ACC
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4                              'h00000AD0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5                              'h00000AD4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6                              'h00000AD8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7                              'h00000ADC
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8                              'h00000AE0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                              'h00000AE4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1                              'h00000AE8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2                              'h00000AEC
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3                              'h00000AF0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4                              'h00000AF4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5                              'h00000AF8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6                              'h00000AFC
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7                              'h00000B00
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8                              'h00000B04
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                              'h00000B08
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1                              'h00000B0C
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2                              'h00000B10
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3                              'h00000B14
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4                              'h00000B18
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5                              'h00000B1C
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6                              'h00000B20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7                              'h00000B24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8                              'h00000B28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                              'h00000B2C
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1                              'h00000B30
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2                              'h00000B34
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3                              'h00000B38
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4                              'h00000B3C
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5                              'h00000B40
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6                              'h00000B44
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7                              'h00000B48
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8                              'h00000B4C
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                           29:28
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                           25:24
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                           21:20
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                           17:16
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                           13:12
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                             9:8
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                             5:4
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                             1:0
`define CH1_DQ0_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                      32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0                                     'h00000B50
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1                                     'h00000B54
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2                                     'h00000B58
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3                                     'h00000B5C
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4                                     'h00000B60
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5                                     'h00000B64
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6                                     'h00000B68
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7                                     'h00000B6C
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8                                     'h00000B70
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0                                     'h00000B74
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1                                     'h00000B78
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2                                     'h00000B7C
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3                                     'h00000B80
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4                                     'h00000B84
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5                                     'h00000B88
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6                                     'h00000B8C
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7                                     'h00000B90
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8                                     'h00000B94
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0                                     'h00000B98
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1                                     'h00000B9C
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2                                     'h00000BA0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3                                     'h00000BA4
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4                                     'h00000BA8
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5                                     'h00000BAC
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6                                     'h00000BB0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7                                     'h00000BB4
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8                                     'h00000BB8
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0                                     'h00000BBC
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1                                     'h00000BC0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2                                     'h00000BC4
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3                                     'h00000BC8
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4                                     'h00000BCC
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5                                     'h00000BD0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6                                     'h00000BD4
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7                                     'h00000BD8
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8                                     'h00000BDC
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_DDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                               'h00000BE0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1                               'h00000BE4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2                               'h00000BE8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3                               'h00000BEC
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4                               'h00000BF0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5                               'h00000BF4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6                               'h00000BF8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7                               'h00000BFC
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8                               'h00000C00
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                               'h00000C04
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1                               'h00000C08
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2                               'h00000C0C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3                               'h00000C10
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4                               'h00000C14
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5                               'h00000C18
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6                               'h00000C1C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7                               'h00000C20
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8                               'h00000C24
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                               'h00000C28
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1                               'h00000C2C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2                               'h00000C30
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3                               'h00000C34
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4                               'h00000C38
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5                               'h00000C3C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6                               'h00000C40
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7                               'h00000C44
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8                               'h00000C48
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                               'h00000C4C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1                               'h00000C50
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2                               'h00000C54
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3                               'h00000C58
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4                               'h00000C5C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5                               'h00000C60
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6                               'h00000C64
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7                               'h00000C68
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8                               'h00000C6C
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ0_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0                                     'h00000C70
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1                                     'h00000C74
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2                                     'h00000C78
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3                                     'h00000C7C
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4                                     'h00000C80
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5                                     'h00000C84
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6                                     'h00000C88
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7                                     'h00000C8C
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8                                     'h00000C90
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0                                     'h00000C94
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1                                     'h00000C98
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2                                     'h00000C9C
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3                                     'h00000CA0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4                                     'h00000CA4
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5                                     'h00000CA8
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6                                     'h00000CAC
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7                                     'h00000CB0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8                                     'h00000CB4
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0                                     'h00000CB8
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1                                     'h00000CBC
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2                                     'h00000CC0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3                                     'h00000CC4
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4                                     'h00000CC8
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5                                     'h00000CCC
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6                                     'h00000CD0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7                                     'h00000CD4
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8                                     'h00000CD8
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0                                     'h00000CDC
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1                                     'h00000CE0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2                                     'h00000CE4
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3                                     'h00000CE8
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4                                     'h00000CEC
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5                                     'h00000CF0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6                                     'h00000CF4
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7                                     'h00000CF8
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8                                     'h00000CFC
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ0_SWI_DQS_TX_QDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                               'h00000D00
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1                               'h00000D04
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2                               'h00000D08
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3                               'h00000D0C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4                               'h00000D10
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5                               'h00000D14
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6                               'h00000D18
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7                               'h00000D1C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8                               'h00000D20
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                               'h00000D24
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1                               'h00000D28
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2                               'h00000D2C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3                               'h00000D30
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4                               'h00000D34
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5                               'h00000D38
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6                               'h00000D3C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7                               'h00000D40
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8                               'h00000D44
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                               'h00000D48
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1                               'h00000D4C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2                               'h00000D50
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3                               'h00000D54
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4                               'h00000D58
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5                               'h00000D5C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6                               'h00000D60
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7                               'h00000D64
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8                               'h00000D68
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                               'h00000D6C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1                               'h00000D70
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2                               'h00000D74
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3                               'h00000D78
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4                               'h00000D7C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5                               'h00000D80
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6                               'h00000D84
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7                               'h00000D88
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8                               'h00000D8C
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              4
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              0
`define CH1_DQ0_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                    'h00000D90
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1                                    'h00000D94
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R0_CFG_1___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                    'h00000D98
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1                                    'h00000D9C
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M0_R1_CFG_1___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                    'h00000DA0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1                                    'h00000DA4
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R0_CFG_1___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                    'h00000DA8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1                                    'h00000DAC
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__GEAR                                     7:6
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__EN                                         8
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ0_SWI_DQS_TX_LPDE_M1_R1_CFG_1___POR                            32'h00000100

`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0                                         'h00000DB0
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                       8:6
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                          5
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                      11:9
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                      4
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                      3
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                      2:0
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_0___POR                                 32'h00000041

`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1                                         'h00000DB4
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__TX_IMPD                                       8:6
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__SW_OVR                                          5
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__RX_IMPD                                      11:9
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_T                                      4
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_C                                      3
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1__OVRD_SEL                                      2:0
`define CH1_DQ0_SWI_DQS_TX_IO_M0_CFG_1___POR                                 32'h00000041

`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0                                         'h00000DB8
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                       8:6
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                          5
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                      11:9
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                      4
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                      3
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                      2:0
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_0___POR                                 32'h00000041

`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1                                         'h00000DBC
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__TX_IMPD                                       8:6
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__SW_OVR                                          5
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__RX_IMPD                                      11:9
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_T                                      4
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_C                                      3
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1__OVRD_SEL                                      2:0
`define CH1_DQ0_SWI_DQS_TX_IO_M1_CFG_1___POR                                 32'h00000041

`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                    'h00000DC0
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                   13
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                    10:5
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                     4:0
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                   12
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                     11
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                            32'h00000001

`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                    'h00000DC4
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                   13
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                    10:5
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                     4:0
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                   12
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                     11
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                            32'h00000001

`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                    'h00000DC8
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                   13
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                    10:5
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                     4:0
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                   12
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                     11
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                            32'h00000001

`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                    'h00000DCC
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                   13
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                    10:5
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                     4:0
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                   12
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                     11
`define CH1_DQ0_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                            32'h00000001

`define CH1_DQ1_SWI_TOP_CFG                                                    'h00000000
`define CH1_DQ1_SWI_TOP_CFG__WCS_SW_OVR_VAL                                             1
`define CH1_DQ1_SWI_TOP_CFG__WCS_SW_OVR                                                 0
`define CH1_DQ1_SWI_TOP_CFG__TRAINING_MODE                                              9
`define CH1_DQ1_SWI_TOP_CFG__RCS_SW_OVR_VAL                                             3
`define CH1_DQ1_SWI_TOP_CFG__RCS_SW_OVR                                                 2
`define CH1_DQ1_SWI_TOP_CFG__FIFO_CLR                                                   8
`define CH1_DQ1_SWI_TOP_CFG___POR                                            32'h00000000

`define CH1_DQ1_SWI_TOP_STA                                                    'h00000004
`define CH1_DQ1_SWI_TOP_STA__WCS                                                        0
`define CH1_DQ1_SWI_TOP_STA__RCS                                                        1
`define CH1_DQ1_SWI_TOP_STA___POR                                            32'h00000000

`define CH1_DQ1_SWI_DQ_RX_BSCAN_STA                                            'h00000008
`define CH1_DQ1_SWI_DQ_RX_BSCAN_STA__VAL                                              8:0
`define CH1_DQ1_SWI_DQ_RX_BSCAN_STA___POR                                    32'h00000000

`define CH1_DQ1_SWI_DQ_RX_M0_CFG                                               'h0000000C
`define CH1_DQ1_SWI_DQ_RX_M0_CFG__RGB_MODE                                            2:0
`define CH1_DQ1_SWI_DQ_RX_M0_CFG__FGB_MODE                                            7:4
`define CH1_DQ1_SWI_DQ_RX_M0_CFG___POR                                       32'h00000074

`define CH1_DQ1_SWI_DQ_RX_M1_CFG                                               'h00000010
`define CH1_DQ1_SWI_DQ_RX_M1_CFG__RGB_MODE                                            2:0
`define CH1_DQ1_SWI_DQ_RX_M1_CFG__FGB_MODE                                            7:4
`define CH1_DQ1_SWI_DQ_RX_M1_CFG___POR                                       32'h00000074

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0                                       'h00000014
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1                                       'h00000018
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2                                       'h0000001C
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3                                       'h00000020
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4                                       'h00000024
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5                                       'h00000028
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6                                       'h0000002C
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7                                       'h00000030
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8                                       'h00000034
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0                                       'h00000038
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1                                       'h0000003C
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2                                       'h00000040
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3                                       'h00000044
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4                                       'h00000048
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5                                       'h0000004C
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6                                       'h00000050
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7                                       'h00000054
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8                                       'h00000058
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0                                       'h0000005C
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1                                       'h00000060
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2                                       'h00000064
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3                                       'h00000068
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4                                       'h0000006C
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5                                       'h00000070
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6                                       'h00000074
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7                                       'h00000078
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8                                       'h0000007C
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0                                       'h00000080
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1                                       'h00000084
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2                                       'h00000088
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3                                       'h0000008C
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4                                       'h00000090
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5                                       'h00000094
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6                                       'h00000098
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7                                       'h0000009C
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8                                       'h000000A0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                   7:0
`define CH1_DQ1_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_IO_STA                                               'h000000A4
`define CH1_DQ1_SWI_DQ_RX_IO_STA__CORE_IG                                            31:0
`define CH1_DQ1_SWI_DQ_RX_IO_STA___POR                                       32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0                                       'h000000A8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1                                       'h000000AC
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2                                       'h000000B0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3                                       'h000000B4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4                                       'h000000B8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5                                       'h000000BC
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6                                       'h000000C0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7                                       'h000000C4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8                                       'h000000C8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0                                       'h000000CC
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1                                       'h000000D0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2                                       'h000000D4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3                                       'h000000D8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4                                       'h000000DC
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5                                       'h000000E0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6                                       'h000000E4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7                                       'h000000E8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8                                       'h000000EC
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0                                       'h000000F0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1                                       'h000000F4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2                                       'h000000F8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3                                       'h000000FC
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4                                       'h00000100
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5                                       'h00000104
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6                                       'h00000108
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7                                       'h0000010C
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8                                       'h00000110
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0                                       'h00000114
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1                                       'h00000118
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2                                       'h0000011C
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3                                       'h00000120
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4                                       'h00000124
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5                                       'h00000128
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6                                       'h0000012C
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7                                       'h00000130
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8                                       'h00000134
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                   17
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                  19
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                  18
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                    16
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                 7:4
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                              15:12
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                               11:8
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                  3:0
`define CH1_DQ1_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                   'h00000138
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                   'h0000013C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                   'h00000140
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                   'h00000144
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                   'h00000148
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                   'h0000014C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                   'h00000150
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                   'h00000154
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                   'h00000158
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                   'h0000015C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                   'h00000160
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                   'h00000164
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                   'h00000168
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                   'h0000016C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                   'h00000170
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                   'h00000174
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                   'h00000178
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                   'h0000017C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                   'h00000180
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                   'h00000184
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                   'h00000188
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                   'h0000018C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                   'h00000190
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                   'h00000194
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                   'h00000198
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                   'h0000019C
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                   'h000001A0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                   'h000001A4
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                   'h000001A8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                   'h000001AC
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                   'h000001B0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                   'h000001B4
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                   'h000001B8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                   'h000001BC
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                   'h000001C0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                   'h000001C4
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                 9:8
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                              25:24
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                              17:16
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                  1:0
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                               15:10
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                              31:26
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                              23:18
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                  7:2
`define CH1_DQ1_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                           32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_0                                             'h000001C8
`define CH1_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_0___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_1                                             'h000001CC
`define CH1_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_1___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_2                                             'h000001D0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_2___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_3                                             'h000001D4
`define CH1_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_3___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_4                                             'h000001D8
`define CH1_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_4___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_5                                             'h000001DC
`define CH1_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_5___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_6                                             'h000001E0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_6___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_7                                             'h000001E4
`define CH1_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_7___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_RX_SA_STA_8                                             'h000001E8
`define CH1_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                           1
`define CH1_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                          3
`define CH1_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                          2
`define CH1_DQ1_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                            0
`define CH1_DQ1_SWI_DQ_RX_SA_STA_8___POR                                     32'h00000000

`define CH1_DQ1_SWI_DQ_TX_BSCAN_CFG                                            'h000001EC
`define CH1_DQ1_SWI_DQ_TX_BSCAN_CFG__VAL                                              8:0
`define CH1_DQ1_SWI_DQ_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                  'h000001F0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                  'h000001F4
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                  'h000001F8
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                  'h000001FC
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                  'h00000200
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                  'h00000204
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                  'h00000208
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                  'h0000020C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                  'h00000210
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                  'h00000214
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                  'h00000218
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                  'h0000021C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                  'h00000220
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                  'h00000224
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                  'h00000228
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                  'h0000022C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                  'h00000230
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                  'h00000234
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                            5:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                          32'h00000001

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                  'h00000238
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                  'h0000023C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                  'h00000240
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                  'h00000244
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                  'h00000248
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                  'h0000024C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                  'h00000250
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                  'h00000254
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                  'h00000258
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                  'h0000025C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                  'h00000260
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                  'h00000264
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                  'h00000268
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                  'h0000026C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                  'h00000270
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                  'h00000274
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                  'h00000278
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                  'h0000027C
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                            6:0
`define CH1_DQ1_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                          32'h00000002

`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                     'h00000280
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                     'h00000284
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                     'h00000288
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                     'h0000028C
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                   'h00000290
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                   'h00000294
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                   'h00000298
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                   'h0000029C
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                   'h000002A0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                   'h000002A4
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                   'h000002A8
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                   'h000002AC
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                   'h000002B0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                   'h000002B4
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                   'h000002B8
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                   'h000002BC
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                   'h000002C0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                   'h000002C4
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                   'h000002C8
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                   'h000002CC
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_DQ1_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG                                      'h000002D0
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG                                      'h000002D4
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG                                      'h000002D8
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG                                      'h000002DC
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH1_DQ1_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH1_DQ1_SWI_DQ_TX_RT_M0_R0_CFG                                         'h000002E0
`define CH1_DQ1_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       8:0
`define CH1_DQ1_SWI_DQ_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH1_DQ1_SWI_DQ_TX_RT_M0_R1_CFG                                         'h000002E4
`define CH1_DQ1_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       8:0
`define CH1_DQ1_SWI_DQ_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH1_DQ1_SWI_DQ_TX_RT_M1_R0_CFG                                         'h000002E8
`define CH1_DQ1_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       8:0
`define CH1_DQ1_SWI_DQ_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH1_DQ1_SWI_DQ_TX_RT_M1_R1_CFG                                         'h000002EC
`define CH1_DQ1_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       8:0
`define CH1_DQ1_SWI_DQ_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0                                      'h000002F0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1                                      'h000002F4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2                                      'h000002F8
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3                                      'h000002FC
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4                                      'h00000300
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5                                      'h00000304
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6                                      'h00000308
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7                                      'h0000030C
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8                                      'h00000310
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0                                      'h00000314
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1                                      'h00000318
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2                                      'h0000031C
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3                                      'h00000320
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4                                      'h00000324
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5                                      'h00000328
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6                                      'h0000032C
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7                                      'h00000330
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8                                      'h00000334
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0                                      'h00000338
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1                                      'h0000033C
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2                                      'h00000340
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3                                      'h00000344
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4                                      'h00000348
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5                                      'h0000034C
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6                                      'h00000350
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7                                      'h00000354
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8                                      'h00000358
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0                                      'h0000035C
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1                                      'h00000360
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2                                      'h00000364
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3                                      'h00000368
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4                                      'h0000036C
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5                                      'h00000370
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6                                      'h00000374
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7                                      'h00000378
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8                                      'h0000037C
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                   7
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                   6
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                   5
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                   4
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000380
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                'h00000384
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                'h00000388
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                'h0000038C
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                'h00000390
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                'h00000394
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                'h00000398
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                'h0000039C
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                'h000003A0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                'h000003A4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                'h000003A8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                'h000003AC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                'h000003B0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                'h000003B4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                'h000003B8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                'h000003BC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                'h000003C0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                'h000003C4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                'h000003C8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                'h000003CC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                'h000003D0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                'h000003D4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                'h000003D8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                'h000003DC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                'h000003E0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                'h000003E4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                'h000003E8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                'h000003EC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                'h000003F0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                'h000003F4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                'h000003F8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                'h000003FC
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                'h00000400
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                'h00000404
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                'h00000408
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                'h0000040C
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                           30:28
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                           26:24
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                           22:20
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                           18:16
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           14:12
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            10:8
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             6:4
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             2:0
`define CH1_DQ1_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000410
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                               'h00000414
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                               'h00000418
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                               'h0000041C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                               'h00000420
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                               'h00000424
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                               'h00000428
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                               'h0000042C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                               'h00000430
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000434
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                               'h00000438
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                               'h0000043C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                               'h00000440
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                               'h00000444
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                               'h00000448
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                               'h0000044C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                               'h00000450
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                               'h00000454
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000458
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                               'h0000045C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                               'h00000460
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                               'h00000464
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                               'h00000468
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                               'h0000046C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                               'h00000470
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                               'h00000474
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                               'h00000478
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h0000047C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                               'h00000480
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                               'h00000484
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                               'h00000488
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                               'h0000048C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                               'h00000490
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                               'h00000494
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                               'h00000498
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                               'h0000049C
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                            29:28
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                            25:24
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                            21:20
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                            17:16
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                            13:12
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                              9:8
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                              5:4
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                              1:0
`define CH1_DQ1_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0                                      'h000004A0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1                                      'h000004A4
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2                                      'h000004A8
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3                                      'h000004AC
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4                                      'h000004B0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5                                      'h000004B4
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6                                      'h000004B8
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7                                      'h000004BC
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8                                      'h000004C0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0                                      'h000004C4
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1                                      'h000004C8
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2                                      'h000004CC
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3                                      'h000004D0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4                                      'h000004D4
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5                                      'h000004D8
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6                                      'h000004DC
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7                                      'h000004E0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8                                      'h000004E4
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0                                      'h000004E8
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1                                      'h000004EC
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2                                      'h000004F0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3                                      'h000004F4
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4                                      'h000004F8
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5                                      'h000004FC
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6                                      'h00000500
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7                                      'h00000504
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8                                      'h00000508
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0                                      'h0000050C
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1                                      'h00000510
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2                                      'h00000514
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3                                      'h00000518
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4                                      'h0000051C
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5                                      'h00000520
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6                                      'h00000524
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7                                      'h00000528
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8                                      'h0000052C
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                   3
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                   2
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000530
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                'h00000534
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                'h00000538
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                'h0000053C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                'h00000540
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                'h00000544
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                'h00000548
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                'h0000054C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                'h00000550
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000554
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                'h00000558
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                'h0000055C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                'h00000560
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                'h00000564
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                'h00000568
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                'h0000056C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                'h00000570
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                'h00000574
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000578
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                'h0000057C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                'h00000580
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                'h00000584
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                'h00000588
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                'h0000058C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                'h00000590
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                'h00000594
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                'h00000598
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                'h0000059C
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                'h000005A0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                'h000005A4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                'h000005A8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                'h000005AC
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                'h000005B0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                'h000005B4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                'h000005B8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                'h000005BC
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                           13:12
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             9:8
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                             5:4
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                             1:0
`define CH1_DQ1_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0                                      'h000005C0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1                                      'h000005C4
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2                                      'h000005C8
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3                                      'h000005CC
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4                                      'h000005D0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5                                      'h000005D4
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6                                      'h000005D8
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7                                      'h000005DC
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8                                      'h000005E0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0                                      'h000005E4
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1                                      'h000005E8
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2                                      'h000005EC
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3                                      'h000005F0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4                                      'h000005F4
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5                                      'h000005F8
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6                                      'h000005FC
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7                                      'h00000600
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8                                      'h00000604
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0                                      'h00000608
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1                                      'h0000060C
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2                                      'h00000610
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3                                      'h00000614
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4                                      'h00000618
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5                                      'h0000061C
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6                                      'h00000620
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7                                      'h00000624
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8                                      'h00000628
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0                                      'h0000062C
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1                                      'h00000630
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2                                      'h00000634
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3                                      'h00000638
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4                                      'h0000063C
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5                                      'h00000640
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6                                      'h00000644
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7                                      'h00000648
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8                                      'h0000064C
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                   1
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                   0
`define CH1_DQ1_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                              32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000650
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                'h00000654
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                'h00000658
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                'h0000065C
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                'h00000660
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                'h00000664
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                'h00000668
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                'h0000066C
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                'h00000670
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000674
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                'h00000678
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                'h0000067C
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                'h00000680
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                'h00000684
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                'h00000688
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                'h0000068C
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                'h00000690
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                'h00000694
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000698
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                'h0000069C
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                'h000006A0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                'h000006A4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                'h000006A8
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                'h000006AC
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                'h000006B0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                'h000006B4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                'h000006B8
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                'h000006BC
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                'h000006C0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                'h000006C4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                'h000006C8
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                'h000006CC
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                'h000006D0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                'h000006D4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                'h000006D8
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                'h000006DC
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                               4
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                               0
`define CH1_DQ1_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                     'h000006E0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                     'h000006E4
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                     'h000006E8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                     'h000006EC
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                     'h000006F0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                     'h000006F4
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                     'h000006F8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                     'h000006FC
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                     'h00000700
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                     'h00000704
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                     'h00000708
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                     'h0000070C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                     'h00000710
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                     'h00000714
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                     'h00000718
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                     'h0000071C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                     'h00000720
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                     'h00000724
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                     'h00000728
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                     'h0000072C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                     'h00000730
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                     'h00000734
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                     'h00000738
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                     'h0000073C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                     'h00000740
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                     'h00000744
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                     'h00000748
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                     'h0000074C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                     'h00000750
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                     'h00000754
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                     'h00000758
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                     'h0000075C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                     'h00000760
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                     'h00000764
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                     'h00000768
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                     'h0000076C
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                      7:6
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                          8
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                  5:0
`define CH1_DQ1_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                             32'h00000100

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0                                          'h00000770
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_0___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1                                          'h00000774
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_1___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2                                          'h00000778
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_2___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3                                          'h0000077C
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_3___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4                                          'h00000780
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_4___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5                                          'h00000784
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_5___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6                                          'h00000788
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_6___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7                                          'h0000078C
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_7___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8                                          'h00000790
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M0_CFG_8___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0                                          'h00000794
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_0___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1                                          'h00000798
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_1___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2                                          'h0000079C
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_2___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3                                          'h000007A0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_3___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4                                          'h000007A4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_4___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5                                          'h000007A8
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_5___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6                                          'h000007AC
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_6___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7                                          'h000007B0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_7___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8                                          'h000007B4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                        8:6
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                           5
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                       11:9
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                        4
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                         3
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                       2:0
`define CH1_DQ1_SWI_DQ_TX_IO_M1_CFG_8___POR                                  32'h00000040

`define CH1_DQ1_SWI_DQS_RX_M0_CFG                                              'h000007B8
`define CH1_DQ1_SWI_DQS_RX_M0_CFG__WCK_MODE                                             8
`define CH1_DQ1_SWI_DQS_RX_M0_CFG__RGB_MODE                                           2:0
`define CH1_DQ1_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                   13:12
`define CH1_DQ1_SWI_DQS_RX_M0_CFG__FGB_MODE                                           7:4
`define CH1_DQ1_SWI_DQS_RX_M0_CFG___POR                                      32'h00000074

`define CH1_DQ1_SWI_DQS_RX_M1_CFG                                              'h000007BC
`define CH1_DQ1_SWI_DQS_RX_M1_CFG__WCK_MODE                                             8
`define CH1_DQ1_SWI_DQS_RX_M1_CFG__RGB_MODE                                           2:0
`define CH1_DQ1_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                   13:12
`define CH1_DQ1_SWI_DQS_RX_M1_CFG__FGB_MODE                                           7:4
`define CH1_DQ1_SWI_DQS_RX_M1_CFG___POR                                      32'h00000074

`define CH1_DQ1_SWI_DQS_RX_BSCAN_STA                                           'h000007C0
`define CH1_DQ1_SWI_DQS_RX_BSCAN_STA__VAL                                             3:0
`define CH1_DQ1_SWI_DQS_RX_BSCAN_STA___POR                                   32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                  'h000007C4
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                   7:6
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                       8
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                               5:0
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                          32'h00000100

`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                  'h000007C8
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                   7:6
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                       8
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                               5:0
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                          32'h00000100

`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                  'h000007CC
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                   7:6
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                       8
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                               5:0
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                          32'h00000100

`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                  'h000007D0
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                   7:6
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                       8
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                               5:0
`define CH1_DQ1_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                          32'h00000100

`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG                                    'h000007D4
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG                                    'h000007D8
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG                                    'h000007DC
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG                                    'h000007E0
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                    'h000007E4
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                    'h000007E8
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                    'h000007EC
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                    'h000007F0
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                 'h000007F4
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                 'h000007F8
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                 'h000007FC
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                 'h00000800
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                 'h00000804
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                 'h00000808
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                 'h0000080C
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                 'h00000810
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                13:10
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                  9:6
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                     14
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                  5:0
`define CH1_DQ1_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                         32'h00000040

`define CH1_DQ1_SWI_DQS_RX_PI_STA                                              'h00000814
`define CH1_DQ1_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                         0
`define CH1_DQ1_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                         1
`define CH1_DQ1_SWI_DQS_RX_PI_STA___POR                                      32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0                                      'h00000818
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1                                      'h0000081C
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0                                      'h00000820
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1                                      'h00000824
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0                                      'h00000828
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1                                      'h0000082C
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0                                      'h00000830
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1                                      'h00000834
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_T                                15:8
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1__DLY_CTRL_C                                 7:0
`define CH1_DQ1_SWI_DQS_RX_IO_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                    'h00000838
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                    23
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                   22
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                  21
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                  18:16
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                        20
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                 19
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                  7:4
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                  3:0
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                15:12
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                 11:8
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                            32'h004A7777

`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                    'h0000083C
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                    23
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                   22
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                  21
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                  18:16
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                        20
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                 19
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                  7:4
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                  3:0
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                15:12
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                 11:8
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                            32'h004A7777

`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                    'h00000840
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                    23
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                   22
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                  21
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                  18:16
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                        20
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                 19
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                  7:4
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                  3:0
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                15:12
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                 11:8
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                            32'h004A7777

`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                    'h00000844
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                    23
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                   22
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                  21
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                  18:16
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                        20
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                 19
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                  7:4
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                  3:0
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                15:12
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                 11:8
`define CH1_DQ1_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                            32'h004A7777

`define CH1_DQ1_SWI_DQS_RX_IO_STA                                              'h00000848
`define CH1_DQ1_SWI_DQS_RX_IO_STA__CORE_IG                                           31:0
`define CH1_DQ1_SWI_DQS_RX_IO_STA___POR                                      32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0                                      'h0000084C
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1                                      'h00000850
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0                                      'h00000854
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1                                      'h00000858
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M0_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0                                      'h0000085C
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1                                      'h00000860
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R0_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0                                      'h00000864
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1                                      'h00000868
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                  17
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                 19
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                 18
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                   16
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                7:4
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_270                             15:12
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_180                              11:8
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                 3:0
`define CH1_DQ1_SWI_DQS_RX_SA_M1_R1_CFG_1___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG                                          'h0000086C
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                           4
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                    2
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                     0
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                    3
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                     1
`define CH1_DQ1_SWI_DQS_RX_SA_CMN_CFG___POR                                  32'h00000005

`define CH1_DQ1_SWI_DQS_TX_M0_CFG                                              'h00000870
`define CH1_DQ1_SWI_DQS_TX_M0_CFG__WGB_MODE                                           7:4
`define CH1_DQ1_SWI_DQS_TX_M0_CFG__TGB_MODE                                           2:0
`define CH1_DQ1_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                       9:8
`define CH1_DQ1_SWI_DQS_TX_M0_CFG___POR                                      32'h00000087

`define CH1_DQ1_SWI_DQS_TX_M1_CFG                                              'h00000874
`define CH1_DQ1_SWI_DQS_TX_M1_CFG__WGB_MODE                                           7:4
`define CH1_DQ1_SWI_DQS_TX_M1_CFG__TGB_MODE                                           2:0
`define CH1_DQ1_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                       9:8
`define CH1_DQ1_SWI_DQS_TX_M1_CFG___POR                                      32'h00000087

`define CH1_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG                                      'h00000878
`define CH1_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                           1
`define CH1_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                           0
`define CH1_DQ1_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                              32'h00000000

`define CH1_DQ1_SWI_DQS_TX_BSCAN_CFG                                           'h0000087C
`define CH1_DQ1_SWI_DQS_TX_BSCAN_CFG__VAL                                             3:0
`define CH1_DQ1_SWI_DQS_TX_BSCAN_CFG___POR                                   32'h00000000

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                 'h00000880
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1                                 'h00000884
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_1___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2                                 'h00000888
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_2___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3                                 'h0000088C
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_3___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4                                 'h00000890
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_4___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5                                 'h00000894
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_5___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6                                 'h00000898
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_6___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7                                 'h0000089C
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_7___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8                                 'h000008A0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M0_CFG_8___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                 'h000008A4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1                                 'h000008A8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_1___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2                                 'h000008AC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_2___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3                                 'h000008B0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_3___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4                                 'h000008B4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_4___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5                                 'h000008B8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_5___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6                                 'h000008BC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_6___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7                                 'h000008C0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_7___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8                                 'h000008C4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                           5:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_ANA_M1_CFG_8___POR                         32'h00000001

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                 'h000008C8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1                                 'h000008CC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_1___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2                                 'h000008D0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_2___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3                                 'h000008D4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_3___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4                                 'h000008D8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_4___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5                                 'h000008DC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_5___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6                                 'h000008E0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_6___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7                                 'h000008E4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_7___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8                                 'h000008E8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M0_CFG_8___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                 'h000008EC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1                                 'h000008F0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_1___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2                                 'h000008F4
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_2___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3                                 'h000008F8
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_3___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4                                 'h000008FC
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_4___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5                                 'h00000900
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_5___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6                                 'h00000904
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_6___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7                                 'h00000908
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_7___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8                                 'h0000090C
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                           6:0
`define CH1_DQ1_SWI_DQS_TX_EGRESS_DIG_M1_CFG_8___POR                         32'h00000002

`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                    'h00000910
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                    'h00000914
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                    'h00000918
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                    'h0000091C
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                     5:0
`define CH1_DQ1_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                  'h00000920
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                  'h00000924
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                  'h00000928
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                  'h0000092C
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                  'h00000930
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                  'h00000934
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                  'h00000938
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                  'h0000093C
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                  'h00000940
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                  'h00000944
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                  'h00000948
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                  'h0000094C
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                  'h00000950
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                  'h00000954
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                  'h00000958
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                  'h0000095C
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                      14
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH1_DQ1_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG                                     'h00000960
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                         14
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG                                     'h00000964
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                         14
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG                                     'h00000968
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                         14
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG                                     'h0000096C
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                    13:10
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                      9:6
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                         14
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                      5:0
`define CH1_DQ1_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                             32'h00000040

`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                    'h00000970
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                    'h00000974
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                    'h00000978
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                    'h0000097C
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                    'h00000980
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                    'h00000984
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                    'h00000988
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                    'h0000098C
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                   13:10
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                     5:0
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                     9:6
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                        14
`define CH1_DQ1_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                            32'h00000040

`define CH1_DQ1_SWI_DQS_TX_RT_M0_R0_CFG                                        'h00000990
`define CH1_DQ1_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                      8:0
`define CH1_DQ1_SWI_DQS_TX_RT_M0_R0_CFG___POR                                32'h00000000

`define CH1_DQ1_SWI_DQS_TX_RT_M0_R1_CFG                                        'h00000994
`define CH1_DQ1_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                      8:0
`define CH1_DQ1_SWI_DQS_TX_RT_M0_R1_CFG___POR                                32'h00000000

`define CH1_DQ1_SWI_DQS_TX_RT_M1_R0_CFG                                        'h00000998
`define CH1_DQ1_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                      8:0
`define CH1_DQ1_SWI_DQS_TX_RT_M1_R0_CFG___POR                                32'h00000000

`define CH1_DQ1_SWI_DQS_TX_RT_M1_R1_CFG                                        'h0000099C
`define CH1_DQ1_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                      8:0
`define CH1_DQ1_SWI_DQS_TX_RT_M1_R1_CFG___POR                                32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0                                     'h000009A0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1                                     'h000009A4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2                                     'h000009A8
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3                                     'h000009AC
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4                                     'h000009B0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5                                     'h000009B4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6                                     'h000009B8
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7                                     'h000009BC
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8                                     'h000009C0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0                                     'h000009C4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1                                     'h000009C8
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2                                     'h000009CC
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3                                     'h000009D0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4                                     'h000009D4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5                                     'h000009D8
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6                                     'h000009DC
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7                                     'h000009E0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8                                     'h000009E4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0                                     'h000009E8
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1                                     'h000009EC
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2                                     'h000009F0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3                                     'h000009F4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4                                     'h000009F8
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5                                     'h000009FC
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6                                     'h00000A00
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7                                     'h00000A04
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8                                     'h00000A08
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0                                     'h00000A0C
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1                                     'h00000A10
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2                                     'h00000A14
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3                                     'h00000A18
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4                                     'h00000A1C
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5                                     'h00000A20
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6                                     'h00000A24
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7                                     'h00000A28
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8                                     'h00000A2C
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                  7
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                  6
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                  5
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                  4
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_SDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                               'h00000A30
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1                               'h00000A34
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2                               'h00000A38
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3                               'h00000A3C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4                               'h00000A40
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5                               'h00000A44
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6                               'h00000A48
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7                               'h00000A4C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8                               'h00000A50
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                               'h00000A54
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1                               'h00000A58
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2                               'h00000A5C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3                               'h00000A60
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4                               'h00000A64
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5                               'h00000A68
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6                               'h00000A6C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7                               'h00000A70
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8                               'h00000A74
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                               'h00000A78
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1                               'h00000A7C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2                               'h00000A80
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3                               'h00000A84
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4                               'h00000A88
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5                               'h00000A8C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6                               'h00000A90
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7                               'h00000A94
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8                               'h00000A98
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                               'h00000A9C
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1                               'h00000AA0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2                               'h00000AA4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3                               'h00000AA8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4                               'h00000AAC
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5                               'h00000AB0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6                               'h00000AB4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7                               'h00000AB8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8                               'h00000ABC
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                          30:28
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                          26:24
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                          22:20
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                          18:16
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          14:12
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                           10:8
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            6:4
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            2:0
`define CH1_DQ1_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                              'h00000AC0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1                              'h00000AC4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2                              'h00000AC8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3                              'h00000ACC
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4                              'h00000AD0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5                              'h00000AD4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6                              'h00000AD8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7                              'h00000ADC
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8                              'h00000AE0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                              'h00000AE4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1                              'h00000AE8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2                              'h00000AEC
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3                              'h00000AF0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4                              'h00000AF4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5                              'h00000AF8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6                              'h00000AFC
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7                              'h00000B00
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8                              'h00000B04
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                              'h00000B08
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1                              'h00000B0C
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2                              'h00000B10
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3                              'h00000B14
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4                              'h00000B18
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5                              'h00000B1C
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6                              'h00000B20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7                              'h00000B24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8                              'h00000B28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                              'h00000B2C
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1                              'h00000B30
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2                              'h00000B34
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3                              'h00000B38
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4                              'h00000B3C
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5                              'h00000B40
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6                              'h00000B44
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7                              'h00000B48
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8                              'h00000B4C
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                           29:28
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                           25:24
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                           21:20
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                           17:16
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                           13:12
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                             9:8
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                             5:4
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                             1:0
`define CH1_DQ1_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                      32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0                                     'h00000B50
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1                                     'h00000B54
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2                                     'h00000B58
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3                                     'h00000B5C
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4                                     'h00000B60
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5                                     'h00000B64
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6                                     'h00000B68
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7                                     'h00000B6C
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8                                     'h00000B70
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0                                     'h00000B74
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1                                     'h00000B78
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2                                     'h00000B7C
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3                                     'h00000B80
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4                                     'h00000B84
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5                                     'h00000B88
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6                                     'h00000B8C
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7                                     'h00000B90
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8                                     'h00000B94
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0                                     'h00000B98
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1                                     'h00000B9C
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2                                     'h00000BA0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3                                     'h00000BA4
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4                                     'h00000BA8
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5                                     'h00000BAC
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6                                     'h00000BB0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7                                     'h00000BB4
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8                                     'h00000BB8
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0                                     'h00000BBC
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1                                     'h00000BC0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2                                     'h00000BC4
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3                                     'h00000BC8
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4                                     'h00000BCC
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5                                     'h00000BD0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6                                     'h00000BD4
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7                                     'h00000BD8
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8                                     'h00000BDC
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                  3
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                  2
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_DDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                               'h00000BE0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1                               'h00000BE4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2                               'h00000BE8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3                               'h00000BEC
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4                               'h00000BF0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5                               'h00000BF4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6                               'h00000BF8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7                               'h00000BFC
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8                               'h00000C00
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                               'h00000C04
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1                               'h00000C08
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2                               'h00000C0C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3                               'h00000C10
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4                               'h00000C14
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5                               'h00000C18
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6                               'h00000C1C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7                               'h00000C20
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8                               'h00000C24
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                               'h00000C28
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1                               'h00000C2C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2                               'h00000C30
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3                               'h00000C34
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4                               'h00000C38
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5                               'h00000C3C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6                               'h00000C40
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7                               'h00000C44
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8                               'h00000C48
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                               'h00000C4C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1                               'h00000C50
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2                               'h00000C54
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3                               'h00000C58
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4                               'h00000C5C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5                               'h00000C60
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6                               'h00000C64
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7                               'h00000C68
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8                               'h00000C6C
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                          13:12
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                            9:8
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                            5:4
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                            1:0
`define CH1_DQ1_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0                                     'h00000C70
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1                                     'h00000C74
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2                                     'h00000C78
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3                                     'h00000C7C
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4                                     'h00000C80
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5                                     'h00000C84
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6                                     'h00000C88
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7                                     'h00000C8C
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8                                     'h00000C90
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0                                     'h00000C94
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1                                     'h00000C98
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2                                     'h00000C9C
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3                                     'h00000CA0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4                                     'h00000CA4
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5                                     'h00000CA8
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6                                     'h00000CAC
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7                                     'h00000CB0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8                                     'h00000CB4
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M0_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0                                     'h00000CB8
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1                                     'h00000CBC
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2                                     'h00000CC0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3                                     'h00000CC4
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4                                     'h00000CC8
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5                                     'h00000CCC
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6                                     'h00000CD0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7                                     'h00000CD4
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8                                     'h00000CD8
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R0_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0                                     'h00000CDC
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1                                     'h00000CE0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_1___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2                                     'h00000CE4
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_2___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3                                     'h00000CE8
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_3___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4                                     'h00000CEC
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_4___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5                                     'h00000CF0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_5___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6                                     'h00000CF4
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_6___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7                                     'h00000CF8
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_7___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8                                     'h00000CFC
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                  1
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                  0
`define CH1_DQ1_SWI_DQS_TX_QDR_M1_R1_CFG_8___POR                             32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                               'h00000D00
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1                               'h00000D04
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2                               'h00000D08
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3                               'h00000D0C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4                               'h00000D10
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5                               'h00000D14
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6                               'h00000D18
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7                               'h00000D1C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8                               'h00000D20
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                               'h00000D24
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1                               'h00000D28
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2                               'h00000D2C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3                               'h00000D30
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4                               'h00000D34
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5                               'h00000D38
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6                               'h00000D3C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7                               'h00000D40
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8                               'h00000D44
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                               'h00000D48
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1                               'h00000D4C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2                               'h00000D50
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3                               'h00000D54
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4                               'h00000D58
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5                               'h00000D5C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6                               'h00000D60
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7                               'h00000D64
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8                               'h00000D68
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                               'h00000D6C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1                               'h00000D70
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_1___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2                               'h00000D74
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_2___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3                               'h00000D78
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_3___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4                               'h00000D7C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_4___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5                               'h00000D80
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_5___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6                               'h00000D84
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_6___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7                               'h00000D88
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_7___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8                               'h00000D8C
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              4
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              0
`define CH1_DQ1_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_8___POR                       32'h00000000

`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                    'h00000D90
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1                                    'h00000D94
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R0_CFG_1___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                    'h00000D98
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1                                    'h00000D9C
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M0_R1_CFG_1___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                    'h00000DA0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1                                    'h00000DA4
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R0_CFG_1___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                    'h00000DA8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1                                    'h00000DAC
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__GEAR                                     7:6
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__EN                                         8
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                 5:0
`define CH1_DQ1_SWI_DQS_TX_LPDE_M1_R1_CFG_1___POR                            32'h00000100

`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0                                         'h00000DB0
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                       8:6
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                          5
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                      11:9
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                      4
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                      3
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                      2:0
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_0___POR                                 32'h00000041

`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1                                         'h00000DB4
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__TX_IMPD                                       8:6
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__SW_OVR                                          5
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__RX_IMPD                                      11:9
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_T                                      4
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_VAL_C                                      3
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1__OVRD_SEL                                      2:0
`define CH1_DQ1_SWI_DQS_TX_IO_M0_CFG_1___POR                                 32'h00000041

`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0                                         'h00000DB8
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                       8:6
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                          5
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                      11:9
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                      4
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                      3
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                      2:0
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_0___POR                                 32'h00000041

`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1                                         'h00000DBC
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__TX_IMPD                                       8:6
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__SW_OVR                                          5
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__RX_IMPD                                      11:9
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_T                                      4
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_VAL_C                                      3
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1__OVRD_SEL                                      2:0
`define CH1_DQ1_SWI_DQS_TX_IO_M1_CFG_1___POR                                 32'h00000041

`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                    'h00000DC0
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                   13
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                    10:5
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                     4:0
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                   12
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                     11
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                            32'h00000001

`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                    'h00000DC4
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                   13
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                    10:5
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                     4:0
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                   12
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                     11
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                            32'h00000001

`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                    'h00000DC8
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                   13
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                    10:5
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                     4:0
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                   12
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                     11
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                            32'h00000001

`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                    'h00000DCC
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                   13
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                    10:5
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                     4:0
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                   12
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                     11
`define CH1_DQ1_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                            32'h00000001

`define CH1_CA_SWI_TOP_CFG                                                     'h00000000
`define CH1_CA_SWI_TOP_CFG__WCS_SW_OVR_VAL                                              1
`define CH1_CA_SWI_TOP_CFG__WCS_SW_OVR                                                  0
`define CH1_CA_SWI_TOP_CFG__TRAINING_MODE                                               9
`define CH1_CA_SWI_TOP_CFG__RCS_SW_OVR_VAL                                              3
`define CH1_CA_SWI_TOP_CFG__RCS_SW_OVR                                                  2
`define CH1_CA_SWI_TOP_CFG__FIFO_CLR                                                    8
`define CH1_CA_SWI_TOP_CFG___POR                                             32'h00000000

`define CH1_CA_SWI_TOP_STA                                                     'h00000004
`define CH1_CA_SWI_TOP_STA__WCS                                                         0
`define CH1_CA_SWI_TOP_STA__RCS                                                         1
`define CH1_CA_SWI_TOP_STA___POR                                             32'h00000000

`define CH1_CA_SWI_DQ_RX_BSCAN_STA                                             'h00000008
`define CH1_CA_SWI_DQ_RX_BSCAN_STA__VAL                                              10:0
`define CH1_CA_SWI_DQ_RX_BSCAN_STA___POR                                     32'h00000000

`define CH1_CA_SWI_DQ_RX_M0_CFG                                                'h0000000C
`define CH1_CA_SWI_DQ_RX_M0_CFG__RGB_MODE                                             2:0
`define CH1_CA_SWI_DQ_RX_M0_CFG__FGB_MODE                                             7:4
`define CH1_CA_SWI_DQ_RX_M0_CFG___POR                                        32'h00000074

`define CH1_CA_SWI_DQ_RX_M1_CFG                                                'h00000010
`define CH1_CA_SWI_DQ_RX_M1_CFG__RGB_MODE                                             2:0
`define CH1_CA_SWI_DQ_RX_M1_CFG__FGB_MODE                                             7:4
`define CH1_CA_SWI_DQ_RX_M1_CFG___POR                                        32'h00000074

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_0                                        'h00000014
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_0__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_1                                        'h00000018
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_1__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_2                                        'h0000001C
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_2__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_3                                        'h00000020
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_3__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_4                                        'h00000024
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_4__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_5                                        'h00000028
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_5__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_6                                        'h0000002C
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_6__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_7                                        'h00000030
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_7__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_8                                        'h00000034
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_8__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_9                                        'h00000038
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_9__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_10                                       'h0000003C
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_10__RESERVED0                                   7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R0_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_0                                        'h00000040
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_0__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_1                                        'h00000044
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_1__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_2                                        'h00000048
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_2__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_3                                        'h0000004C
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_3__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_4                                        'h00000050
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_4__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_5                                        'h00000054
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_5__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_6                                        'h00000058
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_6__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_7                                        'h0000005C
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_7__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_8                                        'h00000060
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_8__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_9                                        'h00000064
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_9__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_10                                       'h00000068
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_10__RESERVED0                                   7:0
`define CH1_CA_SWI_DQ_RX_IO_M0_R1_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_0                                        'h0000006C
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_0__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_1                                        'h00000070
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_1__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_2                                        'h00000074
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_2__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_3                                        'h00000078
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_3__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_4                                        'h0000007C
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_4__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_5                                        'h00000080
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_5__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_6                                        'h00000084
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_6__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_7                                        'h00000088
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_7__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_8                                        'h0000008C
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_8__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_9                                        'h00000090
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_9__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_10                                       'h00000094
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_10__RESERVED0                                   7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R0_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_0                                        'h00000098
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_0__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_1                                        'h0000009C
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_1__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_2                                        'h000000A0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_2__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_3                                        'h000000A4
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_3__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_4                                        'h000000A8
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_4__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_5                                        'h000000AC
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_5__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_6                                        'h000000B0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_6__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_7                                        'h000000B4
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_7__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_8                                        'h000000B8
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_8__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_9                                        'h000000BC
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_9__RESERVED0                                    7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_10                                       'h000000C0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_10__RESERVED0                                   7:0
`define CH1_CA_SWI_DQ_RX_IO_M1_R1_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_IO_STA                                                'h000000C4
`define CH1_CA_SWI_DQ_RX_IO_STA__CORE_IG                                             31:0
`define CH1_CA_SWI_DQ_RX_IO_STA___POR                                        32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0                                        'h000000C8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1                                        'h000000CC
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2                                        'h000000D0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3                                        'h000000D4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4                                        'h000000D8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5                                        'h000000DC
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6                                        'h000000E0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7                                        'h000000E4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8                                        'h000000E8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9                                        'h000000EC
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10                                       'h000000F0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R0_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0                                        'h000000F4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1                                        'h000000F8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2                                        'h000000FC
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3                                        'h00000100
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4                                        'h00000104
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5                                        'h00000108
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6                                        'h0000010C
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7                                        'h00000110
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8                                        'h00000114
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9                                        'h00000118
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10                                       'h0000011C
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQ_RX_SA_M0_R1_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0                                        'h00000120
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1                                        'h00000124
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2                                        'h00000128
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3                                        'h0000012C
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4                                        'h00000130
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5                                        'h00000134
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6                                        'h00000138
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7                                        'h0000013C
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8                                        'h00000140
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9                                        'h00000144
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10                                       'h00000148
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R0_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0                                        'h0000014C
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_0___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1                                        'h00000150
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_1___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2                                        'h00000154
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_2___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3                                        'h00000158
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_3___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4                                        'h0000015C
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_4___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5                                        'h00000160
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_5___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6                                        'h00000164
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_6___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7                                        'h00000168
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_7___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8                                        'h0000016C
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_8___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9                                        'h00000170
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_90                                    17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_270                                   19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_180                                   18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_DIR_0                                     16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_90                                  7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_270                               15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_180                                11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9__CAL_CODE_0                                   3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_9___POR                                32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10                                       'h00000174
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQ_RX_SA_M1_R1_CFG_10___POR                               32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0                                    'h00000178
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_0___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1                                    'h0000017C
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_1___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2                                    'h00000180
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_2___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3                                    'h00000184
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_3___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4                                    'h00000188
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_4___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5                                    'h0000018C
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_5___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6                                    'h00000190
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_6___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7                                    'h00000194
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_7___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8                                    'h00000198
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_8___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9                                    'h0000019C
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_9___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10                                   'h000001A0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_90                                 9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_270                              25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_180                              17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__GEAR_0                                  1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_90                               15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_270                              31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_180                              23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10__CTRL_0                                  7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R0_CFG_10___POR                           32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0                                    'h000001A4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_0___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1                                    'h000001A8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_1___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2                                    'h000001AC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_2___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3                                    'h000001B0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_3___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4                                    'h000001B4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_4___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5                                    'h000001B8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_5___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6                                    'h000001BC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_6___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7                                    'h000001C0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_7___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8                                    'h000001C4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_8___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9                                    'h000001C8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_9___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10                                   'h000001CC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_90                                 9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_270                              25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_180                              17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__GEAR_0                                  1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_90                               15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_270                              31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_180                              23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10__CTRL_0                                  7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M0_R1_CFG_10___POR                           32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0                                    'h000001D0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_0___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1                                    'h000001D4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_1___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2                                    'h000001D8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_2___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3                                    'h000001DC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_3___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4                                    'h000001E0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_4___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5                                    'h000001E4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_5___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6                                    'h000001E8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_6___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7                                    'h000001EC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_7___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8                                    'h000001F0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_8___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9                                    'h000001F4
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_9___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10                                   'h000001F8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_90                                 9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_270                              25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_180                              17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__GEAR_0                                  1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_90                               15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_270                              31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_180                              23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10__CTRL_0                                  7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R0_CFG_10___POR                           32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0                                    'h000001FC
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_0___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1                                    'h00000200
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_1___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2                                    'h00000204
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_2___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3                                    'h00000208
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_3___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4                                    'h0000020C
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_4___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5                                    'h00000210
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_5___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6                                    'h00000214
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_6___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7                                    'h00000218
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_7___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8                                    'h0000021C
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_8___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9                                    'h00000220
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_90                                  9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_270                               25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_180                               17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__GEAR_0                                   1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_90                                15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_270                               31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_180                               23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9__CTRL_0                                   7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_9___POR                            32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10                                   'h00000224
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_90                                 9:8
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_270                              25:24
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_180                              17:16
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__GEAR_0                                  1:0
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_90                               15:10
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_270                              31:26
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_180                              23:18
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10__CTRL_0                                  7:2
`define CH1_CA_SWI_DQ_RX_SA_DLY_M1_R1_CFG_10___POR                           32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_0                                              'h00000228
`define CH1_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_0__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_0___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_1                                              'h0000022C
`define CH1_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_1__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_1___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_2                                              'h00000230
`define CH1_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_2__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_2___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_3                                              'h00000234
`define CH1_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_3__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_3___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_4                                              'h00000238
`define CH1_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_4__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_4___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_5                                              'h0000023C
`define CH1_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_5__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_5___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_6                                              'h00000240
`define CH1_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_6__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_6___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_7                                              'h00000244
`define CH1_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_7__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_7___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_8                                              'h00000248
`define CH1_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_8__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_8___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_9                                              'h0000024C
`define CH1_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_90                                            1
`define CH1_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_270                                           3
`define CH1_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_180                                           2
`define CH1_CA_SWI_DQ_RX_SA_STA_9__SA_OUT_0                                             0
`define CH1_CA_SWI_DQ_RX_SA_STA_9___POR                                      32'h00000000

`define CH1_CA_SWI_DQ_RX_SA_STA_10                                             'h00000250
`define CH1_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_90                                           1
`define CH1_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_270                                          3
`define CH1_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_180                                          2
`define CH1_CA_SWI_DQ_RX_SA_STA_10__SA_OUT_0                                            0
`define CH1_CA_SWI_DQ_RX_SA_STA_10___POR                                     32'h00000000

`define CH1_CA_SWI_DQ_TX_BSCAN_CFG                                             'h00000254
`define CH1_CA_SWI_DQ_TX_BSCAN_CFG__VAL                                              10:0
`define CH1_CA_SWI_DQ_TX_BSCAN_CFG___POR                                     32'h00000000

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0                                   'h00000258
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_0___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1                                   'h0000025C
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_1___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2                                   'h00000260
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_2___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3                                   'h00000264
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_3___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4                                   'h00000268
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_4___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5                                   'h0000026C
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_5___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6                                   'h00000270
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_6___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7                                   'h00000274
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_7___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8                                   'h00000278
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_8___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9                                   'h0000027C
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_9___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10                                  'h00000280
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10__EGRESS_MODE                            5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M0_CFG_10___POR                          32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0                                   'h00000284
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_0___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1                                   'h00000288
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_1___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2                                   'h0000028C
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_2___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3                                   'h00000290
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_3___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4                                   'h00000294
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_4___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5                                   'h00000298
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_5___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6                                   'h0000029C
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_6___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7                                   'h000002A0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_7___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8                                   'h000002A4
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_8___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9                                   'h000002A8
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9__EGRESS_MODE                             5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_9___POR                           32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10                                  'h000002AC
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10__EGRESS_MODE                            5:0
`define CH1_CA_SWI_DQ_TX_EGRESS_ANA_M1_CFG_10___POR                          32'h00000001

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0                                   'h000002B0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_0___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1                                   'h000002B4
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_1___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2                                   'h000002B8
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_2___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3                                   'h000002BC
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_3___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4                                   'h000002C0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_4___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5                                   'h000002C4
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_5___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6                                   'h000002C8
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_6___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7                                   'h000002CC
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_7___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8                                   'h000002D0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_8___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9                                   'h000002D4
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_9___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10                                  'h000002D8
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10__EGRESS_MODE                            6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M0_CFG_10___POR                          32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0                                   'h000002DC
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_0___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1                                   'h000002E0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_1___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2                                   'h000002E4
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_2___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3                                   'h000002E8
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_3___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4                                   'h000002EC
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_4___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5                                   'h000002F0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_5___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6                                   'h000002F4
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_6___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7                                   'h000002F8
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_7___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8                                   'h000002FC
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_8___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9                                   'h00000300
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9__EGRESS_MODE                             6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_9___POR                           32'h00000002

`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10                                  'h00000304
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10__EGRESS_MODE                            6:0
`define CH1_CA_SWI_DQ_TX_EGRESS_DIG_M1_CFG_10___POR                          32'h00000002

`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG                                      'h00000308
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__EN                                          14
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R0_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG                                      'h0000030C
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__EN                                          14
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQ_TX_ODR_PI_M0_R1_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG                                      'h00000310
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__EN                                          14
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R0_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG                                      'h00000314
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__EN                                          14
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQ_TX_ODR_PI_M1_R1_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG                                    'h00000318
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG                                    'h0000031C
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M0_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG                                    'h00000320
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG                                    'h00000324
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_0_M1_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG                                    'h00000328
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG                                    'h0000032C
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M0_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG                                    'h00000330
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG                                    'h00000334
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_QDR_PI_1_M1_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG                                    'h00000338
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG                                    'h0000033C
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M0_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG                                    'h00000340
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG                                    'h00000344
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_0_M1_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG                                    'h00000348
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG                                    'h0000034C
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M0_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG                                    'h00000350
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R0_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG                                    'h00000354
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__XCPL                                   13:10
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__GEAR                                     9:6
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__EN                                        14
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG__CODE                                     5:0
`define CH1_CA_SWI_DQ_TX_DDR_PI_1_M1_R1_CFG___POR                            32'h00000040

`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG                                       'h00000358
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__XCPL                                      13:10
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__GEAR                                        9:6
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__EN                                           14
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG__CODE                                        5:0
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R0_CFG___POR                               32'h00000040

`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG                                       'h0000035C
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__XCPL                                      13:10
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__GEAR                                        9:6
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__EN                                           14
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG__CODE                                        5:0
`define CH1_CA_SWI_DQ_TX_PI_RT_M0_R1_CFG___POR                               32'h00000040

`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG                                       'h00000360
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__XCPL                                      13:10
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__GEAR                                        9:6
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__EN                                           14
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG__CODE                                        5:0
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R0_CFG___POR                               32'h00000040

`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG                                       'h00000364
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__XCPL                                      13:10
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__GEAR                                        9:6
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__EN                                           14
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG__CODE                                        5:0
`define CH1_CA_SWI_DQ_TX_PI_RT_M1_R1_CFG___POR                               32'h00000040

`define CH1_CA_SWI_DQ_TX_RT_M0_R0_CFG                                          'h00000368
`define CH1_CA_SWI_DQ_TX_RT_M0_R0_CFG__PIPE_EN                                       10:0
`define CH1_CA_SWI_DQ_TX_RT_M0_R0_CFG___POR                                  32'h00000000

`define CH1_CA_SWI_DQ_TX_RT_M0_R1_CFG                                          'h0000036C
`define CH1_CA_SWI_DQ_TX_RT_M0_R1_CFG__PIPE_EN                                       10:0
`define CH1_CA_SWI_DQ_TX_RT_M0_R1_CFG___POR                                  32'h00000000

`define CH1_CA_SWI_DQ_TX_RT_M1_R0_CFG                                          'h00000370
`define CH1_CA_SWI_DQ_TX_RT_M1_R0_CFG__PIPE_EN                                       10:0
`define CH1_CA_SWI_DQ_TX_RT_M1_R0_CFG___POR                                  32'h00000000

`define CH1_CA_SWI_DQ_TX_RT_M1_R1_CFG                                          'h00000374
`define CH1_CA_SWI_DQ_TX_RT_M1_R1_CFG__PIPE_EN                                       10:0
`define CH1_CA_SWI_DQ_TX_RT_M1_R1_CFG___POR                                  32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0                                       'h00000378
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1                                       'h0000037C
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2                                       'h00000380
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3                                       'h00000384
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4                                       'h00000388
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5                                       'h0000038C
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6                                       'h00000390
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7                                       'h00000394
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8                                       'h00000398
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9                                       'h0000039C
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10                                      'h000003A0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0                                       'h000003A4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1                                       'h000003A8
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2                                       'h000003AC
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3                                       'h000003B0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4                                       'h000003B4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5                                       'h000003B8
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6                                       'h000003BC
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7                                       'h000003C0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8                                       'h000003C4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9                                       'h000003C8
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10                                      'h000003CC
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_SDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0                                       'h000003D0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1                                       'h000003D4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2                                       'h000003D8
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3                                       'h000003DC
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4                                       'h000003E0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5                                       'h000003E4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6                                       'h000003E8
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7                                       'h000003EC
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8                                       'h000003F0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9                                       'h000003F4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10                                      'h000003F8
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0                                       'h000003FC
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1                                       'h00000400
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2                                       'h00000404
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3                                       'h00000408
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4                                       'h0000040C
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5                                       'h00000410
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6                                       'h00000414
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7                                       'h00000418
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8                                       'h0000041C
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9                                       'h00000420
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P7                                    7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P6                                    6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P5                                    5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P4                                    4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10                                      'h00000424
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_SDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0                                 'h00000428
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1                                 'h0000042C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2                                 'h00000430
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3                                 'h00000434
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4                                 'h00000438
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5                                 'h0000043C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6                                 'h00000440
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7                                 'h00000444
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8                                 'h00000448
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9                                 'h0000044C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10                                'h00000450
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0                                 'h00000454
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1                                 'h00000458
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2                                 'h0000045C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3                                 'h00000460
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4                                 'h00000464
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5                                 'h00000468
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6                                 'h0000046C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7                                 'h00000470
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8                                 'h00000474
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9                                 'h00000478
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10                                'h0000047C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0                                 'h00000480
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1                                 'h00000484
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2                                 'h00000488
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3                                 'h0000048C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4                                 'h00000490
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5                                 'h00000494
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6                                 'h00000498
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7                                 'h0000049C
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8                                 'h000004A0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9                                 'h000004A4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10                                'h000004A8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0                                 'h000004AC
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1                                 'h000004B0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2                                 'h000004B4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3                                 'h000004B8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4                                 'h000004BC
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5                                 'h000004C0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6                                 'h000004C4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7                                 'h000004C8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8                                 'h000004CC
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9                                 'h000004D0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P7                            30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P6                            26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P5                            22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P4                            18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P3                            14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P2                             10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                              6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                              2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10                                'h000004D4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQ_TX_SDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0                                'h000004D8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1                                'h000004DC
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_1___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2                                'h000004E0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_2___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3                                'h000004E4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_3___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4                                'h000004E8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_4___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5                                'h000004EC
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_5___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6                                'h000004F0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_6___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7                                'h000004F4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_7___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8                                'h000004F8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_8___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9                                'h000004FC
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_9___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10                               'h00000500
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P7                            29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P6                            25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P5                            21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P4                            17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P3                            13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P2                              9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P1                              5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10__DLY_P0                              1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R0_CFG_10___POR                       32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0                                'h00000504
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1                                'h00000508
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_1___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2                                'h0000050C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_2___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3                                'h00000510
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_3___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4                                'h00000514
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_4___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5                                'h00000518
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_5___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6                                'h0000051C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_6___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7                                'h00000520
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_7___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8                                'h00000524
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_8___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9                                'h00000528
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_9___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10                               'h0000052C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P7                            29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P6                            25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P5                            21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P4                            17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P3                            13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P2                              9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P1                              5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10__DLY_P0                              1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M0_R1_CFG_10___POR                       32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0                                'h00000530
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1                                'h00000534
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_1___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2                                'h00000538
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_2___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3                                'h0000053C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_3___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4                                'h00000540
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_4___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5                                'h00000544
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_5___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6                                'h00000548
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_6___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7                                'h0000054C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_7___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8                                'h00000550
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_8___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9                                'h00000554
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_9___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10                               'h00000558
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P7                            29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P6                            25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P5                            21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P4                            17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P3                            13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P2                              9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P1                              5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10__DLY_P0                              1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R0_CFG_10___POR                       32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0                                'h0000055C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1                                'h00000560
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_1___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2                                'h00000564
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_2___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3                                'h00000568
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_3___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4                                'h0000056C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_4___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5                                'h00000570
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_5___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6                                'h00000574
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_6___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7                                'h00000578
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_7___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8                                'h0000057C
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_8___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9                                'h00000580
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P7                             29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P6                             25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P5                             21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P4                             17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P3                             13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P2                               9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P1                               5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9__DLY_P0                               1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_9___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10                               'h00000584
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P7                            29:28
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P6                            25:24
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P5                            21:20
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P4                            17:16
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P3                            13:12
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P2                              9:8
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P1                              5:4
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10__DLY_P0                              1:0
`define CH1_CA_SWI_DQ_TX_SDR_FC_DLY_M1_R1_CFG_10___POR                       32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0                                       'h00000588
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1                                       'h0000058C
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2                                       'h00000590
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3                                       'h00000594
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4                                       'h00000598
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5                                       'h0000059C
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6                                       'h000005A0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7                                       'h000005A4
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8                                       'h000005A8
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9                                       'h000005AC
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10                                      'h000005B0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0                                       'h000005B4
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1                                       'h000005B8
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2                                       'h000005BC
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3                                       'h000005C0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4                                       'h000005C4
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5                                       'h000005C8
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6                                       'h000005CC
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7                                       'h000005D0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8                                       'h000005D4
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9                                       'h000005D8
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10                                      'h000005DC
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_DDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0                                       'h000005E0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1                                       'h000005E4
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2                                       'h000005E8
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3                                       'h000005EC
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4                                       'h000005F0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5                                       'h000005F4
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6                                       'h000005F8
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7                                       'h000005FC
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8                                       'h00000600
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9                                       'h00000604
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10                                      'h00000608
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0                                       'h0000060C
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1                                       'h00000610
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2                                       'h00000614
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3                                       'h00000618
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4                                       'h0000061C
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5                                       'h00000620
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6                                       'h00000624
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7                                       'h00000628
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8                                       'h0000062C
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9                                       'h00000630
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P3                                    3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P2                                    2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10                                      'h00000634
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_DDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0                                 'h00000638
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1                                 'h0000063C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2                                 'h00000640
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3                                 'h00000644
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4                                 'h00000648
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5                                 'h0000064C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6                                 'h00000650
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7                                 'h00000654
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8                                 'h00000658
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9                                 'h0000065C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10                                'h00000660
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0                                 'h00000664
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1                                 'h00000668
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2                                 'h0000066C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3                                 'h00000670
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4                                 'h00000674
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5                                 'h00000678
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6                                 'h0000067C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7                                 'h00000680
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8                                 'h00000684
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9                                 'h00000688
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10                                'h0000068C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0                                 'h00000690
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1                                 'h00000694
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2                                 'h00000698
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3                                 'h0000069C
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4                                 'h000006A0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5                                 'h000006A4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6                                 'h000006A8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7                                 'h000006AC
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8                                 'h000006B0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9                                 'h000006B4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10                                'h000006B8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0                                 'h000006BC
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1                                 'h000006C0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2                                 'h000006C4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3                                 'h000006C8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4                                 'h000006CC
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5                                 'h000006D0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6                                 'h000006D4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7                                 'h000006D8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8                                 'h000006DC
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9                                 'h000006E0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P3                            13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P2                              9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                              5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                              1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10                                'h000006E4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQ_TX_DDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0                                       'h000006E8
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1                                       'h000006EC
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2                                       'h000006F0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3                                       'h000006F4
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4                                       'h000006F8
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5                                       'h000006FC
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6                                       'h00000700
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7                                       'h00000704
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8                                       'h00000708
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9                                       'h0000070C
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10                                      'h00000710
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0                                       'h00000714
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1                                       'h00000718
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2                                       'h0000071C
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3                                       'h00000720
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4                                       'h00000724
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5                                       'h00000728
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6                                       'h0000072C
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7                                       'h00000730
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8                                       'h00000734
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9                                       'h00000738
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10                                      'h0000073C
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_QDR_M0_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0                                       'h00000740
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1                                       'h00000744
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2                                       'h00000748
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3                                       'h0000074C
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4                                       'h00000750
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5                                       'h00000754
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6                                       'h00000758
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7                                       'h0000075C
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8                                       'h00000760
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9                                       'h00000764
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10                                      'h00000768
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R0_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0                                       'h0000076C
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1                                       'h00000770
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_1___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2                                       'h00000774
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_2___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3                                       'h00000778
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_3___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4                                       'h0000077C
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_4___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5                                       'h00000780
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_5___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6                                       'h00000784
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_6___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7                                       'h00000788
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_7___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8                                       'h0000078C
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_8___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9                                       'h00000790
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9__PIPE_EN_P1                                    1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9__PIPE_EN_P0                                    0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_9___POR                               32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10                                      'h00000794
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQ_TX_QDR_M1_R1_CFG_10___POR                              32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0                                 'h00000798
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1                                 'h0000079C
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2                                 'h000007A0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3                                 'h000007A4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4                                 'h000007A8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5                                 'h000007AC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6                                 'h000007B0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7                                 'h000007B4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8                                 'h000007B8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9                                 'h000007BC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10                                'h000007C0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10__X_SEL_P1                               4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10__X_SEL_P0                               0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0                                 'h000007C4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1                                 'h000007C8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2                                 'h000007CC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3                                 'h000007D0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4                                 'h000007D4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5                                 'h000007D8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6                                 'h000007DC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7                                 'h000007E0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8                                 'h000007E4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9                                 'h000007E8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10                                'h000007EC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10__X_SEL_P1                               4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10__X_SEL_P0                               0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M0_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0                                 'h000007F0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1                                 'h000007F4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2                                 'h000007F8
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3                                 'h000007FC
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4                                 'h00000800
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5                                 'h00000804
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6                                 'h00000808
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7                                 'h0000080C
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8                                 'h00000810
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9                                 'h00000814
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10                                'h00000818
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10__X_SEL_P1                               4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10__X_SEL_P0                               0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R0_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0                                 'h0000081C
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_0___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1                                 'h00000820
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_1___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2                                 'h00000824
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_2___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3                                 'h00000828
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_3___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4                                 'h0000082C
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_4___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5                                 'h00000830
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_5___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6                                 'h00000834
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_6___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7                                 'h00000838
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_7___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8                                 'h0000083C
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_8___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9                                 'h00000840
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9__X_SEL_P1                                4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9__X_SEL_P0                                0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_9___POR                         32'h00000000

`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10                                'h00000844
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10__X_SEL_P1                               4
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10__X_SEL_P0                               0
`define CH1_CA_SWI_DQ_TX_QDR_X_SEL_M1_R1_CFG_10___POR                        32'h00000000

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0                                      'h00000848
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_0___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1                                      'h0000084C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_1___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2                                      'h00000850
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_2___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3                                      'h00000854
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_3___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4                                      'h00000858
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_4___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5                                      'h0000085C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_5___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6                                      'h00000860
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_6___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7                                      'h00000864
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_7___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8                                      'h00000868
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_8___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9                                      'h0000086C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_9___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10                                     'h00000870
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__GEAR                                      7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__EN                                          8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R0_CFG_10___POR                             32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0                                      'h00000874
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_0___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1                                      'h00000878
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_1___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2                                      'h0000087C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_2___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3                                      'h00000880
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_3___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4                                      'h00000884
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_4___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5                                      'h00000888
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_5___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6                                      'h0000088C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_6___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7                                      'h00000890
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_7___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8                                      'h00000894
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_8___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9                                      'h00000898
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_9___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10                                     'h0000089C
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__GEAR                                      7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__EN                                          8
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M0_R1_CFG_10___POR                             32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0                                      'h000008A0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_0___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1                                      'h000008A4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_1___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2                                      'h000008A8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_2___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3                                      'h000008AC
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_3___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4                                      'h000008B0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_4___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5                                      'h000008B4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_5___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6                                      'h000008B8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_6___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7                                      'h000008BC
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_7___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8                                      'h000008C0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_8___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9                                      'h000008C4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_9___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10                                     'h000008C8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__GEAR                                      7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__EN                                          8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R0_CFG_10___POR                             32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0                                      'h000008CC
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_0___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1                                      'h000008D0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_1___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2                                      'h000008D4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_2___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3                                      'h000008D8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_3___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4                                      'h000008DC
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_4___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5                                      'h000008E0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_5___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6                                      'h000008E4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_6___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7                                      'h000008E8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_7___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8                                      'h000008EC
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_8___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9                                      'h000008F0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__GEAR                                       7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__EN                                           8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9__CTRL_BIN                                   5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_9___POR                              32'h00000100

`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10                                     'h000008F4
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__GEAR                                      7:6
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__EN                                          8
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQ_TX_LPDE_M1_R1_CFG_10___POR                             32'h00000100

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0                                           'h000008F8
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_0___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1                                           'h000008FC
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_1___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2                                           'h00000900
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_2___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3                                           'h00000904
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_3___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4                                           'h00000908
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_4___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5                                           'h0000090C
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_5___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6                                           'h00000910
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_6___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7                                           'h00000914
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_7___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8                                           'h00000918
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_8___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9                                           'h0000091C
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_9___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10                                          'h00000920
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__TX_IMPD                                        8:6
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__SW_OVR                                           5
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__RX_IMPD                                       11:9
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__RESERVED0                                        4
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__OVRD_VAL                                         3
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10__OVRD_SEL                                       2:0
`define CH1_CA_SWI_DQ_TX_IO_M0_CFG_10___POR                                  32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0                                           'h00000924
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_0___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1                                           'h00000928
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_1___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2                                           'h0000092C
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_2___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3                                           'h00000930
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_3___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4                                           'h00000934
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_4___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5                                           'h00000938
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_5___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6                                           'h0000093C
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_6___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7                                           'h00000940
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_7___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8                                           'h00000944
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_8___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9                                           'h00000948
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__TX_IMPD                                         8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__SW_OVR                                            5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__RX_IMPD                                        11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__RESERVED0                                         4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__OVRD_VAL                                          3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9__OVRD_SEL                                        2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_9___POR                                   32'h00000040

`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10                                          'h0000094C
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__TX_IMPD                                        8:6
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__SW_OVR                                           5
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__RX_IMPD                                       11:9
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__RESERVED0                                        4
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__OVRD_VAL                                         3
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10__OVRD_SEL                                       2:0
`define CH1_CA_SWI_DQ_TX_IO_M1_CFG_10___POR                                  32'h00000040

`define CH1_CA_SWI_DQS_RX_M0_CFG                                               'h00000950
`define CH1_CA_SWI_DQS_RX_M0_CFG__WCK_MODE                                              8
`define CH1_CA_SWI_DQS_RX_M0_CFG__RGB_MODE                                            2:0
`define CH1_CA_SWI_DQS_RX_M0_CFG__PRE_FILTER_SEL                                    13:12
`define CH1_CA_SWI_DQS_RX_M0_CFG__FGB_MODE                                            7:4
`define CH1_CA_SWI_DQS_RX_M0_CFG___POR                                       32'h00000074

`define CH1_CA_SWI_DQS_RX_M1_CFG                                               'h00000954
`define CH1_CA_SWI_DQS_RX_M1_CFG__WCK_MODE                                              8
`define CH1_CA_SWI_DQS_RX_M1_CFG__RGB_MODE                                            2:0
`define CH1_CA_SWI_DQS_RX_M1_CFG__PRE_FILTER_SEL                                    13:12
`define CH1_CA_SWI_DQS_RX_M1_CFG__FGB_MODE                                            7:4
`define CH1_CA_SWI_DQS_RX_M1_CFG___POR                                       32'h00000074

`define CH1_CA_SWI_DQS_RX_BSCAN_STA                                            'h00000958
`define CH1_CA_SWI_DQS_RX_BSCAN_STA__VAL                                              1:0
`define CH1_CA_SWI_DQS_RX_BSCAN_STA___POR                                    32'h00000000

`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG                                   'h0000095C
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__GEAR                                    7:6
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__EN                                        8
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG__CTRL_BIN                                5:0
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R0_CFG___POR                           32'h00000100

`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG                                   'h00000960
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__GEAR                                    7:6
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__EN                                        8
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG__CTRL_BIN                                5:0
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M0_R1_CFG___POR                           32'h00000100

`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG                                   'h00000964
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__GEAR                                    7:6
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__EN                                        8
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG__CTRL_BIN                                5:0
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R0_CFG___POR                           32'h00000100

`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG                                   'h00000968
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__GEAR                                    7:6
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__EN                                        8
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG__CTRL_BIN                                5:0
`define CH1_CA_SWI_DQS_RX_SDR_LPDE_M1_R1_CFG___POR                           32'h00000100

`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG                                     'h0000096C
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG                                     'h00000970
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_REN_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG                                     'h00000974
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG                                     'h00000978
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_REN_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG                                     'h0000097C
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG                                     'h00000980
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_RCS_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG                                     'h00000984
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG                                     'h00000988
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_RX_RCS_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG                                  'h0000098C
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R0_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG                                  'h00000990
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M0_R1_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG                                  'h00000994
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R0_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG                                  'h00000998
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_0_M1_R1_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG                                  'h0000099C
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R0_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG                                  'h000009A0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M0_R1_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG                                  'h000009A4
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R0_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG                                  'h000009A8
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__XCPL                                 13:10
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__GEAR                                   9:6
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__EN                                      14
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG__CODE                                   5:0
`define CH1_CA_SWI_DQS_RX_RDQS_PI_1_M1_R1_CFG___POR                          32'h00000040

`define CH1_CA_SWI_DQS_RX_PI_STA                                               'h000009AC
`define CH1_CA_SWI_DQS_RX_PI_STA__REN_PI_PHASE                                          0
`define CH1_CA_SWI_DQS_RX_PI_STA__RCS_PI_PHASE                                          1
`define CH1_CA_SWI_DQS_RX_PI_STA___POR                                       32'h00000000

`define CH1_CA_SWI_DQS_RX_IO_M0_R0_CFG_0                                       'h000009B0
`define CH1_CA_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_T                                 15:8
`define CH1_CA_SWI_DQS_RX_IO_M0_R0_CFG_0__DLY_CTRL_C                                  7:0
`define CH1_CA_SWI_DQS_RX_IO_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_IO_M0_R1_CFG_0                                       'h000009B4
`define CH1_CA_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_T                                 15:8
`define CH1_CA_SWI_DQS_RX_IO_M0_R1_CFG_0__DLY_CTRL_C                                  7:0
`define CH1_CA_SWI_DQS_RX_IO_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_IO_M1_R0_CFG_0                                       'h000009B8
`define CH1_CA_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_T                                 15:8
`define CH1_CA_SWI_DQS_RX_IO_M1_R0_CFG_0__DLY_CTRL_C                                  7:0
`define CH1_CA_SWI_DQS_RX_IO_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_IO_M1_R1_CFG_0                                       'h000009BC
`define CH1_CA_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_T                                 15:8
`define CH1_CA_SWI_DQS_RX_IO_M1_R1_CFG_0__DLY_CTRL_C                                  7:0
`define CH1_CA_SWI_DQS_RX_IO_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG                                     'h000009C0
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SW_OVR                                     23
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__SE_MODE                                    22
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__RXCAL_EN                                   21
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__FB_EN                                   18:16
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__EN                                         20
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__DCPATH_EN                                  19
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_T                                   7:4
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_P_C                                   3:0
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_T                                 15:12
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG__CAL_N_C                                  11:8
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R0_CFG___POR                             32'h004A7777

`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG                                     'h000009C4
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SW_OVR                                     23
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__SE_MODE                                    22
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__RXCAL_EN                                   21
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__FB_EN                                   18:16
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__EN                                         20
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__DCPATH_EN                                  19
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_T                                   7:4
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_P_C                                   3:0
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_T                                 15:12
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG__CAL_N_C                                  11:8
`define CH1_CA_SWI_DQS_RX_IO_CMN_M0_R1_CFG___POR                             32'h004A7777

`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG                                     'h000009C8
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SW_OVR                                     23
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__SE_MODE                                    22
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__RXCAL_EN                                   21
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__FB_EN                                   18:16
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__EN                                         20
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__DCPATH_EN                                  19
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_T                                   7:4
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_P_C                                   3:0
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_T                                 15:12
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG__CAL_N_C                                  11:8
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R0_CFG___POR                             32'h004A7777

`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG                                     'h000009CC
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SW_OVR                                     23
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__SE_MODE                                    22
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__RXCAL_EN                                   21
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__FB_EN                                   18:16
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__EN                                         20
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__DCPATH_EN                                  19
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_T                                   7:4
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_P_C                                   3:0
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_T                                 15:12
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG__CAL_N_C                                  11:8
`define CH1_CA_SWI_DQS_RX_IO_CMN_M1_R1_CFG___POR                             32'h004A7777

`define CH1_CA_SWI_DQS_RX_IO_STA                                               'h000009D0
`define CH1_CA_SWI_DQS_RX_IO_STA__CORE_IG                                            31:0
`define CH1_CA_SWI_DQS_RX_IO_STA___POR                                       32'h00000000

`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0                                       'h000009D4
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQS_RX_SA_M0_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0                                       'h000009D8
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQS_RX_SA_M0_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0                                       'h000009DC
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQS_RX_SA_M1_R0_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0                                       'h000009E0
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_90                                   17
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_270                                  19
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_180                                  18
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_DIR_0                                    16
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_90                                 7:4
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_270                              15:12
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_180                               11:8
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0__CAL_CODE_0                                  3:0
`define CH1_CA_SWI_DQS_RX_SA_M1_R1_CFG_0___POR                               32'h00000000

`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG                                           'h000009E4
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG__SW_OVR                                            4
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_90_270                                     2
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG__OVR_EN_0_180                                      0
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_90_270                                     3
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG__CAL_EN_0_180                                      1
`define CH1_CA_SWI_DQS_RX_SA_CMN_CFG___POR                                   32'h00000005

`define CH1_CA_SWI_DQS_TX_M0_CFG                                               'h000009E8
`define CH1_CA_SWI_DQS_TX_M0_CFG__WGB_MODE                                            7:4
`define CH1_CA_SWI_DQS_TX_M0_CFG__TGB_MODE                                            2:0
`define CH1_CA_SWI_DQS_TX_M0_CFG__CK2WCK_RATIO                                        9:8
`define CH1_CA_SWI_DQS_TX_M0_CFG___POR                                       32'h00000087

`define CH1_CA_SWI_DQS_TX_M1_CFG                                               'h000009EC
`define CH1_CA_SWI_DQS_TX_M1_CFG__WGB_MODE                                            7:4
`define CH1_CA_SWI_DQS_TX_M1_CFG__TGB_MODE                                            2:0
`define CH1_CA_SWI_DQS_TX_M1_CFG__CK2WCK_RATIO                                        9:8
`define CH1_CA_SWI_DQS_TX_M1_CFG___POR                                       32'h00000087

`define CH1_CA_SWI_DQS_TX_BSCAN_CTRL_CFG                                       'h000009F0
`define CH1_CA_SWI_DQS_TX_BSCAN_CTRL_CFG__OE                                            1
`define CH1_CA_SWI_DQS_TX_BSCAN_CTRL_CFG__IE                                            0
`define CH1_CA_SWI_DQS_TX_BSCAN_CTRL_CFG___POR                               32'h00000000

`define CH1_CA_SWI_DQS_TX_BSCAN_CFG                                            'h000009F4
`define CH1_CA_SWI_DQS_TX_BSCAN_CFG__VAL                                              1:0
`define CH1_CA_SWI_DQS_TX_BSCAN_CFG___POR                                    32'h00000000

`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0                                  'h000009F8
`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0__EGRESS_MODE                            5:0
`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M0_CFG_0___POR                          32'h00000001

`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0                                  'h000009FC
`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0__EGRESS_MODE                            5:0
`define CH1_CA_SWI_DQS_TX_EGRESS_ANA_M1_CFG_0___POR                          32'h00000001

`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0                                  'h00000A00
`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0__EGRESS_MODE                            6:0
`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M0_CFG_0___POR                          32'h00000002

`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0                                  'h00000A04
`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0__EGRESS_MODE                            6:0
`define CH1_CA_SWI_DQS_TX_EGRESS_DIG_M1_CFG_0___POR                          32'h00000002

`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG                                     'h00000A08
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG                                     'h00000A0C
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_TX_ODR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG                                     'h00000A10
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG                                     'h00000A14
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG__CODE                                      5:0
`define CH1_CA_SWI_DQS_TX_ODR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG                                   'h00000A18
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG                                   'h00000A1C
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG                                   'h00000A20
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG                                   'h00000A24
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG                                   'h00000A28
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG                                   'h00000A2C
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG                                   'h00000A30
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG                                   'h00000A34
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_QDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG                                   'h00000A38
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG                                   'h00000A3C
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M0_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG                                   'h00000A40
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG                                   'h00000A44
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_0_M1_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG                                   'h00000A48
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG                                   'h00000A4C
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M0_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG                                   'h00000A50
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R0_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG                                   'h00000A54
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__XCPL                                  13:10
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__GEAR                                    9:6
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__EN                                       14
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG__CODE                                    5:0
`define CH1_CA_SWI_DQS_TX_DDR_PI_1_M1_R1_CFG___POR                           32'h00000040

`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG                                      'h00000A58
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__EN                                          14
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R0_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG                                      'h00000A5C
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__EN                                          14
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQS_TX_PI_RT_M0_R1_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG                                      'h00000A60
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__EN                                          14
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R0_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG                                      'h00000A64
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__XCPL                                     13:10
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__GEAR                                       9:6
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__EN                                          14
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG__CODE                                       5:0
`define CH1_CA_SWI_DQS_TX_PI_RT_M1_R1_CFG___POR                              32'h00000040

`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG                                     'h00000A68
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG                                     'h00000A6C
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_SDR_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG                                     'h00000A70
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG                                     'h00000A74
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_SDR_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG                                     'h00000A78
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG                                     'h00000A7C
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_DFI_PI_M0_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG                                     'h00000A80
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R0_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG                                     'h00000A84
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__XCPL                                    13:10
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__RSVD                                      5:0
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__GEAR                                      9:6
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG__EN                                         14
`define CH1_CA_SWI_DQS_TX_DFI_PI_M1_R1_CFG___POR                             32'h00000040

`define CH1_CA_SWI_DQS_TX_RT_M0_R0_CFG                                         'h00000A88
`define CH1_CA_SWI_DQS_TX_RT_M0_R0_CFG__PIPE_EN                                         0
`define CH1_CA_SWI_DQS_TX_RT_M0_R0_CFG___POR                                 32'h00000000

`define CH1_CA_SWI_DQS_TX_RT_M0_R1_CFG                                         'h00000A8C
`define CH1_CA_SWI_DQS_TX_RT_M0_R1_CFG__PIPE_EN                                         0
`define CH1_CA_SWI_DQS_TX_RT_M0_R1_CFG___POR                                 32'h00000000

`define CH1_CA_SWI_DQS_TX_RT_M1_R0_CFG                                         'h00000A90
`define CH1_CA_SWI_DQS_TX_RT_M1_R0_CFG__PIPE_EN                                         0
`define CH1_CA_SWI_DQS_TX_RT_M1_R0_CFG___POR                                 32'h00000000

`define CH1_CA_SWI_DQS_TX_RT_M1_R1_CFG                                         'h00000A94
`define CH1_CA_SWI_DQS_TX_RT_M1_R1_CFG__PIPE_EN                                         0
`define CH1_CA_SWI_DQS_TX_RT_M1_R1_CFG___POR                                 32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0                                      'h00000A98
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_SDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0                                      'h00000A9C
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_SDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0                                      'h00000AA0
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_SDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0                                      'h00000AA4
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P7                                   7
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P6                                   6
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P5                                   5
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P4                                   4
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_SDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0                                'h00000AA8
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0                                'h00000AAC
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0                                'h00000AB0
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0                                'h00000AB4
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P7                           30:28
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P6                           26:24
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P5                           22:20
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P4                           18:16
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           14:12
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                            10:8
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             6:4
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             2:0
`define CH1_CA_SWI_DQS_TX_SDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0                               'h00000AB8
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P7                            29:28
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P6                            25:24
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P5                            21:20
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P4                            17:16
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P3                            13:12
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P2                              9:8
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P1                              5:4
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0__DLY_P0                              1:0
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R0_CFG_0___POR                       32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0                               'h00000ABC
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P7                            29:28
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P6                            25:24
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P5                            21:20
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P4                            17:16
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P3                            13:12
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P2                              9:8
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P1                              5:4
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0__DLY_P0                              1:0
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M0_R1_CFG_0___POR                       32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0                               'h00000AC0
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P7                            29:28
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P6                            25:24
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P5                            21:20
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P4                            17:16
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P3                            13:12
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P2                              9:8
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P1                              5:4
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0__DLY_P0                              1:0
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R0_CFG_0___POR                       32'h00000000

`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0                               'h00000AC4
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P7                            29:28
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P6                            25:24
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P5                            21:20
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P4                            17:16
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P3                            13:12
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P2                              9:8
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P1                              5:4
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0__DLY_P0                              1:0
`define CH1_CA_SWI_DQS_TX_SDR_FC_DLY_M1_R1_CFG_0___POR                       32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0                                      'h00000AC8
`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_DDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0                                      'h00000ACC
`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_DDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0                                      'h00000AD0
`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_DDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0                                      'h00000AD4
`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P3                                   3
`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P2                                   2
`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_DDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0                                'h00000AD8
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0                                'h00000ADC
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0                                'h00000AE0
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0                                'h00000AE4
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P3                           13:12
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P2                             9:8
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                             5:4
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                             1:0
`define CH1_CA_SWI_DQS_TX_DDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0                                      'h00000AE8
`define CH1_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_QDR_M0_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0                                      'h00000AEC
`define CH1_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_QDR_M0_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0                                      'h00000AF0
`define CH1_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_QDR_M1_R0_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0                                      'h00000AF4
`define CH1_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P1                                   1
`define CH1_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0__PIPE_EN_P0                                   0
`define CH1_CA_SWI_DQS_TX_QDR_M1_R1_CFG_0___POR                              32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0                                'h00000AF8
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P1                               4
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0__X_SEL_P0                               0
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0                                'h00000AFC
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P1                               4
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0__X_SEL_P0                               0
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M0_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0                                'h00000B00
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P1                               4
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0__X_SEL_P0                               0
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R0_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0                                'h00000B04
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P1                               4
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0__X_SEL_P0                               0
`define CH1_CA_SWI_DQS_TX_QDR_X_SEL_M1_R1_CFG_0___POR                        32'h00000000

`define CH1_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0                                     'h00000B08
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__GEAR                                      7:6
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__EN                                          8
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R0_CFG_0___POR                             32'h00000100

`define CH1_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0                                     'h00000B0C
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__GEAR                                      7:6
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__EN                                          8
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQS_TX_LPDE_M0_R1_CFG_0___POR                             32'h00000100

`define CH1_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0                                     'h00000B10
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__GEAR                                      7:6
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__EN                                          8
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R0_CFG_0___POR                             32'h00000100

`define CH1_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0                                     'h00000B14
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__GEAR                                      7:6
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__EN                                          8
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0__CTRL_BIN                                  5:0
`define CH1_CA_SWI_DQS_TX_LPDE_M1_R1_CFG_0___POR                             32'h00000100

`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0                                          'h00000B18
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__TX_IMPD                                        8:6
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__SW_OVR                                           5
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__RX_IMPD                                       11:9
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_T                                       4
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_VAL_C                                       3
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0__OVRD_SEL                                       2:0
`define CH1_CA_SWI_DQS_TX_IO_M0_CFG_0___POR                                  32'h00000041

`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0                                          'h00000B1C
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__TX_IMPD                                        8:6
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__SW_OVR                                           5
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__RX_IMPD                                       11:9
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_T                                       4
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_VAL_C                                       3
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0__OVRD_SEL                                       2:0
`define CH1_CA_SWI_DQS_TX_IO_M1_CFG_0___POR                                  32'h00000041

`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG                                     'h00000B20
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__SE_MODE                                    13
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__PCAL                                     10:5
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__NCAL                                      4:0
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__LPBK_EN                                    12
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG__BS_EN                                      11
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R0_CFG___POR                             32'h00000001

`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG                                     'h00000B24
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__SE_MODE                                    13
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__PCAL                                     10:5
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__NCAL                                      4:0
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__LPBK_EN                                    12
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG__BS_EN                                      11
`define CH1_CA_SWI_DQS_TX_IO_CMN_M0_R1_CFG___POR                             32'h00000001

`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG                                     'h00000B28
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__SE_MODE                                    13
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__PCAL                                     10:5
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__NCAL                                      4:0
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__LPBK_EN                                    12
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG__BS_EN                                      11
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R0_CFG___POR                             32'h00000001

`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG                                     'h00000B2C
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__SE_MODE                                    13
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__PCAL                                     10:5
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__NCAL                                      4:0
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__LPBK_EN                                    12
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG__BS_EN                                      11
`define CH1_CA_SWI_DQS_TX_IO_CMN_M1_R1_CFG___POR                             32'h00000001
