/*
:name: class_test_5
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
virtual class automatic Foo; endclass