/*
:name: class_member_test_19
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function void subr(bool x[N]);
endclass