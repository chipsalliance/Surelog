/*
:name: 22.12--line-illegal-5
:description: Missing filename 
:should_fail_because: filename is missing 
:tags: 22.12
:type: preprocessing
*/
`line 1
