/*
:name: class_test_33
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class zzxy;
extern function void set_port(dbg_pkg::analysis_port app);
endclass