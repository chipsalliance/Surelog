/*
:name: empty_test_1
:description: Test
:should_fail: 0
:tags: 5.3 5.4
*/
    