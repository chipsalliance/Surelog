/*
:name: parameter_type
:description: parameter type tests
:should_fail: 0
:tags: 6.20.3
*/
module top #(type T = real);
endmodule
