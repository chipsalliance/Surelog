

package bp_common_pkg;

  `include "bp_common_me_if.vh"

endpackage : bp_common_pkg

