/*
:name: parameter_real
:description: parameter with real value test
:tags: 6.20.2
*/
module top();
	parameter p = 4.76;
endmodule
