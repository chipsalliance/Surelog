/*
:name: timescale-directive
:description: Set timescale
:tags: 5.6.4
*/

`timescale 1 ns / 1 ps

module ts();
endmodule
