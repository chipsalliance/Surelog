/*
:name: realtime
:description: realtime type tests
:should_fail: 0
:tags: 6.12
*/
module top();
	realtime a = 0.5;
endmodule
