`include "tb_env.sv"

program test;

tb_env env = new;

initial
begin
   env.cfg.perf_on = 1;
   env.run();
end

endprogram
