package toto1_1;





class blah1_7;
endclass












class blah2_21;
endclass





`include "middle.v"









class blah3_38;
endclass








endpackage




package toto2_53;





class blah21_59;
endclass




class blah22_65;
endclass




endpackage



module inb_75 ();
endmodule


package toto3_79;


endpackage

module gap2_84();
endmodule





























module gap3_115();
endmodule


package toto4_119;

class blah31_121;
endclass












class blah31_135;
endclass















class blah32_152;
endclass













class blah31_167;
endclass





endpackage






module gap4_181();












endmodule
