`define DDR_ANA_CKE_DRVR_LPBK_BS_EN_FIELD        11
`define DDR_ANA_CKE_DRVR_LPBK_LPBK_EN_FIELD      12
