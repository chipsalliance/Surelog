mem[   0] = 32'he3a00000;
mem[   1] = 32'he13ff000;
mem[   2] = 32'he3a00001;
mem[   3] = 32'hee030f10;
mem[   4] = 32'he3a00001;
mem[   5] = 32'hee020f10;
mem[   6] = 32'he3a0d801;
mem[   7] = 32'heb000000;
mem[   8] = 32'heafffffe;
mem[   9] = 32'he3a01201;
mem[  10] = 32'he3a03002;
mem[  11] = 32'he59f0084;
mem[  12] = 32'he92d40f0;
mem[  13] = 32'he3a02003;
mem[  14] = 32'he5813000;
mem[  15] = 32'he3a0c001;
mem[  16] = 32'he3a03000;
mem[  17] = 32'he1a06001;
mem[  18] = 32'he1a012a3;
mem[  19] = 32'he7901101;
mem[  20] = 32'he203401f;
mem[  21] = 32'he011141c;
mem[  22] = 32'h1a00000e;
mem[  23] = 32'he5862000;
mem[  24] = 32'he1a01082;
mem[  25] = 32'he3110001;
mem[  26] = 32'h0a000008;
mem[  27] = 32'he2414003;
mem[  28] = 32'he1a050a4;
mem[  29] = 32'he355003f;
mem[  30] = 32'h8a000006;
mem[  31] = 32'he1a04324;
mem[  32] = 32'he7907104;
mem[  33] = 32'he205501f;
mem[  34] = 32'he187551c;
mem[  35] = 32'he7805104;
mem[  36] = 32'he0811002;
mem[  37] = 32'heafffff2;
mem[  38] = 32'he2833001;
mem[  39] = 32'he3530040;
mem[  40] = 32'he2822002;
mem[  41] = 32'h1affffe7;
mem[  42] = 32'he3a00000;
mem[  43] = 32'he3a03201;
mem[  44] = 32'he5830000;
mem[  45] = 32'he8bd80f0;
mem[  46] = 32'h000000bc;
mem[  47] = 32'h00000000;
mem[  48] = 32'h00000000;
