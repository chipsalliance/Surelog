/*
:name: string
:description: string type tests
:should_fail: 0
:tags: 6.16
*/
module top();
	string a;
endmodule
