HAL/vmm_hw_rtl.sv