/*
:name: class_test_59
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class pp_class;
`ifdef DEBUGGER
`endif
endclass