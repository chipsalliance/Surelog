/*
:name: stop_task
:description: $stop test
:should_fail: 0
:tags: 20.2
*/
module top();

initial
	$stop;

endmodule
