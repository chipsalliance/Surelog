module dut();

   top top();

   
endmodule

