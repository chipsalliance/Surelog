/*
:name: typedef_test_7
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef struct { int i, j, k; bool b, c, d; } mystruct;