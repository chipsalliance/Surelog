/*
:name: class_test_4
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
virtual class Foo; endclass