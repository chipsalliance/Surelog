/*
:name: enum_test_0
:description: Test
:tags: 6.19
*/
typedef enum myenum_fwd;