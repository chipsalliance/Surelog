module simple_if (logic a);

endmodule
