/*
:name: 22.4--include_basic
:description: Test
:should_fail: 0
:tags: 22.4
:type: preprocessing parsing
*/
`include <dummy_include.sv>
module top ();
endmodule
