/*
:name: queues-basic
:description: Test queues support
:should_fail: 0
:tags: 7.10
*/
module top ();

int q[$];

endmodule
