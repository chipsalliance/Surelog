/*
:name: parameter_port_list
:description: parameter port list tests
:should_fail: 0
:tags: 6.20.2
*/
module top #(p = 12);
endmodule
