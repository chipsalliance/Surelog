/*
:name: class_member_test_26
:description: Test
:tags: 8.3
*/
class myclass;
pure virtual function integer subroutine;
pure virtual function integer compute(int a, bit b);
endclass