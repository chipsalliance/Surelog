/*
:name: class_test_24
:description: Test
:tags: 6.15 8.3
*/
class Foo implements Bar, Blah, Baz; endclass