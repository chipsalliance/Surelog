`define DDR_ANA_SA_2PH_OVR_EN_0_180_RANGE            0
`define DDR_ANA_SA_2PH_CAL_EN_0_180_RANGE            1
`define DDR_ANA_SA_2PH_SW_OVR_RANGE                  4
