/*
:name: associative-arrays-string
:description: Test associative arrays support
:tags: 7.8.2 7.8
*/
module top ();

int arr [ string ];

endmodule
