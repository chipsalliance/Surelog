/*
:name: desc_test_8
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
package mypkg;
endpackage
`endif
