/*
module dut (input i, output o);
  wire i;
  reg o;
  assign o = i;
endmodule
*/

module dut (i, o);
  input i;
  output o;
  wire i;
  reg o;
  assign o = i;
endmodule
