// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: desc_test_10
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef FPGA
`ifndef DEBUGGER
interface myinterface;
endinterface
`endif
`endif
