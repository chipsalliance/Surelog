/*
:name: associative-arrays-class
:description: Test associative arrays support
:tags: 7.8.3 7.8
*/
module top ();

class C;
    int x;
endclass

int arr [ C ];

endmodule
