/*
:name: class_member_test_48
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
virtual splinterface grinterface;
virtual interface foo_if bar_if;
endclass