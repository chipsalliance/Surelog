/*
:name: typedef_test_5
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef union { int i; bool b; } bint;