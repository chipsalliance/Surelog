/*
:name: typedef_test_10
:description: Test
:tags: 6.18
*/
typedef bit data_t;

typedef data_t my_array_t [ * ];
