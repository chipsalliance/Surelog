/*
:name: preproc_test_9
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`define LONG_MACRO(
    a, b, c)
