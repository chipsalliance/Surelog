/*
:name: defs 
:description: Utility for testing `include directive
:should_fail: 0
:tags: 22.4
*/

`define define_var "define_var"
`define TWO_PLUS_TWO 5
