/*
:name: preproc_test_0
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`define TRUTH
