`define DDR_ANA_SA_4PH_EN_0_180_RANGE                0
`define DDR_ANA_SA_4PH_CAL_EN_0_180_RANGE            1
`define DDR_ANA_SA_4PH_EN_90_270_RANGE               2
`define DDR_ANA_SA_4PH_CAL_EN_90_270_RANGE           3
`define DDR_ANA_SA_4PH_SW_OVR_RANGE                  4
