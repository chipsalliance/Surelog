/*
:name: class_member_test_45
:description: Test
:tags: 8.3
*/
class constructible;
extern function new();
endclass