/*
:name: desc_test_8
:description: Test
:type: preprocessing
:should_fail: 0
:tags: 5.6.4
*/
`ifdef DEBUGGER
package mypkg;
endpackage
`endif
