// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: typedef_test_16
:description: Test
:tags: 6.18
*/
typedef struct packed {
  logic [4:0] some_member;
} mystruct_t;

module test;
endmodule
