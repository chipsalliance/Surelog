


/*


  Leaf


*/


class leaf_13;
endclass

