// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: string-basic
:description: Basic string example
:tags: 5.9 5.3
*/
module top();

  initial begin;
    $display("one line");
  end

endmodule
