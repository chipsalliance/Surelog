module top(b);
input b;
reg [31:0] reg_32 = 32'bX;
endmodule

