// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: class_test_56
:description: Test
:tags: 6.15 8.3
*/
typedef int data_type_or_module_type;

class Driver;
  data_type_or_module_type foo1;
  data_type_or_module_type foo2 = 1'b1;
  data_type_or_module_type foo3, foo4;
  data_type_or_module_type foo5 = 5, foo6 = 6;
endclass

module test;
endmodule
