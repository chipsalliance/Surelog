module add(
  input [31:0] a,b,
  output signed [31:0] sum
);
assign sum = a + b ;
endmodule // add
