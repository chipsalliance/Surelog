// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: string_tolower
:description: string.tolower()  tests
:tags: 6.16.5
*/
module top();
	string a = "Test";
	string b = a.tolower();
endmodule
