`define DDR_ANA_PROG_DLY_SE_CTRL_BIN_RANGE                5:0
`define DDR_ANA_PROG_DLY_SE_GEAR_RANGE                    7:6
`define DDR_ANA_PROG_DLY_SE_EN_RANGE                      8

