/*
:name: class_member_test_29
:description: Test
:tags: 8.3
*/
class myclass;
function void shifter;
  for ( ; shft_idx < n_bits; ) begin
  end
endfunction
endclass