/*
:name: realtime_task
:description: $realtime test
:should_fail: 0
:tags: 20.3
*/
module top();

initial
	$display($realtime);

endmodule
