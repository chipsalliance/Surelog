/*
:name: class_member_test_6
:description: Test
:tags: 8.3
*/
class myclass;
extern protected task subtask(arg_type arg);
endclass