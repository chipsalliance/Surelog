module top();
 
    (* keep , syn_keep *) wire       [31:0]   execute_RS1 /* synthesis syn_keep = 1 */ ;
    (* async_reg = "true" *) reg                 system_rsp_valid;
    (* anyconst *)	reg	[LGFLEN:0]	fw_first_addr;

endmodule

