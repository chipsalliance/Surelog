`define DDR_ANA_DQ_DRVR_LPBK_OVRD_SEL_FIELD    2:0
`define DDR_ANA_DQ_DRVR_LPBK_OVRD_VAL_FIELD      3
`define DDR_ANA_DQ_DRVR_LPBK_RSVD_FIELD          4
`define DDR_ANA_DQ_DRVR_LPBK_SW_OVR_FIELD        5
`define DDR_ANA_DQ_DRVR_LPBK_TX_IMPD_FIELD     8:6
`define DDR_ANA_DQ_DRVR_LPBK_RX_IMPD_FIELD    11:9
