module badtop();
   import pkg2::*;
   mod m();
   top p();
   
endmodule
