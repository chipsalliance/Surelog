/*
:name: desc_test_5
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
`elsif BORED
`elsif MORE_BORED
`else
`endif
