/*
:name: string_bintoa
:description: string.bintoa()  tests
:tags: 6.16.14
*/
module top();
	string a;
	initial
		a.bintoa(12);
endmodule
