module top();

(* preserve *) reg my_reg1, my_reg2;

reg no_attrib;

endmodule // top
