/*
:name: class_test_17
:description: Test
:tags: 6.15 8.3
*/
class Foo #(type IFType=virtual x_if);
endclass