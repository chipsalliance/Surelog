/*
:name: class_test_31
:description: Test
:tags: 6.15 8.3
*/
typedef class myclass_fwd;