module top(output string o);
//string o;
   initial begin
      o = "abcd";
   end
endmodule
