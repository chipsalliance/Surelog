/*
:name: chandle
:description: chandle type tests
:should_fail: 0
:tags: 6.14
*/
module top();
	chandle a;
endmodule
