module top (input i, output o);
wire i;
reg o;
assign o = i;
endmodule


