/*
:name: dummy_include
:description: Utility for testing `include directive
:should_fail: 0
:tags: 22.4
*/
