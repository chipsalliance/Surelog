/*
:name: 22.12--line-illegal-3
:description: `line number parameter test
:should_fail_because: the number parameter shall be a positive integer that specifies the new line number
:tags: 22.12
:type: preprocessing
*/
`line -12 "somefile" 3
