module dut;
   chandle c;
endmodule
