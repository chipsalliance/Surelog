// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.10--celldefine-basic-1
:description: Test
:tags: 22.10
:type: preprocessing
*/
`celldefine
`endcelldefine
