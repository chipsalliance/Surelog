module top(b);
input b;
wire a = 100_000.0;
endmodule

