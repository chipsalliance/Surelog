// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: typedef_test_11
:description: Test
:tags: 6.18
*/
typedef bit data_t;

typedef data_t my_array_t [bit];

module test;
endmodule
