/*
:name: shortreal
:description: shortreal type tests
:should_fail: 0
:tags: 6.12
*/
module top();
	shortreal a = 0.5;
endmodule
