/*
:name: 22.3--resetall_basic
:description: Test
:should_fail: 0
:tags: 22.3
:type: preprocessing parsing
*/
`resetall
module top ();
endmodule
