module top();

	

	
endmodule