/*
:name: class_member_test_21
:description: Test
:tags: 8.3
*/
class myclass;
extern function sometype #(N+1) subr(ducktype #(3) x);
endclass