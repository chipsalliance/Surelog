/*
:name: 22.12--line-complex
:description: Test
:should_fail: 0
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 2
`line 123 "someother" 1
`line 8273 "somefile" 0
`resetall
`line 5 "foo" 2
