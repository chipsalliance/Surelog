/*
:name: 22.12--line-illegal-2
:description: filename parameter test
:should_fail_because: the filename parameter shall be a string literal
:tags: 22.12
:type: preprocessing
*/
`line 1 somefile 2
