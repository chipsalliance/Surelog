/*
:name: typedef_test_8__bad
:description: Test
:should_fail_because: some_other_type is not defined
:tags: 6.18
:type: simulation
*/
typedef some_other_type myalias;
