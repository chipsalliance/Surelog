module CELL1 (); 
endmodule

