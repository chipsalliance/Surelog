// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: arrays
:description: Basic arrays test
:tags: 5.11
*/
module top();
  int n[1:2][1:3] = '{'{0,1,2},'{3{4}}};
endmodule
