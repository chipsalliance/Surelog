/*
:name: module_definition
:description: module definition test
:should_fail: 0
:tags: 23.2
*/
module top();

endmodule
