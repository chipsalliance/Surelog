/*
:name: empty_test_2
:description: Test
:type: preprocessing
:tags: 5.3 5.4
*/
			