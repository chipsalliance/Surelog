/*
:name: nettype
:description: user-defined nettype tests
:tags: 6.6.7
*/
module top();
	nettype real real_net;
endmodule
