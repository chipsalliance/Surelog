/*
:name: display_task
:description: $display test
:tags: 21.2
:type: simulation parsing
*/
module top();

initial begin
	int val = 1234;
	$display(val);
end

endmodule
