/*
:name: typedef_test_3
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef reg[1:0] quartet[1:0];