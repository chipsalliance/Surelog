/*
:name: class_test_62
:description: Test
:tags: 6.15 8.3
*/
class pp_class;
  int num_packets;
`ifdef DEBUGGER
`endif
  int router_size;
endclass