/*
:name: time_task
:description: $time test
:tags: 20.3
*/
module top();

initial
	$display($time);

endmodule
