/*
 * Copyright (c) 2001 Stephen Williams (steve@icarus.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

/*
 * This problem shows the case of a function with no input ports,
 * and also a function with a parameter (not a port).
 */

module main;

   function [3:0] test;

      parameter a = 3;
      reg [a:0] out;

      begin
	 out = a;
	 test[3:0] = out[3:0];
      end

   endfunction

   reg [3:0] tmp;
   initial begin
      tmp = test();
      if (tmp !== 4'b0011) begin
	 $display("FAILED -- tmp == %b", tmp);
	 $finish;
      end

      $display("PASSED");
   end

endmodule // main

