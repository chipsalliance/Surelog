/*
:name: string
:description: string type tests
:tags: 6.16
*/
module top();
	string a;
endmodule
