/*
:name: class_member_test_34
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
virtual function integer subroutine;
  input a;
  subroutine = a+42;
endfunction
endclass