/*
:name: 22.12--line-illegal-1
:description: `line test
:should_fail_because: the level parameter shall be 0, 1, or 2
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile" 3
