

module top();
  import pack::*;
  initial begin
    $error("");
  end
  
  
endmodule
