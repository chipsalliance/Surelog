/*
:name: class_test_16
:description: Test
:tags: 6.15 8.3
*/
class Foo #(IFType=virtual x_if);
endclass