/*
:name: 22.5.1--define_expansion_23
:description: Test
:should_fail: 1
:tags: 22.5.1
:type: preprocessing
*/
`define define "illegal"
