/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  IC6.1.8-64b.500.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 17877
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_prog_dly_se_4g_small_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_sim_lib, Cell -
//wphy_prog_dly_se_4g_small_tb, View - schematic
// LAST TIME SAVED: Feb  1 21:48:21 2021
// NETLIST TIME: Feb  1 23:42:58 2021
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wphy_ips_lib", "wphy_prog_dly_se_4g" "systemVerilog"

`timescale 1ps/1fs

`endif //SYNTHESIS 
module wphy_prog_dly_se_4g_small ( outb,   ena, gear, i_ctrl, in 
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


  input  [5:0] i_ctrl;
  input in;
  input  [1:0] gear;
  
  input ena;
  output outb;
  
`ifdef SYNTHESIS
`else 

  reg  outb_int = 1'b0;
  real delay_total  = 0.0;
  reg assert_en=1'b0;
  real posedge_in=0.0;
  real posedge_in_pre=0.0;
  real period_in=1000.0;
  reg tmp_flag=0;
  wire pwr_ok;

  assign pwr_ok = ~vss & vdda;

  assign signals_ok = ((^i_ctrl)!==1'bz) && ((^i_ctrl)!==1'bx) &&  
                      ((^gear)!==1'bz) && ((^gear)!==1'bx) ;


  initial begin
   if ($value$plusargs("WPHY_ANA_ASSERT_EN=%f", assert_en)) begin
      assert_en=assert_en;
   end
  end

  initial begin
    case(gear)
      //0: delay_total = 40+6*i_ctrl;
      1: delay_total = 39+3*i_ctrl;
      2: delay_total = 27+2*i_ctrl;
      3: delay_total = 22+1*i_ctrl;
      default: delay_total = 0.0;
    endcase

    if(ena)
      outb_int <=  #(delay_total) ~in;
    else
      outb_int <= 1'bz;

  end

  //assign en_int = ena | (|gear);

  always @(i_ctrl,gear) begin
    case(gear)
      //0: delay_total = 40+6*i_ctrl;
      1: delay_total = 39+3*i_ctrl;
      2: delay_total = 27+2*i_ctrl;
      3: delay_total = 22+1*i_ctrl;
      default: delay_total = 0.0;
    endcase
  end

  always @(in,ena,delay_total) begin
    #0;
    if(ena)
      outb_int <=  #(delay_total) ~in;
    else
      outb_int <= 1'b1;
  end

  assign outb = (pwr_ok & signals_ok & (~ena | gear!==2'b00)) ? (ena) ? outb_int : 1'b1 : 1'bx;


  always @(posedge in) begin
      posedge_in = $realtime;
      period_in = posedge_in - posedge_in_pre; 
      posedge_in_pre = posedge_in;
  
      if(period_in<delay_total & ena & assert_en) begin
        $display("WPHY_ANA_ERROR: input period to slow for delay selected in %m at %t",$realtime);
        tmp_flag=1;
      end
      else begin
        tmp_flag=0;
        period_in=1000.0;
      end
  end

  always @(in,ena) begin
   #0;
     if(ena) begin
       if(gear===2'b00 & assert_en) begin
          $display("WPHY_ANA_ERROR: Gear=0 is not allowed for small programmable delay in %m at %t",$realtime);
       end
     end

  end


`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
`endif //SYNTHESIS
