/*
:name: 22.10--celldefine-basic-1
:description: Test
:tags: 22.10
:type: preprocessing
*/
`celldefine
`endcelldefine
