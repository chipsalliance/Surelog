/*
:name: desc_test_0
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifdef DEBUGGER
`endif
