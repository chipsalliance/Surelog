module omsp_alu(alu_out, alu_out_add, alu_stat, alu_stat_wr, dbg_halt_st, exec_cycle, inst_alu, inst_bw, inst_jmp, inst_so, op_dst, op_src, status);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire N;
  wire Z;
  wire [16:0] alu_add;
  output [15:0] alu_out;
  output [15:0] alu_out_add;
  wire [16:0] alu_out_nxt;
  wire [16:0] alu_shift;
  output [3:0] alu_stat;
  output [3:0] alu_stat_wr;
  wire [16:0] alu_swpb;
  wire [16:0] alu_sxt;
  input dbg_halt_st;
  input exec_cycle;
  input [11:0] inst_alu;
  input inst_bw;
  input [7:0] inst_jmp;
  input [7:0] inst_so;
  input [15:0] op_dst;
  wire [16:0] op_dst_in;
  input [15:0] op_src;
  input [3:0] status;
  \$_AND_  _0785_ (
    .A(exec_cycle),
    .B(inst_alu[0]),
    .Y(_0783_)
  );
  \$_XOR_  _0786_ (
    .A(_0783_),
    .B(op_src[0]),
    .Y(_0784_)
  );
  \$_INV_  _0787_ (
    .A(_0784_),
    .Y(_0000_)
  );
  \$_INV_  _0788_ (
    .A(status[2]),
    .Y(_0001_)
  );
  \$_AND_  _0789_ (
    .A(_0001_),
    .B(inst_jmp[4]),
    .Y(_0002_)
  );
  \$_INV_  _0790_ (
    .A(status[0]),
    .Y(_0003_)
  );
  \$_AND_  _0791_ (
    .A(inst_jmp[3]),
    .B(_0003_),
    .Y(_0004_)
  );
  \$_OR_  _0792_ (
    .A(_0004_),
    .B(_0002_),
    .Y(_0005_)
  );
  \$_AND_  _0793_ (
    .A(inst_jmp[0]),
    .B(status[1]),
    .Y(_0006_)
  );
  \$_AND_  _0794_ (
    .A(inst_jmp[2]),
    .B(status[0]),
    .Y(_0007_)
  );
  \$_INV_  _0795_ (
    .A(status[1]),
    .Y(_0008_)
  );
  \$_AND_  _0796_ (
    .A(_0008_),
    .B(inst_jmp[1]),
    .Y(_0009_)
  );
  \$_OR_  _0797_ (
    .A(_0009_),
    .B(_0007_),
    .Y(_0010_)
  );
  \$_OR_  _0798_ (
    .A(_0010_),
    .B(_0006_),
    .Y(_0011_)
  );
  \$_OR_  _0799_ (
    .A(_0011_),
    .B(_0005_),
    .Y(_0012_)
  );
  \$_XOR_  _0800_ (
    .A(status[3]),
    .B(status[2]),
    .Y(_0013_)
  );
  \$_MUX_  _0801_ (
    .A(inst_jmp[6]),
    .B(inst_jmp[5]),
    .S(_0013_),
    .Y(_0014_)
  );
  \$_OR_  _0802_ (
    .A(_0014_),
    .B(_0012_),
    .Y(_0015_)
  );
  \$_OR_  _0803_ (
    .A(_0015_),
    .B(_0000_),
    .Y(_0016_)
  );
  \$_XOR_  _0804_ (
    .A(_0016_),
    .B(op_dst[0]),
    .Y(_0017_)
  );
  \$_INV_  _0805_ (
    .A(_0017_),
    .Y(alu_add[0])
  );
  \$_INV_  _0806_ (
    .A(inst_jmp[4]),
    .Y(_0018_)
  );
  \$_OR_  _0807_ (
    .A(status[2]),
    .B(_0018_),
    .Y(_0019_)
  );
  \$_INV_  _0808_ (
    .A(inst_jmp[3]),
    .Y(_0020_)
  );
  \$_OR_  _0809_ (
    .A(_0020_),
    .B(status[0]),
    .Y(_0021_)
  );
  \$_AND_  _0810_ (
    .A(_0021_),
    .B(_0019_),
    .Y(_0022_)
  );
  \$_INV_  _0811_ (
    .A(_0006_),
    .Y(_0023_)
  );
  \$_INV_  _0812_ (
    .A(inst_jmp[2]),
    .Y(_0024_)
  );
  \$_OR_  _0813_ (
    .A(_0024_),
    .B(_0003_),
    .Y(_0025_)
  );
  \$_INV_  _0814_ (
    .A(inst_jmp[1]),
    .Y(_0026_)
  );
  \$_OR_  _0815_ (
    .A(status[1]),
    .B(_0026_),
    .Y(_0027_)
  );
  \$_AND_  _0816_ (
    .A(_0027_),
    .B(_0025_),
    .Y(_0028_)
  );
  \$_AND_  _0817_ (
    .A(_0028_),
    .B(_0023_),
    .Y(_0029_)
  );
  \$_AND_  _0818_ (
    .A(_0029_),
    .B(_0022_),
    .Y(_0030_)
  );
  \$_INV_  _0819_ (
    .A(_0014_),
    .Y(_0031_)
  );
  \$_AND_  _0820_ (
    .A(_0031_),
    .B(_0030_),
    .Y(_0032_)
  );
  \$_INV_  _0821_ (
    .A(op_src[10]),
    .Y(_0033_)
  );
  \$_XOR_  _0822_ (
    .A(_0783_),
    .B(_0033_),
    .Y(_0034_)
  );
  \$_AND_  _0823_ (
    .A(inst_bw),
    .B(exec_cycle),
    .Y(_0035_)
  );
  \$_OR_  _0824_ (
    .A(_0035_),
    .B(_0034_),
    .Y(_0036_)
  );
  \$_INV_  _0825_ (
    .A(_0036_),
    .Y(_0037_)
  );
  \$_AND_  _0826_ (
    .A(_0037_),
    .B(_0032_),
    .Y(_0038_)
  );
  \$_INV_  _0827_ (
    .A(_0035_),
    .Y(_0039_)
  );
  \$_AND_  _0828_ (
    .A(_0039_),
    .B(op_dst[10]),
    .Y(_0040_)
  );
  \$_INV_  _0829_ (
    .A(_0040_),
    .Y(_0041_)
  );
  \$_XOR_  _0830_ (
    .A(_0041_),
    .B(_0038_),
    .Y(_0042_)
  );
  \$_INV_  _0831_ (
    .A(_0042_),
    .Y(_0043_)
  );
  \$_INV_  _0832_ (
    .A(op_src[9]),
    .Y(_0044_)
  );
  \$_XOR_  _0833_ (
    .A(_0783_),
    .B(_0044_),
    .Y(_0045_)
  );
  \$_OR_  _0834_ (
    .A(_0045_),
    .B(_0035_),
    .Y(_0046_)
  );
  \$_INV_  _0835_ (
    .A(_0046_),
    .Y(_0047_)
  );
  \$_AND_  _0836_ (
    .A(_0047_),
    .B(_0032_),
    .Y(_0048_)
  );
  \$_AND_  _0837_ (
    .A(_0039_),
    .B(op_dst[9]),
    .Y(_0049_)
  );
  \$_AND_  _0838_ (
    .A(_0049_),
    .B(_0048_),
    .Y(_0050_)
  );
  \$_INV_  _0839_ (
    .A(_0050_),
    .Y(_0051_)
  );
  \$_INV_  _0840_ (
    .A(_0049_),
    .Y(_0052_)
  );
  \$_XOR_  _0841_ (
    .A(_0052_),
    .B(_0048_),
    .Y(_0053_)
  );
  \$_INV_  _0842_ (
    .A(op_src[8]),
    .Y(_0054_)
  );
  \$_XOR_  _0843_ (
    .A(_0783_),
    .B(_0054_),
    .Y(_0055_)
  );
  \$_OR_  _0844_ (
    .A(_0055_),
    .B(_0035_),
    .Y(_0056_)
  );
  \$_INV_  _0845_ (
    .A(_0056_),
    .Y(_0057_)
  );
  \$_AND_  _0846_ (
    .A(_0057_),
    .B(_0032_),
    .Y(_0058_)
  );
  \$_AND_  _0847_ (
    .A(_0039_),
    .B(op_dst[8]),
    .Y(_0059_)
  );
  \$_AND_  _0848_ (
    .A(_0059_),
    .B(_0058_),
    .Y(_0060_)
  );
  \$_INV_  _0849_ (
    .A(_0060_),
    .Y(_0061_)
  );
  \$_INV_  _0850_ (
    .A(_0059_),
    .Y(_0062_)
  );
  \$_XOR_  _0851_ (
    .A(_0062_),
    .B(_0058_),
    .Y(_0063_)
  );
  \$_INV_  _0852_ (
    .A(op_src[7]),
    .Y(_0064_)
  );
  \$_XOR_  _0853_ (
    .A(_0783_),
    .B(_0064_),
    .Y(_0065_)
  );
  \$_INV_  _0854_ (
    .A(_0065_),
    .Y(_0066_)
  );
  \$_AND_  _0855_ (
    .A(_0066_),
    .B(_0032_),
    .Y(_0067_)
  );
  \$_AND_  _0856_ (
    .A(_0067_),
    .B(op_dst[7]),
    .Y(_0068_)
  );
  \$_INV_  _0857_ (
    .A(_0068_),
    .Y(_0069_)
  );
  \$_INV_  _0858_ (
    .A(op_dst[7]),
    .Y(_0070_)
  );
  \$_XOR_  _0859_ (
    .A(_0067_),
    .B(_0070_),
    .Y(_0071_)
  );
  \$_INV_  _0860_ (
    .A(op_src[6]),
    .Y(_0072_)
  );
  \$_XOR_  _0861_ (
    .A(_0783_),
    .B(_0072_),
    .Y(_0073_)
  );
  \$_INV_  _0862_ (
    .A(_0073_),
    .Y(_0074_)
  );
  \$_AND_  _0863_ (
    .A(_0074_),
    .B(_0032_),
    .Y(_0075_)
  );
  \$_AND_  _0864_ (
    .A(_0075_),
    .B(op_dst[6]),
    .Y(_0076_)
  );
  \$_INV_  _0865_ (
    .A(_0076_),
    .Y(_0077_)
  );
  \$_INV_  _0866_ (
    .A(op_dst[6]),
    .Y(_0078_)
  );
  \$_XOR_  _0867_ (
    .A(_0075_),
    .B(_0078_),
    .Y(_0079_)
  );
  \$_INV_  _0868_ (
    .A(op_src[5]),
    .Y(_0080_)
  );
  \$_XOR_  _0869_ (
    .A(_0783_),
    .B(_0080_),
    .Y(_0081_)
  );
  \$_INV_  _0870_ (
    .A(_0081_),
    .Y(_0082_)
  );
  \$_AND_  _0871_ (
    .A(_0082_),
    .B(_0032_),
    .Y(_0083_)
  );
  \$_AND_  _0872_ (
    .A(_0083_),
    .B(op_dst[5]),
    .Y(_0084_)
  );
  \$_INV_  _0873_ (
    .A(_0084_),
    .Y(_0085_)
  );
  \$_INV_  _0874_ (
    .A(op_dst[5]),
    .Y(_0086_)
  );
  \$_XOR_  _0875_ (
    .A(_0083_),
    .B(_0086_),
    .Y(_0087_)
  );
  \$_INV_  _0876_ (
    .A(op_src[4]),
    .Y(_0088_)
  );
  \$_XOR_  _0877_ (
    .A(_0783_),
    .B(_0088_),
    .Y(_0089_)
  );
  \$_INV_  _0878_ (
    .A(_0089_),
    .Y(_0090_)
  );
  \$_AND_  _0879_ (
    .A(_0090_),
    .B(_0032_),
    .Y(_0091_)
  );
  \$_AND_  _0880_ (
    .A(_0091_),
    .B(op_dst[4]),
    .Y(_0092_)
  );
  \$_INV_  _0881_ (
    .A(_0092_),
    .Y(_0093_)
  );
  \$_INV_  _0882_ (
    .A(op_dst[4]),
    .Y(_0094_)
  );
  \$_XOR_  _0883_ (
    .A(_0091_),
    .B(_0094_),
    .Y(_0095_)
  );
  \$_INV_  _0884_ (
    .A(op_src[3]),
    .Y(_0096_)
  );
  \$_XOR_  _0885_ (
    .A(_0783_),
    .B(_0096_),
    .Y(_0097_)
  );
  \$_INV_  _0886_ (
    .A(_0097_),
    .Y(_0098_)
  );
  \$_AND_  _0887_ (
    .A(_0098_),
    .B(_0032_),
    .Y(_0099_)
  );
  \$_AND_  _0888_ (
    .A(_0099_),
    .B(op_dst[3]),
    .Y(_0100_)
  );
  \$_INV_  _0889_ (
    .A(_0100_),
    .Y(_0101_)
  );
  \$_INV_  _0890_ (
    .A(op_dst[3]),
    .Y(_0102_)
  );
  \$_XOR_  _0891_ (
    .A(_0099_),
    .B(_0102_),
    .Y(_0103_)
  );
  \$_INV_  _0892_ (
    .A(op_dst[2]),
    .Y(_0104_)
  );
  \$_INV_  _0893_ (
    .A(op_src[2]),
    .Y(_0105_)
  );
  \$_XOR_  _0894_ (
    .A(_0783_),
    .B(_0105_),
    .Y(_0106_)
  );
  \$_INV_  _0895_ (
    .A(_0106_),
    .Y(_0107_)
  );
  \$_AND_  _0896_ (
    .A(_0107_),
    .B(_0032_),
    .Y(_0108_)
  );
  \$_INV_  _0897_ (
    .A(_0108_),
    .Y(_0109_)
  );
  \$_OR_  _0898_ (
    .A(_0109_),
    .B(_0104_),
    .Y(_0110_)
  );
  \$_XOR_  _0899_ (
    .A(_0108_),
    .B(_0104_),
    .Y(_0111_)
  );
  \$_INV_  _0900_ (
    .A(op_dst[1]),
    .Y(_0112_)
  );
  \$_XOR_  _0901_ (
    .A(_0783_),
    .B(op_src[1]),
    .Y(_0113_)
  );
  \$_INV_  _0902_ (
    .A(_0113_),
    .Y(_0114_)
  );
  \$_OR_  _0903_ (
    .A(_0114_),
    .B(_0015_),
    .Y(_0115_)
  );
  \$_OR_  _0904_ (
    .A(_0115_),
    .B(_0112_),
    .Y(_0116_)
  );
  \$_XOR_  _0905_ (
    .A(_0115_),
    .B(op_dst[1]),
    .Y(_0117_)
  );
  \$_INV_  _0906_ (
    .A(op_dst[0]),
    .Y(_0118_)
  );
  \$_OR_  _0907_ (
    .A(_0016_),
    .B(_0118_),
    .Y(_0119_)
  );
  \$_OR_  _0908_ (
    .A(_0119_),
    .B(_0117_),
    .Y(_0120_)
  );
  \$_AND_  _0909_ (
    .A(_0120_),
    .B(_0116_),
    .Y(_0121_)
  );
  \$_OR_  _0910_ (
    .A(_0121_),
    .B(_0111_),
    .Y(_0122_)
  );
  \$_AND_  _0911_ (
    .A(_0122_),
    .B(_0110_),
    .Y(_0123_)
  );
  \$_OR_  _0912_ (
    .A(_0123_),
    .B(_0103_),
    .Y(_0124_)
  );
  \$_AND_  _0913_ (
    .A(_0124_),
    .B(_0101_),
    .Y(_0125_)
  );
  \$_OR_  _0914_ (
    .A(_0125_),
    .B(_0095_),
    .Y(_0126_)
  );
  \$_AND_  _0915_ (
    .A(_0126_),
    .B(_0093_),
    .Y(_0127_)
  );
  \$_OR_  _0916_ (
    .A(_0127_),
    .B(_0087_),
    .Y(_0128_)
  );
  \$_AND_  _0917_ (
    .A(_0128_),
    .B(_0085_),
    .Y(_0129_)
  );
  \$_OR_  _0918_ (
    .A(_0129_),
    .B(_0079_),
    .Y(_0130_)
  );
  \$_AND_  _0919_ (
    .A(_0130_),
    .B(_0077_),
    .Y(_0131_)
  );
  \$_OR_  _0920_ (
    .A(_0131_),
    .B(_0071_),
    .Y(_0132_)
  );
  \$_AND_  _0921_ (
    .A(_0132_),
    .B(_0069_),
    .Y(_0133_)
  );
  \$_OR_  _0922_ (
    .A(_0133_),
    .B(_0063_),
    .Y(_0134_)
  );
  \$_AND_  _0923_ (
    .A(_0134_),
    .B(_0061_),
    .Y(_0135_)
  );
  \$_OR_  _0924_ (
    .A(_0135_),
    .B(_0053_),
    .Y(_0136_)
  );
  \$_AND_  _0925_ (
    .A(_0136_),
    .B(_0051_),
    .Y(_0137_)
  );
  \$_XOR_  _0926_ (
    .A(_0137_),
    .B(_0043_),
    .Y(_0138_)
  );
  \$_INV_  _0927_ (
    .A(_0138_),
    .Y(alu_add[10])
  );
  \$_INV_  _0928_ (
    .A(op_src[11]),
    .Y(_0139_)
  );
  \$_XOR_  _0929_ (
    .A(_0783_),
    .B(_0139_),
    .Y(_0140_)
  );
  \$_OR_  _0930_ (
    .A(_0140_),
    .B(_0035_),
    .Y(_0141_)
  );
  \$_INV_  _0931_ (
    .A(_0141_),
    .Y(_0142_)
  );
  \$_AND_  _0932_ (
    .A(_0142_),
    .B(_0032_),
    .Y(_0143_)
  );
  \$_AND_  _0933_ (
    .A(_0039_),
    .B(op_dst[11]),
    .Y(_0144_)
  );
  \$_INV_  _0934_ (
    .A(_0144_),
    .Y(_0145_)
  );
  \$_XOR_  _0935_ (
    .A(_0145_),
    .B(_0143_),
    .Y(_0146_)
  );
  \$_AND_  _0936_ (
    .A(_0040_),
    .B(_0038_),
    .Y(_0147_)
  );
  \$_INV_  _0937_ (
    .A(_0147_),
    .Y(_0148_)
  );
  \$_OR_  _0938_ (
    .A(_0137_),
    .B(_0042_),
    .Y(_0149_)
  );
  \$_AND_  _0939_ (
    .A(_0149_),
    .B(_0148_),
    .Y(_0150_)
  );
  \$_XOR_  _0940_ (
    .A(_0150_),
    .B(_0146_),
    .Y(alu_add[11])
  );
  \$_INV_  _0941_ (
    .A(op_src[12]),
    .Y(_0151_)
  );
  \$_XOR_  _0942_ (
    .A(_0783_),
    .B(_0151_),
    .Y(_0152_)
  );
  \$_OR_  _0943_ (
    .A(_0152_),
    .B(_0035_),
    .Y(_0153_)
  );
  \$_INV_  _0944_ (
    .A(_0153_),
    .Y(_0154_)
  );
  \$_AND_  _0945_ (
    .A(_0154_),
    .B(_0032_),
    .Y(_0155_)
  );
  \$_AND_  _0946_ (
    .A(_0039_),
    .B(op_dst[12]),
    .Y(_0156_)
  );
  \$_INV_  _0947_ (
    .A(_0156_),
    .Y(_0157_)
  );
  \$_XOR_  _0948_ (
    .A(_0157_),
    .B(_0155_),
    .Y(_0158_)
  );
  \$_AND_  _0949_ (
    .A(_0144_),
    .B(_0143_),
    .Y(_0159_)
  );
  \$_INV_  _0950_ (
    .A(_0159_),
    .Y(_0160_)
  );
  \$_OR_  _0951_ (
    .A(_0150_),
    .B(_0146_),
    .Y(_0161_)
  );
  \$_AND_  _0952_ (
    .A(_0161_),
    .B(_0160_),
    .Y(_0162_)
  );
  \$_XOR_  _0953_ (
    .A(_0162_),
    .B(_0158_),
    .Y(alu_add[12])
  );
  \$_INV_  _0954_ (
    .A(op_src[13]),
    .Y(_0163_)
  );
  \$_XOR_  _0955_ (
    .A(_0783_),
    .B(_0163_),
    .Y(_0164_)
  );
  \$_OR_  _0956_ (
    .A(_0164_),
    .B(_0035_),
    .Y(_0165_)
  );
  \$_INV_  _0957_ (
    .A(_0165_),
    .Y(_0166_)
  );
  \$_AND_  _0958_ (
    .A(_0166_),
    .B(_0032_),
    .Y(_0167_)
  );
  \$_AND_  _0959_ (
    .A(_0039_),
    .B(op_dst[13]),
    .Y(_0168_)
  );
  \$_INV_  _0960_ (
    .A(_0168_),
    .Y(_0169_)
  );
  \$_XOR_  _0961_ (
    .A(_0169_),
    .B(_0167_),
    .Y(_0170_)
  );
  \$_AND_  _0962_ (
    .A(_0156_),
    .B(_0155_),
    .Y(_0171_)
  );
  \$_INV_  _0963_ (
    .A(_0171_),
    .Y(_0172_)
  );
  \$_OR_  _0964_ (
    .A(_0162_),
    .B(_0158_),
    .Y(_0173_)
  );
  \$_AND_  _0965_ (
    .A(_0173_),
    .B(_0172_),
    .Y(_0174_)
  );
  \$_XOR_  _0966_ (
    .A(_0174_),
    .B(_0170_),
    .Y(alu_add[13])
  );
  \$_INV_  _0967_ (
    .A(op_src[14]),
    .Y(_0175_)
  );
  \$_XOR_  _0968_ (
    .A(_0783_),
    .B(_0175_),
    .Y(_0176_)
  );
  \$_OR_  _0969_ (
    .A(_0176_),
    .B(_0035_),
    .Y(_0177_)
  );
  \$_INV_  _0970_ (
    .A(_0177_),
    .Y(_0178_)
  );
  \$_AND_  _0971_ (
    .A(_0178_),
    .B(_0032_),
    .Y(_0179_)
  );
  \$_AND_  _0972_ (
    .A(_0039_),
    .B(op_dst[14]),
    .Y(_0180_)
  );
  \$_INV_  _0973_ (
    .A(_0180_),
    .Y(_0181_)
  );
  \$_XOR_  _0974_ (
    .A(_0181_),
    .B(_0179_),
    .Y(_0182_)
  );
  \$_AND_  _0975_ (
    .A(_0168_),
    .B(_0167_),
    .Y(_0183_)
  );
  \$_INV_  _0976_ (
    .A(_0183_),
    .Y(_0184_)
  );
  \$_OR_  _0977_ (
    .A(_0174_),
    .B(_0170_),
    .Y(_0185_)
  );
  \$_AND_  _0978_ (
    .A(_0185_),
    .B(_0184_),
    .Y(_0186_)
  );
  \$_XOR_  _0979_ (
    .A(_0186_),
    .B(_0182_),
    .Y(alu_add[14])
  );
  \$_INV_  _0980_ (
    .A(op_src[15]),
    .Y(_0187_)
  );
  \$_XOR_  _0981_ (
    .A(_0783_),
    .B(_0187_),
    .Y(_0188_)
  );
  \$_OR_  _0982_ (
    .A(_0188_),
    .B(_0035_),
    .Y(_0189_)
  );
  \$_INV_  _0983_ (
    .A(_0189_),
    .Y(_0190_)
  );
  \$_AND_  _0984_ (
    .A(_0190_),
    .B(_0032_),
    .Y(_0191_)
  );
  \$_AND_  _0985_ (
    .A(_0039_),
    .B(op_dst[15]),
    .Y(_0192_)
  );
  \$_INV_  _0986_ (
    .A(_0192_),
    .Y(_0193_)
  );
  \$_XOR_  _0987_ (
    .A(_0193_),
    .B(_0191_),
    .Y(_0194_)
  );
  \$_AND_  _0988_ (
    .A(_0180_),
    .B(_0179_),
    .Y(_0195_)
  );
  \$_INV_  _0989_ (
    .A(_0195_),
    .Y(_0196_)
  );
  \$_OR_  _0990_ (
    .A(_0186_),
    .B(_0182_),
    .Y(_0197_)
  );
  \$_AND_  _0991_ (
    .A(_0197_),
    .B(_0196_),
    .Y(_0198_)
  );
  \$_XOR_  _0992_ (
    .A(_0198_),
    .B(_0194_),
    .Y(alu_add[15])
  );
  \$_INV_  _0993_ (
    .A(_0119_),
    .Y(_0199_)
  );
  \$_XOR_  _0994_ (
    .A(_0199_),
    .B(_0117_),
    .Y(_0200_)
  );
  \$_INV_  _0995_ (
    .A(_0200_),
    .Y(alu_add[1])
  );
  \$_INV_  _0996_ (
    .A(_0111_),
    .Y(_0201_)
  );
  \$_XOR_  _0997_ (
    .A(_0121_),
    .B(_0201_),
    .Y(_0202_)
  );
  \$_INV_  _0998_ (
    .A(_0202_),
    .Y(alu_add[2])
  );
  \$_INV_  _0999_ (
    .A(_0103_),
    .Y(_0203_)
  );
  \$_XOR_  _1000_ (
    .A(_0123_),
    .B(_0203_),
    .Y(_0204_)
  );
  \$_INV_  _1001_ (
    .A(_0204_),
    .Y(alu_add[3])
  );
  \$_INV_  _1002_ (
    .A(_0095_),
    .Y(_0205_)
  );
  \$_XOR_  _1003_ (
    .A(_0125_),
    .B(_0205_),
    .Y(_0206_)
  );
  \$_INV_  _1004_ (
    .A(_0206_),
    .Y(alu_add[4])
  );
  \$_INV_  _1005_ (
    .A(_0087_),
    .Y(_0207_)
  );
  \$_XOR_  _1006_ (
    .A(_0127_),
    .B(_0207_),
    .Y(_0208_)
  );
  \$_INV_  _1007_ (
    .A(_0208_),
    .Y(alu_add[5])
  );
  \$_INV_  _1008_ (
    .A(_0079_),
    .Y(_0209_)
  );
  \$_XOR_  _1009_ (
    .A(_0129_),
    .B(_0209_),
    .Y(_0210_)
  );
  \$_INV_  _1010_ (
    .A(_0210_),
    .Y(alu_add[6])
  );
  \$_INV_  _1011_ (
    .A(_0071_),
    .Y(_0211_)
  );
  \$_XOR_  _1012_ (
    .A(_0131_),
    .B(_0211_),
    .Y(_0212_)
  );
  \$_INV_  _1013_ (
    .A(_0212_),
    .Y(alu_add[7])
  );
  \$_INV_  _1014_ (
    .A(_0063_),
    .Y(_0213_)
  );
  \$_XOR_  _1015_ (
    .A(_0133_),
    .B(_0213_),
    .Y(_0214_)
  );
  \$_INV_  _1016_ (
    .A(_0214_),
    .Y(alu_add[8])
  );
  \$_INV_  _1017_ (
    .A(_0053_),
    .Y(_0215_)
  );
  \$_XOR_  _1018_ (
    .A(_0135_),
    .B(_0215_),
    .Y(_0216_)
  );
  \$_INV_  _1019_ (
    .A(_0216_),
    .Y(alu_add[9])
  );
  \$_OR_  _1020_ (
    .A(inst_so[7]),
    .B(dbg_halt_st),
    .Y(_0217_)
  );
  \$_OR_  _1021_ (
    .A(_0217_),
    .B(inst_alu[3]),
    .Y(_0218_)
  );
  \$_AND_  _1022_ (
    .A(inst_alu[2]),
    .B(status[0]),
    .Y(_0219_)
  );
  \$_OR_  _1023_ (
    .A(_0219_),
    .B(inst_alu[1]),
    .Y(_0220_)
  );
  \$_AND_  _1024_ (
    .A(_0220_),
    .B(exec_cycle),
    .Y(_0221_)
  );
  \$_AND_  _1025_ (
    .A(_0221_),
    .B(alu_add[0]),
    .Y(_0222_)
  );
  \$_AND_  _1026_ (
    .A(_0222_),
    .B(alu_add[1]),
    .Y(_0223_)
  );
  \$_AND_  _1027_ (
    .A(_0223_),
    .B(alu_add[2]),
    .Y(_0224_)
  );
  \$_AND_  _1028_ (
    .A(_0224_),
    .B(alu_add[3]),
    .Y(_0225_)
  );
  \$_AND_  _1029_ (
    .A(_0225_),
    .B(alu_add[4]),
    .Y(_0226_)
  );
  \$_AND_  _1030_ (
    .A(_0226_),
    .B(alu_add[5]),
    .Y(_0227_)
  );
  \$_AND_  _1031_ (
    .A(_0227_),
    .B(alu_add[6]),
    .Y(_0228_)
  );
  \$_XOR_  _1032_ (
    .A(_0228_),
    .B(_0212_),
    .Y(_0229_)
  );
  \$_XOR_  _1033_ (
    .A(_0065_),
    .B(op_dst[7]),
    .Y(_0230_)
  );
  \$_AND_  _1034_ (
    .A(_0074_),
    .B(op_dst[6]),
    .Y(_0231_)
  );
  \$_XOR_  _1035_ (
    .A(_0073_),
    .B(op_dst[6]),
    .Y(_0232_)
  );
  \$_INV_  _1036_ (
    .A(_0232_),
    .Y(_0233_)
  );
  \$_AND_  _1037_ (
    .A(_0082_),
    .B(op_dst[5]),
    .Y(_0234_)
  );
  \$_XOR_  _1038_ (
    .A(_0081_),
    .B(op_dst[5]),
    .Y(_0235_)
  );
  \$_INV_  _1039_ (
    .A(_0235_),
    .Y(_0236_)
  );
  \$_AND_  _1040_ (
    .A(_0090_),
    .B(op_dst[4]),
    .Y(_0237_)
  );
  \$_AND_  _1041_ (
    .A(_0237_),
    .B(_0236_),
    .Y(_0238_)
  );
  \$_OR_  _1042_ (
    .A(_0238_),
    .B(_0234_),
    .Y(_0239_)
  );
  \$_AND_  _1043_ (
    .A(_0239_),
    .B(_0233_),
    .Y(_0240_)
  );
  \$_OR_  _1044_ (
    .A(_0240_),
    .B(_0231_),
    .Y(_0241_)
  );
  \$_XOR_  _1045_ (
    .A(_0241_),
    .B(_0230_),
    .Y(_0242_)
  );
  \$_INV_  _1046_ (
    .A(_0242_),
    .Y(_0243_)
  );
  \$_XOR_  _1047_ (
    .A(_0239_),
    .B(_0232_),
    .Y(_0244_)
  );
  \$_INV_  _1048_ (
    .A(_0244_),
    .Y(_0245_)
  );
  \$_XOR_  _1049_ (
    .A(_0237_),
    .B(_0235_),
    .Y(_0246_)
  );
  \$_INV_  _1050_ (
    .A(_0246_),
    .Y(_0247_)
  );
  \$_XOR_  _1051_ (
    .A(_0089_),
    .B(op_dst[4]),
    .Y(_0248_)
  );
  \$_INV_  _1052_ (
    .A(_0248_),
    .Y(_0249_)
  );
  \$_AND_  _1053_ (
    .A(_0098_),
    .B(op_dst[3]),
    .Y(_0250_)
  );
  \$_XOR_  _1054_ (
    .A(_0097_),
    .B(op_dst[3]),
    .Y(_0251_)
  );
  \$_INV_  _1055_ (
    .A(_0251_),
    .Y(_0252_)
  );
  \$_AND_  _1056_ (
    .A(_0107_),
    .B(op_dst[2]),
    .Y(_0253_)
  );
  \$_XOR_  _1057_ (
    .A(_0106_),
    .B(op_dst[2]),
    .Y(_0254_)
  );
  \$_INV_  _1058_ (
    .A(_0254_),
    .Y(_0255_)
  );
  \$_AND_  _1059_ (
    .A(_0113_),
    .B(op_dst[1]),
    .Y(_0256_)
  );
  \$_XOR_  _1060_ (
    .A(_0113_),
    .B(_0112_),
    .Y(_0257_)
  );
  \$_INV_  _1061_ (
    .A(_0257_),
    .Y(_0258_)
  );
  \$_AND_  _1062_ (
    .A(_0784_),
    .B(op_dst[0]),
    .Y(_0259_)
  );
  \$_AND_  _1063_ (
    .A(_0259_),
    .B(_0258_),
    .Y(_0260_)
  );
  \$_OR_  _1064_ (
    .A(_0260_),
    .B(_0256_),
    .Y(_0261_)
  );
  \$_AND_  _1065_ (
    .A(_0261_),
    .B(_0255_),
    .Y(_0262_)
  );
  \$_OR_  _1066_ (
    .A(_0262_),
    .B(_0253_),
    .Y(_0263_)
  );
  \$_AND_  _1067_ (
    .A(_0263_),
    .B(_0252_),
    .Y(_0264_)
  );
  \$_OR_  _1068_ (
    .A(_0264_),
    .B(_0250_),
    .Y(_0265_)
  );
  \$_XOR_  _1069_ (
    .A(_0263_),
    .B(_0251_),
    .Y(_0266_)
  );
  \$_INV_  _1070_ (
    .A(_0266_),
    .Y(_0267_)
  );
  \$_XOR_  _1071_ (
    .A(_0261_),
    .B(_0254_),
    .Y(_0268_)
  );
  \$_INV_  _1072_ (
    .A(_0268_),
    .Y(_0269_)
  );
  \$_XOR_  _1073_ (
    .A(_0259_),
    .B(_0257_),
    .Y(_0270_)
  );
  \$_INV_  _1074_ (
    .A(_0270_),
    .Y(_0271_)
  );
  \$_XOR_  _1075_ (
    .A(_0784_),
    .B(_0118_),
    .Y(_0272_)
  );
  \$_INV_  _1076_ (
    .A(_0272_),
    .Y(_0273_)
  );
  \$_AND_  _1077_ (
    .A(_0273_),
    .B(status[0]),
    .Y(_0274_)
  );
  \$_AND_  _1078_ (
    .A(_0274_),
    .B(_0271_),
    .Y(_0275_)
  );
  \$_AND_  _1079_ (
    .A(_0275_),
    .B(_0269_),
    .Y(_0276_)
  );
  \$_AND_  _1080_ (
    .A(_0276_),
    .B(_0267_),
    .Y(_0277_)
  );
  \$_XOR_  _1081_ (
    .A(_0277_),
    .B(_0265_),
    .Y(_0278_)
  );
  \$_XOR_  _1082_ (
    .A(_0276_),
    .B(_0266_),
    .Y(_0279_)
  );
  \$_XOR_  _1083_ (
    .A(_0275_),
    .B(_0268_),
    .Y(_0280_)
  );
  \$_XOR_  _1084_ (
    .A(_0274_),
    .B(_0270_),
    .Y(_0281_)
  );
  \$_AND_  _1085_ (
    .A(_0281_),
    .B(_0280_),
    .Y(_0282_)
  );
  \$_OR_  _1086_ (
    .A(_0282_),
    .B(_0279_),
    .Y(_0283_)
  );
  \$_XOR_  _1087_ (
    .A(_0283_),
    .B(_0278_),
    .Y(_0284_)
  );
  \$_INV_  _1088_ (
    .A(_0284_),
    .Y(_0285_)
  );
  \$_AND_  _1089_ (
    .A(_0285_),
    .B(_0249_),
    .Y(_0286_)
  );
  \$_AND_  _1090_ (
    .A(_0286_),
    .B(_0247_),
    .Y(_0287_)
  );
  \$_AND_  _1091_ (
    .A(_0287_),
    .B(_0245_),
    .Y(_0288_)
  );
  \$_XOR_  _1092_ (
    .A(_0288_),
    .B(_0243_),
    .Y(_0289_)
  );
  \$_INV_  _1093_ (
    .A(_0289_),
    .Y(_0290_)
  );
  \$_AND_  _1094_ (
    .A(_0066_),
    .B(op_dst[7]),
    .Y(_0291_)
  );
  \$_INV_  _1095_ (
    .A(_0230_),
    .Y(_0292_)
  );
  \$_AND_  _1096_ (
    .A(_0241_),
    .B(_0292_),
    .Y(_0293_)
  );
  \$_OR_  _1097_ (
    .A(_0293_),
    .B(_0291_),
    .Y(_0294_)
  );
  \$_AND_  _1098_ (
    .A(_0288_),
    .B(_0243_),
    .Y(_0295_)
  );
  \$_XOR_  _1099_ (
    .A(_0295_),
    .B(_0294_),
    .Y(_0296_)
  );
  \$_INV_  _1100_ (
    .A(_0296_),
    .Y(_0297_)
  );
  \$_XOR_  _1101_ (
    .A(_0287_),
    .B(_0245_),
    .Y(_0298_)
  );
  \$_XOR_  _1102_ (
    .A(_0286_),
    .B(_0246_),
    .Y(_0299_)
  );
  \$_INV_  _1103_ (
    .A(_0299_),
    .Y(_0300_)
  );
  \$_OR_  _1104_ (
    .A(_0300_),
    .B(_0298_),
    .Y(_0301_)
  );
  \$_AND_  _1105_ (
    .A(_0301_),
    .B(_0289_),
    .Y(_0302_)
  );
  \$_INV_  _1106_ (
    .A(_0302_),
    .Y(_0303_)
  );
  \$_AND_  _1107_ (
    .A(_0303_),
    .B(_0297_),
    .Y(_0304_)
  );
  \$_XOR_  _1108_ (
    .A(_0301_),
    .B(_0290_),
    .Y(_0305_)
  );
  \$_MUX_  _1109_ (
    .A(_0305_),
    .B(_0290_),
    .S(_0304_),
    .Y(_0306_)
  );
  \$_INV_  _1110_ (
    .A(inst_alu[10]),
    .Y(_0307_)
  );
  \$_INV_  _1111_ (
    .A(inst_bw),
    .Y(_0308_)
  );
  \$_MUX_  _1112_ (
    .A(_0064_),
    .B(_0187_),
    .S(_0308_),
    .Y(_0309_)
  );
  \$_MUX_  _1113_ (
    .A(_0309_),
    .B(_0003_),
    .S(inst_so[0]),
    .Y(_0310_)
  );
  \$_MUX_  _1114_ (
    .A(_0310_),
    .B(_0054_),
    .S(_0308_),
    .Y(_0311_)
  );
  \$_OR_  _1115_ (
    .A(_0311_),
    .B(_0307_),
    .Y(_0312_)
  );
  \$_AND_  _1116_ (
    .A(_0292_),
    .B(inst_alu[6]),
    .Y(_0313_)
  );
  \$_INV_  _1117_ (
    .A(_0313_),
    .Y(_0314_)
  );
  \$_INV_  _1118_ (
    .A(inst_alu[5]),
    .Y(_0315_)
  );
  \$_AND_  _1119_ (
    .A(_0065_),
    .B(_0070_),
    .Y(_0316_)
  );
  \$_OR_  _1120_ (
    .A(_0316_),
    .B(_0315_),
    .Y(_0317_)
  );
  \$_AND_  _1121_ (
    .A(_0291_),
    .B(inst_alu[4]),
    .Y(_0318_)
  );
  \$_INV_  _1122_ (
    .A(inst_alu[4]),
    .Y(_0319_)
  );
  \$_AND_  _1123_ (
    .A(_0315_),
    .B(_0319_),
    .Y(_0320_)
  );
  \$_INV_  _1124_ (
    .A(inst_alu[6]),
    .Y(_0321_)
  );
  \$_AND_  _1125_ (
    .A(_0307_),
    .B(_0321_),
    .Y(_0322_)
  );
  \$_INV_  _1126_ (
    .A(inst_so[1]),
    .Y(_0323_)
  );
  \$_INV_  _1127_ (
    .A(inst_so[3]),
    .Y(_0324_)
  );
  \$_AND_  _1128_ (
    .A(_0324_),
    .B(_0323_),
    .Y(_0325_)
  );
  \$_AND_  _1129_ (
    .A(_0325_),
    .B(_0322_),
    .Y(_0326_)
  );
  \$_AND_  _1130_ (
    .A(_0326_),
    .B(_0320_),
    .Y(_0327_)
  );
  \$_AND_  _1131_ (
    .A(_0327_),
    .B(_0066_),
    .Y(_0328_)
  );
  \$_AND_  _1132_ (
    .A(inst_so[1]),
    .B(op_src[15]),
    .Y(_0329_)
  );
  \$_AND_  _1133_ (
    .A(inst_so[3]),
    .B(op_src[7]),
    .Y(_0330_)
  );
  \$_OR_  _1134_ (
    .A(_0330_),
    .B(_0329_),
    .Y(_0331_)
  );
  \$_OR_  _1135_ (
    .A(_0331_),
    .B(_0328_),
    .Y(_0332_)
  );
  \$_OR_  _1136_ (
    .A(_0332_),
    .B(_0318_),
    .Y(_0333_)
  );
  \$_INV_  _1137_ (
    .A(_0333_),
    .Y(_0334_)
  );
  \$_AND_  _1138_ (
    .A(_0334_),
    .B(_0317_),
    .Y(_0335_)
  );
  \$_AND_  _1139_ (
    .A(_0335_),
    .B(_0314_),
    .Y(_0336_)
  );
  \$_AND_  _1140_ (
    .A(_0336_),
    .B(_0312_),
    .Y(_0337_)
  );
  \$_MUX_  _1141_ (
    .A(_0337_),
    .B(_0306_),
    .S(inst_alu[7]),
    .Y(_0338_)
  );
  \$_MUX_  _1142_ (
    .A(_0338_),
    .B(_0229_),
    .S(_0218_),
    .Y(_0339_)
  );
  \$_INV_  _1143_ (
    .A(_0339_),
    .Y(alu_out[7])
  );
  \$_AND_  _1144_ (
    .A(_0228_),
    .B(alu_add[7]),
    .Y(_0340_)
  );
  \$_AND_  _1145_ (
    .A(_0340_),
    .B(alu_add[8]),
    .Y(_0341_)
  );
  \$_AND_  _1146_ (
    .A(_0341_),
    .B(alu_add[9]),
    .Y(_0342_)
  );
  \$_AND_  _1147_ (
    .A(_0342_),
    .B(alu_add[10]),
    .Y(_0343_)
  );
  \$_AND_  _1148_ (
    .A(_0343_),
    .B(alu_add[11]),
    .Y(_0344_)
  );
  \$_AND_  _1149_ (
    .A(_0344_),
    .B(alu_add[12]),
    .Y(_0345_)
  );
  \$_AND_  _1150_ (
    .A(_0345_),
    .B(alu_add[13]),
    .Y(_0346_)
  );
  \$_AND_  _1151_ (
    .A(_0346_),
    .B(alu_add[14]),
    .Y(_0347_)
  );
  \$_XOR_  _1152_ (
    .A(_0347_),
    .B(alu_add[15]),
    .Y(_0348_)
  );
  \$_XOR_  _1153_ (
    .A(_0192_),
    .B(_0189_),
    .Y(_0349_)
  );
  \$_AND_  _1154_ (
    .A(_0180_),
    .B(_0178_),
    .Y(_0350_)
  );
  \$_XOR_  _1155_ (
    .A(_0180_),
    .B(_0177_),
    .Y(_0351_)
  );
  \$_INV_  _1156_ (
    .A(_0351_),
    .Y(_0352_)
  );
  \$_AND_  _1157_ (
    .A(_0168_),
    .B(_0166_),
    .Y(_0353_)
  );
  \$_XOR_  _1158_ (
    .A(_0168_),
    .B(_0165_),
    .Y(_0354_)
  );
  \$_INV_  _1159_ (
    .A(_0354_),
    .Y(_0355_)
  );
  \$_AND_  _1160_ (
    .A(_0156_),
    .B(_0154_),
    .Y(_0356_)
  );
  \$_AND_  _1161_ (
    .A(_0356_),
    .B(_0355_),
    .Y(_0357_)
  );
  \$_OR_  _1162_ (
    .A(_0357_),
    .B(_0353_),
    .Y(_0358_)
  );
  \$_AND_  _1163_ (
    .A(_0358_),
    .B(_0352_),
    .Y(_0359_)
  );
  \$_OR_  _1164_ (
    .A(_0359_),
    .B(_0350_),
    .Y(_0360_)
  );
  \$_XOR_  _1165_ (
    .A(_0360_),
    .B(_0349_),
    .Y(_0361_)
  );
  \$_XOR_  _1166_ (
    .A(_0358_),
    .B(_0351_),
    .Y(_0362_)
  );
  \$_INV_  _1167_ (
    .A(_0362_),
    .Y(_0363_)
  );
  \$_XOR_  _1168_ (
    .A(_0356_),
    .B(_0354_),
    .Y(_0364_)
  );
  \$_INV_  _1169_ (
    .A(_0364_),
    .Y(_0365_)
  );
  \$_XOR_  _1170_ (
    .A(_0156_),
    .B(_0153_),
    .Y(_0366_)
  );
  \$_INV_  _1171_ (
    .A(_0366_),
    .Y(_0367_)
  );
  \$_AND_  _1172_ (
    .A(_0144_),
    .B(_0142_),
    .Y(_0368_)
  );
  \$_XOR_  _1173_ (
    .A(_0144_),
    .B(_0141_),
    .Y(_0369_)
  );
  \$_INV_  _1174_ (
    .A(_0369_),
    .Y(_0370_)
  );
  \$_AND_  _1175_ (
    .A(_0040_),
    .B(_0037_),
    .Y(_0371_)
  );
  \$_XOR_  _1176_ (
    .A(_0040_),
    .B(_0036_),
    .Y(_0372_)
  );
  \$_INV_  _1177_ (
    .A(_0372_),
    .Y(_0373_)
  );
  \$_AND_  _1178_ (
    .A(_0049_),
    .B(_0047_),
    .Y(_0374_)
  );
  \$_XOR_  _1179_ (
    .A(_0049_),
    .B(_0046_),
    .Y(_0375_)
  );
  \$_INV_  _1180_ (
    .A(_0375_),
    .Y(_0376_)
  );
  \$_AND_  _1181_ (
    .A(_0059_),
    .B(_0057_),
    .Y(_0377_)
  );
  \$_AND_  _1182_ (
    .A(_0377_),
    .B(_0376_),
    .Y(_0378_)
  );
  \$_OR_  _1183_ (
    .A(_0378_),
    .B(_0374_),
    .Y(_0379_)
  );
  \$_AND_  _1184_ (
    .A(_0379_),
    .B(_0373_),
    .Y(_0380_)
  );
  \$_OR_  _1185_ (
    .A(_0380_),
    .B(_0371_),
    .Y(_0381_)
  );
  \$_AND_  _1186_ (
    .A(_0381_),
    .B(_0370_),
    .Y(_0382_)
  );
  \$_OR_  _1187_ (
    .A(_0382_),
    .B(_0368_),
    .Y(_0383_)
  );
  \$_XOR_  _1188_ (
    .A(_0381_),
    .B(_0369_),
    .Y(_0384_)
  );
  \$_INV_  _1189_ (
    .A(_0384_),
    .Y(_0385_)
  );
  \$_XOR_  _1190_ (
    .A(_0379_),
    .B(_0372_),
    .Y(_0386_)
  );
  \$_INV_  _1191_ (
    .A(_0386_),
    .Y(_0387_)
  );
  \$_XOR_  _1192_ (
    .A(_0377_),
    .B(_0375_),
    .Y(_0388_)
  );
  \$_INV_  _1193_ (
    .A(_0388_),
    .Y(_0389_)
  );
  \$_XOR_  _1194_ (
    .A(_0059_),
    .B(_0056_),
    .Y(_0390_)
  );
  \$_INV_  _1195_ (
    .A(_0390_),
    .Y(_0391_)
  );
  \$_XOR_  _1196_ (
    .A(_0302_),
    .B(_0296_),
    .Y(_0392_)
  );
  \$_AND_  _1197_ (
    .A(_0392_),
    .B(_0391_),
    .Y(_0393_)
  );
  \$_AND_  _1198_ (
    .A(_0393_),
    .B(_0389_),
    .Y(_0394_)
  );
  \$_AND_  _1199_ (
    .A(_0394_),
    .B(_0387_),
    .Y(_0395_)
  );
  \$_AND_  _1200_ (
    .A(_0395_),
    .B(_0385_),
    .Y(_0396_)
  );
  \$_XOR_  _1201_ (
    .A(_0396_),
    .B(_0383_),
    .Y(_0397_)
  );
  \$_XOR_  _1202_ (
    .A(_0395_),
    .B(_0385_),
    .Y(_0398_)
  );
  \$_XOR_  _1203_ (
    .A(_0394_),
    .B(_0387_),
    .Y(_0399_)
  );
  \$_XOR_  _1204_ (
    .A(_0393_),
    .B(_0388_),
    .Y(_0400_)
  );
  \$_INV_  _1205_ (
    .A(_0400_),
    .Y(_0401_)
  );
  \$_OR_  _1206_ (
    .A(_0401_),
    .B(_0399_),
    .Y(_0402_)
  );
  \$_AND_  _1207_ (
    .A(_0402_),
    .B(_0398_),
    .Y(_0403_)
  );
  \$_XOR_  _1208_ (
    .A(_0403_),
    .B(_0397_),
    .Y(_0404_)
  );
  \$_AND_  _1209_ (
    .A(_0404_),
    .B(_0367_),
    .Y(_0405_)
  );
  \$_AND_  _1210_ (
    .A(_0405_),
    .B(_0365_),
    .Y(_0406_)
  );
  \$_AND_  _1211_ (
    .A(_0406_),
    .B(_0363_),
    .Y(_0407_)
  );
  \$_XOR_  _1212_ (
    .A(_0407_),
    .B(_0361_),
    .Y(_0408_)
  );
  \$_INV_  _1213_ (
    .A(_0408_),
    .Y(_0409_)
  );
  \$_AND_  _1214_ (
    .A(_0192_),
    .B(_0190_),
    .Y(_0410_)
  );
  \$_INV_  _1215_ (
    .A(_0349_),
    .Y(_0411_)
  );
  \$_AND_  _1216_ (
    .A(_0360_),
    .B(_0411_),
    .Y(_0412_)
  );
  \$_OR_  _1217_ (
    .A(_0412_),
    .B(_0410_),
    .Y(_0413_)
  );
  \$_INV_  _1218_ (
    .A(_0413_),
    .Y(_0414_)
  );
  \$_INV_  _1219_ (
    .A(_0361_),
    .Y(_0415_)
  );
  \$_AND_  _1220_ (
    .A(_0407_),
    .B(_0415_),
    .Y(_0416_)
  );
  \$_XOR_  _1221_ (
    .A(_0416_),
    .B(_0414_),
    .Y(_0417_)
  );
  \$_XOR_  _1222_ (
    .A(_0406_),
    .B(_0362_),
    .Y(_0418_)
  );
  \$_XOR_  _1223_ (
    .A(_0405_),
    .B(_0364_),
    .Y(_0419_)
  );
  \$_AND_  _1224_ (
    .A(_0419_),
    .B(_0418_),
    .Y(_0420_)
  );
  \$_OR_  _1225_ (
    .A(_0420_),
    .B(_0408_),
    .Y(_0421_)
  );
  \$_AND_  _1226_ (
    .A(_0421_),
    .B(_0417_),
    .Y(_0422_)
  );
  \$_XOR_  _1227_ (
    .A(_0420_),
    .B(_0408_),
    .Y(_0423_)
  );
  \$_MUX_  _1228_ (
    .A(_0423_),
    .B(_0409_),
    .S(_0422_),
    .Y(_0424_)
  );
  \$_AND_  _1229_ (
    .A(_0411_),
    .B(inst_alu[6]),
    .Y(_0425_)
  );
  \$_INV_  _1230_ (
    .A(_0425_),
    .Y(_0426_)
  );
  \$_AND_  _1231_ (
    .A(_0327_),
    .B(_0190_),
    .Y(_0427_)
  );
  \$_INV_  _1232_ (
    .A(_0427_),
    .Y(_0428_)
  );
  \$_OR_  _1233_ (
    .A(_0310_),
    .B(_0307_),
    .Y(_0429_)
  );
  \$_AND_  _1234_ (
    .A(inst_so[1]),
    .B(op_src[7]),
    .Y(_0430_)
  );
  \$_OR_  _1235_ (
    .A(_0430_),
    .B(_0330_),
    .Y(_0431_)
  );
  \$_INV_  _1236_ (
    .A(_0431_),
    .Y(_0432_)
  );
  \$_AND_  _1237_ (
    .A(_0432_),
    .B(_0429_),
    .Y(_0433_)
  );
  \$_AND_  _1238_ (
    .A(_0433_),
    .B(_0428_),
    .Y(_0434_)
  );
  \$_AND_  _1239_ (
    .A(_0410_),
    .B(inst_alu[4]),
    .Y(_0435_)
  );
  \$_INV_  _1240_ (
    .A(_0435_),
    .Y(_0436_)
  );
  \$_AND_  _1241_ (
    .A(_0193_),
    .B(_0189_),
    .Y(_0437_)
  );
  \$_OR_  _1242_ (
    .A(_0437_),
    .B(_0315_),
    .Y(_0438_)
  );
  \$_AND_  _1243_ (
    .A(_0438_),
    .B(_0436_),
    .Y(_0439_)
  );
  \$_AND_  _1244_ (
    .A(_0439_),
    .B(_0434_),
    .Y(_0440_)
  );
  \$_AND_  _1245_ (
    .A(_0440_),
    .B(_0426_),
    .Y(_0441_)
  );
  \$_INV_  _1246_ (
    .A(_0441_),
    .Y(_0442_)
  );
  \$_MUX_  _1247_ (
    .A(_0442_),
    .B(_0424_),
    .S(inst_alu[7]),
    .Y(_0443_)
  );
  \$_MUX_  _1248_ (
    .A(_0443_),
    .B(_0348_),
    .S(_0218_),
    .Y(alu_out[15])
  );
  \$_XOR_  _1249_ (
    .A(_0225_),
    .B(_0206_),
    .Y(_0444_)
  );
  \$_XOR_  _1250_ (
    .A(_0284_),
    .B(_0249_),
    .Y(_0445_)
  );
  \$_AND_  _1251_ (
    .A(_0249_),
    .B(inst_alu[6]),
    .Y(_0446_)
  );
  \$_INV_  _1252_ (
    .A(_0446_),
    .Y(_0447_)
  );
  \$_AND_  _1253_ (
    .A(_0089_),
    .B(_0094_),
    .Y(_0448_)
  );
  \$_OR_  _1254_ (
    .A(_0448_),
    .B(_0315_),
    .Y(_0449_)
  );
  \$_AND_  _1255_ (
    .A(_0237_),
    .B(inst_alu[4]),
    .Y(_0450_)
  );
  \$_AND_  _1256_ (
    .A(_0327_),
    .B(_0090_),
    .Y(_0451_)
  );
  \$_AND_  _1257_ (
    .A(inst_so[3]),
    .B(op_src[4]),
    .Y(_0452_)
  );
  \$_AND_  _1258_ (
    .A(op_src[5]),
    .B(inst_alu[10]),
    .Y(_0453_)
  );
  \$_AND_  _1259_ (
    .A(inst_so[1]),
    .B(op_src[12]),
    .Y(_0454_)
  );
  \$_OR_  _1260_ (
    .A(_0454_),
    .B(_0453_),
    .Y(_0455_)
  );
  \$_OR_  _1261_ (
    .A(_0455_),
    .B(_0452_),
    .Y(_0456_)
  );
  \$_OR_  _1262_ (
    .A(_0456_),
    .B(_0451_),
    .Y(_0457_)
  );
  \$_OR_  _1263_ (
    .A(_0457_),
    .B(_0450_),
    .Y(_0458_)
  );
  \$_INV_  _1264_ (
    .A(_0458_),
    .Y(_0459_)
  );
  \$_AND_  _1265_ (
    .A(_0459_),
    .B(_0449_),
    .Y(_0460_)
  );
  \$_AND_  _1266_ (
    .A(_0460_),
    .B(_0447_),
    .Y(_0461_)
  );
  \$_MUX_  _1267_ (
    .A(_0461_),
    .B(_0445_),
    .S(inst_alu[7]),
    .Y(_0462_)
  );
  \$_MUX_  _1268_ (
    .A(_0462_),
    .B(_0444_),
    .S(_0218_),
    .Y(_0463_)
  );
  \$_XOR_  _1269_ (
    .A(_0224_),
    .B(_0204_),
    .Y(_0464_)
  );
  \$_INV_  _1270_ (
    .A(_0278_),
    .Y(_0465_)
  );
  \$_AND_  _1271_ (
    .A(_0283_),
    .B(_0465_),
    .Y(_0466_)
  );
  \$_INV_  _1272_ (
    .A(_0282_),
    .Y(_0467_)
  );
  \$_XOR_  _1273_ (
    .A(_0467_),
    .B(_0279_),
    .Y(_0468_)
  );
  \$_MUX_  _1274_ (
    .A(_0468_),
    .B(_0279_),
    .S(_0466_),
    .Y(_0469_)
  );
  \$_AND_  _1275_ (
    .A(_0252_),
    .B(inst_alu[6]),
    .Y(_0470_)
  );
  \$_INV_  _1276_ (
    .A(_0470_),
    .Y(_0471_)
  );
  \$_AND_  _1277_ (
    .A(_0097_),
    .B(_0102_),
    .Y(_0472_)
  );
  \$_OR_  _1278_ (
    .A(_0472_),
    .B(_0315_),
    .Y(_0473_)
  );
  \$_AND_  _1279_ (
    .A(_0250_),
    .B(inst_alu[4]),
    .Y(_0474_)
  );
  \$_AND_  _1280_ (
    .A(_0327_),
    .B(_0098_),
    .Y(_0475_)
  );
  \$_AND_  _1281_ (
    .A(inst_so[3]),
    .B(op_src[3]),
    .Y(_0476_)
  );
  \$_AND_  _1282_ (
    .A(op_src[4]),
    .B(inst_alu[10]),
    .Y(_0477_)
  );
  \$_AND_  _1283_ (
    .A(inst_so[1]),
    .B(op_src[11]),
    .Y(_0478_)
  );
  \$_OR_  _1284_ (
    .A(_0478_),
    .B(_0477_),
    .Y(_0479_)
  );
  \$_OR_  _1285_ (
    .A(_0479_),
    .B(_0476_),
    .Y(_0480_)
  );
  \$_OR_  _1286_ (
    .A(_0480_),
    .B(_0475_),
    .Y(_0481_)
  );
  \$_OR_  _1287_ (
    .A(_0481_),
    .B(_0474_),
    .Y(_0482_)
  );
  \$_INV_  _1288_ (
    .A(_0482_),
    .Y(_0483_)
  );
  \$_AND_  _1289_ (
    .A(_0483_),
    .B(_0473_),
    .Y(_0484_)
  );
  \$_AND_  _1290_ (
    .A(_0484_),
    .B(_0471_),
    .Y(_0485_)
  );
  \$_MUX_  _1291_ (
    .A(_0485_),
    .B(_0469_),
    .S(inst_alu[7]),
    .Y(_0486_)
  );
  \$_MUX_  _1292_ (
    .A(_0486_),
    .B(_0464_),
    .S(_0218_),
    .Y(_0487_)
  );
  \$_XOR_  _1293_ (
    .A(_0221_),
    .B(_0017_),
    .Y(_0488_)
  );
  \$_XOR_  _1294_ (
    .A(_0272_),
    .B(status[0]),
    .Y(_0489_)
  );
  \$_AND_  _1295_ (
    .A(_0273_),
    .B(inst_alu[6]),
    .Y(_0490_)
  );
  \$_INV_  _1296_ (
    .A(_0490_),
    .Y(_0491_)
  );
  \$_AND_  _1297_ (
    .A(_0000_),
    .B(_0118_),
    .Y(_0492_)
  );
  \$_OR_  _1298_ (
    .A(_0492_),
    .B(_0315_),
    .Y(_0493_)
  );
  \$_AND_  _1299_ (
    .A(_0259_),
    .B(inst_alu[4]),
    .Y(_0494_)
  );
  \$_AND_  _1300_ (
    .A(_0327_),
    .B(_0784_),
    .Y(_0495_)
  );
  \$_AND_  _1301_ (
    .A(inst_so[3]),
    .B(op_src[0]),
    .Y(_0496_)
  );
  \$_AND_  _1302_ (
    .A(inst_alu[10]),
    .B(op_src[1]),
    .Y(_0497_)
  );
  \$_AND_  _1303_ (
    .A(inst_so[1]),
    .B(op_src[8]),
    .Y(_0498_)
  );
  \$_OR_  _1304_ (
    .A(_0498_),
    .B(_0497_),
    .Y(_0499_)
  );
  \$_OR_  _1305_ (
    .A(_0499_),
    .B(_0496_),
    .Y(_0500_)
  );
  \$_OR_  _1306_ (
    .A(_0500_),
    .B(_0495_),
    .Y(_0501_)
  );
  \$_OR_  _1307_ (
    .A(_0501_),
    .B(_0494_),
    .Y(_0502_)
  );
  \$_INV_  _1308_ (
    .A(_0502_),
    .Y(_0503_)
  );
  \$_AND_  _1309_ (
    .A(_0503_),
    .B(_0493_),
    .Y(_0504_)
  );
  \$_AND_  _1310_ (
    .A(_0504_),
    .B(_0491_),
    .Y(_0505_)
  );
  \$_MUX_  _1311_ (
    .A(_0505_),
    .B(_0489_),
    .S(inst_alu[7]),
    .Y(_0506_)
  );
  \$_MUX_  _1312_ (
    .A(_0506_),
    .B(_0488_),
    .S(_0218_),
    .Y(_0507_)
  );
  \$_AND_  _1313_ (
    .A(_0507_),
    .B(_0487_),
    .Y(_0508_)
  );
  \$_XOR_  _1314_ (
    .A(_0223_),
    .B(_0202_),
    .Y(_0509_)
  );
  \$_XOR_  _1315_ (
    .A(_0281_),
    .B(_0280_),
    .Y(_0510_)
  );
  \$_MUX_  _1316_ (
    .A(_0510_),
    .B(_0280_),
    .S(_0466_),
    .Y(_0511_)
  );
  \$_AND_  _1317_ (
    .A(_0255_),
    .B(inst_alu[6]),
    .Y(_0512_)
  );
  \$_INV_  _1318_ (
    .A(_0512_),
    .Y(_0513_)
  );
  \$_AND_  _1319_ (
    .A(_0106_),
    .B(_0104_),
    .Y(_0514_)
  );
  \$_OR_  _1320_ (
    .A(_0514_),
    .B(_0315_),
    .Y(_0515_)
  );
  \$_AND_  _1321_ (
    .A(_0253_),
    .B(inst_alu[4]),
    .Y(_0516_)
  );
  \$_AND_  _1322_ (
    .A(_0327_),
    .B(_0107_),
    .Y(_0517_)
  );
  \$_AND_  _1323_ (
    .A(inst_so[3]),
    .B(op_src[2]),
    .Y(_0518_)
  );
  \$_AND_  _1324_ (
    .A(op_src[3]),
    .B(inst_alu[10]),
    .Y(_0519_)
  );
  \$_AND_  _1325_ (
    .A(inst_so[1]),
    .B(op_src[10]),
    .Y(_0520_)
  );
  \$_OR_  _1326_ (
    .A(_0520_),
    .B(_0519_),
    .Y(_0521_)
  );
  \$_OR_  _1327_ (
    .A(_0521_),
    .B(_0518_),
    .Y(_0522_)
  );
  \$_OR_  _1328_ (
    .A(_0522_),
    .B(_0517_),
    .Y(_0523_)
  );
  \$_OR_  _1329_ (
    .A(_0523_),
    .B(_0516_),
    .Y(_0524_)
  );
  \$_INV_  _1330_ (
    .A(_0524_),
    .Y(_0525_)
  );
  \$_AND_  _1331_ (
    .A(_0525_),
    .B(_0515_),
    .Y(_0526_)
  );
  \$_AND_  _1332_ (
    .A(_0526_),
    .B(_0513_),
    .Y(_0527_)
  );
  \$_MUX_  _1333_ (
    .A(_0527_),
    .B(_0511_),
    .S(inst_alu[7]),
    .Y(_0528_)
  );
  \$_MUX_  _1334_ (
    .A(_0528_),
    .B(_0509_),
    .S(_0218_),
    .Y(_0529_)
  );
  \$_XOR_  _1335_ (
    .A(_0222_),
    .B(_0200_),
    .Y(_0530_)
  );
  \$_XOR_  _1336_ (
    .A(_0466_),
    .B(_0281_),
    .Y(_0531_)
  );
  \$_INV_  _1337_ (
    .A(_0531_),
    .Y(_0532_)
  );
  \$_AND_  _1338_ (
    .A(_0258_),
    .B(inst_alu[6]),
    .Y(_0533_)
  );
  \$_INV_  _1339_ (
    .A(_0533_),
    .Y(_0534_)
  );
  \$_AND_  _1340_ (
    .A(_0114_),
    .B(_0112_),
    .Y(_0535_)
  );
  \$_OR_  _1341_ (
    .A(_0535_),
    .B(_0315_),
    .Y(_0536_)
  );
  \$_AND_  _1342_ (
    .A(_0256_),
    .B(inst_alu[4]),
    .Y(_0537_)
  );
  \$_AND_  _1343_ (
    .A(_0327_),
    .B(_0113_),
    .Y(_0538_)
  );
  \$_AND_  _1344_ (
    .A(inst_so[3]),
    .B(op_src[1]),
    .Y(_0539_)
  );
  \$_AND_  _1345_ (
    .A(op_src[2]),
    .B(inst_alu[10]),
    .Y(_0540_)
  );
  \$_AND_  _1346_ (
    .A(inst_so[1]),
    .B(op_src[9]),
    .Y(_0541_)
  );
  \$_OR_  _1347_ (
    .A(_0541_),
    .B(_0540_),
    .Y(_0542_)
  );
  \$_OR_  _1348_ (
    .A(_0542_),
    .B(_0539_),
    .Y(_0543_)
  );
  \$_OR_  _1349_ (
    .A(_0543_),
    .B(_0538_),
    .Y(_0544_)
  );
  \$_OR_  _1350_ (
    .A(_0544_),
    .B(_0537_),
    .Y(_0545_)
  );
  \$_INV_  _1351_ (
    .A(_0545_),
    .Y(_0546_)
  );
  \$_AND_  _1352_ (
    .A(_0546_),
    .B(_0536_),
    .Y(_0547_)
  );
  \$_AND_  _1353_ (
    .A(_0547_),
    .B(_0534_),
    .Y(_0548_)
  );
  \$_MUX_  _1354_ (
    .A(_0548_),
    .B(_0532_),
    .S(inst_alu[7]),
    .Y(_0549_)
  );
  \$_MUX_  _1355_ (
    .A(_0549_),
    .B(_0530_),
    .S(_0218_),
    .Y(_0550_)
  );
  \$_AND_  _1356_ (
    .A(_0550_),
    .B(_0529_),
    .Y(_0551_)
  );
  \$_AND_  _1357_ (
    .A(_0551_),
    .B(_0508_),
    .Y(_0552_)
  );
  \$_AND_  _1358_ (
    .A(_0552_),
    .B(_0463_),
    .Y(_0553_)
  );
  \$_AND_  _1359_ (
    .A(_0553_),
    .B(_0339_),
    .Y(_0554_)
  );
  \$_XOR_  _1360_ (
    .A(_0227_),
    .B(_0210_),
    .Y(_0555_)
  );
  \$_INV_  _1361_ (
    .A(_0298_),
    .Y(_0556_)
  );
  \$_XOR_  _1362_ (
    .A(_0300_),
    .B(_0298_),
    .Y(_0557_)
  );
  \$_MUX_  _1363_ (
    .A(_0557_),
    .B(_0556_),
    .S(_0304_),
    .Y(_0558_)
  );
  \$_AND_  _1364_ (
    .A(_0233_),
    .B(inst_alu[6]),
    .Y(_0559_)
  );
  \$_INV_  _1365_ (
    .A(_0559_),
    .Y(_0560_)
  );
  \$_AND_  _1366_ (
    .A(_0073_),
    .B(_0078_),
    .Y(_0561_)
  );
  \$_OR_  _1367_ (
    .A(_0561_),
    .B(_0315_),
    .Y(_0562_)
  );
  \$_AND_  _1368_ (
    .A(_0231_),
    .B(inst_alu[4]),
    .Y(_0563_)
  );
  \$_AND_  _1369_ (
    .A(_0327_),
    .B(_0074_),
    .Y(_0564_)
  );
  \$_AND_  _1370_ (
    .A(inst_so[3]),
    .B(op_src[6]),
    .Y(_0565_)
  );
  \$_AND_  _1371_ (
    .A(op_src[7]),
    .B(inst_alu[10]),
    .Y(_0566_)
  );
  \$_AND_  _1372_ (
    .A(inst_so[1]),
    .B(op_src[14]),
    .Y(_0567_)
  );
  \$_OR_  _1373_ (
    .A(_0567_),
    .B(_0566_),
    .Y(_0568_)
  );
  \$_OR_  _1374_ (
    .A(_0568_),
    .B(_0565_),
    .Y(_0569_)
  );
  \$_OR_  _1375_ (
    .A(_0569_),
    .B(_0564_),
    .Y(_0570_)
  );
  \$_OR_  _1376_ (
    .A(_0570_),
    .B(_0563_),
    .Y(_0571_)
  );
  \$_INV_  _1377_ (
    .A(_0571_),
    .Y(_0572_)
  );
  \$_AND_  _1378_ (
    .A(_0572_),
    .B(_0562_),
    .Y(_0573_)
  );
  \$_AND_  _1379_ (
    .A(_0573_),
    .B(_0560_),
    .Y(_0574_)
  );
  \$_MUX_  _1380_ (
    .A(_0574_),
    .B(_0558_),
    .S(inst_alu[7]),
    .Y(_0575_)
  );
  \$_MUX_  _1381_ (
    .A(_0575_),
    .B(_0555_),
    .S(_0218_),
    .Y(_0576_)
  );
  \$_XOR_  _1382_ (
    .A(_0226_),
    .B(_0208_),
    .Y(_0577_)
  );
  \$_XOR_  _1383_ (
    .A(_0304_),
    .B(_0300_),
    .Y(_0578_)
  );
  \$_AND_  _1384_ (
    .A(_0236_),
    .B(inst_alu[6]),
    .Y(_0579_)
  );
  \$_INV_  _1385_ (
    .A(_0579_),
    .Y(_0580_)
  );
  \$_AND_  _1386_ (
    .A(_0081_),
    .B(_0086_),
    .Y(_0581_)
  );
  \$_OR_  _1387_ (
    .A(_0581_),
    .B(_0315_),
    .Y(_0582_)
  );
  \$_AND_  _1388_ (
    .A(_0234_),
    .B(inst_alu[4]),
    .Y(_0583_)
  );
  \$_AND_  _1389_ (
    .A(_0327_),
    .B(_0082_),
    .Y(_0584_)
  );
  \$_AND_  _1390_ (
    .A(inst_so[3]),
    .B(op_src[5]),
    .Y(_0585_)
  );
  \$_AND_  _1391_ (
    .A(op_src[6]),
    .B(inst_alu[10]),
    .Y(_0586_)
  );
  \$_AND_  _1392_ (
    .A(inst_so[1]),
    .B(op_src[13]),
    .Y(_0587_)
  );
  \$_OR_  _1393_ (
    .A(_0587_),
    .B(_0586_),
    .Y(_0588_)
  );
  \$_OR_  _1394_ (
    .A(_0588_),
    .B(_0585_),
    .Y(_0589_)
  );
  \$_OR_  _1395_ (
    .A(_0589_),
    .B(_0584_),
    .Y(_0590_)
  );
  \$_OR_  _1396_ (
    .A(_0590_),
    .B(_0583_),
    .Y(_0591_)
  );
  \$_INV_  _1397_ (
    .A(_0591_),
    .Y(_0592_)
  );
  \$_AND_  _1398_ (
    .A(_0592_),
    .B(_0582_),
    .Y(_0593_)
  );
  \$_AND_  _1399_ (
    .A(_0593_),
    .B(_0580_),
    .Y(_0594_)
  );
  \$_MUX_  _1400_ (
    .A(_0594_),
    .B(_0578_),
    .S(inst_alu[7]),
    .Y(_0595_)
  );
  \$_MUX_  _1401_ (
    .A(_0595_),
    .B(_0577_),
    .S(_0218_),
    .Y(_0596_)
  );
  \$_AND_  _1402_ (
    .A(_0596_),
    .B(_0576_),
    .Y(_0597_)
  );
  \$_AND_  _1403_ (
    .A(_0597_),
    .B(_0554_),
    .Y(_0598_)
  );
  \$_AND_  _1404_ (
    .A(_0598_),
    .B(inst_bw),
    .Y(_0599_)
  );
  \$_INV_  _1405_ (
    .A(_0599_),
    .Y(_0600_)
  );
  \$_XOR_  _1406_ (
    .A(_0344_),
    .B(alu_add[12]),
    .Y(_0601_)
  );
  \$_XOR_  _1407_ (
    .A(_0404_),
    .B(_0366_),
    .Y(_0602_)
  );
  \$_AND_  _1408_ (
    .A(_0367_),
    .B(inst_alu[6]),
    .Y(_0603_)
  );
  \$_INV_  _1409_ (
    .A(_0603_),
    .Y(_0604_)
  );
  \$_AND_  _1410_ (
    .A(_0157_),
    .B(_0153_),
    .Y(_0605_)
  );
  \$_OR_  _1411_ (
    .A(_0605_),
    .B(_0315_),
    .Y(_0606_)
  );
  \$_AND_  _1412_ (
    .A(_0356_),
    .B(inst_alu[4]),
    .Y(_0607_)
  );
  \$_AND_  _1413_ (
    .A(_0327_),
    .B(_0154_),
    .Y(_0608_)
  );
  \$_AND_  _1414_ (
    .A(inst_so[1]),
    .B(op_src[4]),
    .Y(_0609_)
  );
  \$_AND_  _1415_ (
    .A(op_src[13]),
    .B(inst_alu[10]),
    .Y(_0610_)
  );
  \$_OR_  _1416_ (
    .A(_0610_),
    .B(_0330_),
    .Y(_0611_)
  );
  \$_OR_  _1417_ (
    .A(_0611_),
    .B(_0609_),
    .Y(_0612_)
  );
  \$_OR_  _1418_ (
    .A(_0612_),
    .B(_0608_),
    .Y(_0613_)
  );
  \$_OR_  _1419_ (
    .A(_0613_),
    .B(_0607_),
    .Y(_0614_)
  );
  \$_INV_  _1420_ (
    .A(_0614_),
    .Y(_0615_)
  );
  \$_AND_  _1421_ (
    .A(_0615_),
    .B(_0606_),
    .Y(_0616_)
  );
  \$_AND_  _1422_ (
    .A(_0616_),
    .B(_0604_),
    .Y(_0617_)
  );
  \$_MUX_  _1423_ (
    .A(_0617_),
    .B(_0602_),
    .S(inst_alu[7]),
    .Y(_0618_)
  );
  \$_INV_  _1424_ (
    .A(_0618_),
    .Y(_0619_)
  );
  \$_MUX_  _1425_ (
    .A(_0619_),
    .B(_0601_),
    .S(_0218_),
    .Y(alu_out[12])
  );
  \$_XOR_  _1426_ (
    .A(_0343_),
    .B(alu_add[11]),
    .Y(_0620_)
  );
  \$_INV_  _1427_ (
    .A(_0398_),
    .Y(_0621_)
  );
  \$_INV_  _1428_ (
    .A(_0397_),
    .Y(_0622_)
  );
  \$_INV_  _1429_ (
    .A(_0403_),
    .Y(_0623_)
  );
  \$_AND_  _1430_ (
    .A(_0623_),
    .B(_0622_),
    .Y(_0624_)
  );
  \$_XOR_  _1431_ (
    .A(_0402_),
    .B(_0621_),
    .Y(_0625_)
  );
  \$_MUX_  _1432_ (
    .A(_0625_),
    .B(_0621_),
    .S(_0624_),
    .Y(_0626_)
  );
  \$_AND_  _1433_ (
    .A(_0370_),
    .B(inst_alu[6]),
    .Y(_0627_)
  );
  \$_INV_  _1434_ (
    .A(_0627_),
    .Y(_0628_)
  );
  \$_AND_  _1435_ (
    .A(_0145_),
    .B(_0141_),
    .Y(_0629_)
  );
  \$_OR_  _1436_ (
    .A(_0629_),
    .B(_0315_),
    .Y(_0630_)
  );
  \$_AND_  _1437_ (
    .A(_0368_),
    .B(inst_alu[4]),
    .Y(_0631_)
  );
  \$_AND_  _1438_ (
    .A(_0327_),
    .B(_0142_),
    .Y(_0632_)
  );
  \$_AND_  _1439_ (
    .A(inst_so[1]),
    .B(op_src[3]),
    .Y(_0633_)
  );
  \$_AND_  _1440_ (
    .A(op_src[12]),
    .B(inst_alu[10]),
    .Y(_0634_)
  );
  \$_OR_  _1441_ (
    .A(_0634_),
    .B(_0330_),
    .Y(_0635_)
  );
  \$_OR_  _1442_ (
    .A(_0635_),
    .B(_0633_),
    .Y(_0636_)
  );
  \$_OR_  _1443_ (
    .A(_0636_),
    .B(_0632_),
    .Y(_0637_)
  );
  \$_OR_  _1444_ (
    .A(_0637_),
    .B(_0631_),
    .Y(_0638_)
  );
  \$_INV_  _1445_ (
    .A(_0638_),
    .Y(_0639_)
  );
  \$_AND_  _1446_ (
    .A(_0639_),
    .B(_0630_),
    .Y(_0640_)
  );
  \$_AND_  _1447_ (
    .A(_0640_),
    .B(_0628_),
    .Y(_0641_)
  );
  \$_MUX_  _1448_ (
    .A(_0641_),
    .B(_0626_),
    .S(inst_alu[7]),
    .Y(_0642_)
  );
  \$_INV_  _1449_ (
    .A(_0642_),
    .Y(_0643_)
  );
  \$_MUX_  _1450_ (
    .A(_0643_),
    .B(_0620_),
    .S(_0218_),
    .Y(alu_out[11])
  );
  \$_XOR_  _1451_ (
    .A(_0340_),
    .B(_0214_),
    .Y(_0644_)
  );
  \$_XOR_  _1452_ (
    .A(_0392_),
    .B(_0390_),
    .Y(_0645_)
  );
  \$_AND_  _1453_ (
    .A(_0391_),
    .B(inst_alu[6]),
    .Y(_0646_)
  );
  \$_INV_  _1454_ (
    .A(_0646_),
    .Y(_0647_)
  );
  \$_AND_  _1455_ (
    .A(_0062_),
    .B(_0056_),
    .Y(_0648_)
  );
  \$_OR_  _1456_ (
    .A(_0648_),
    .B(_0315_),
    .Y(_0649_)
  );
  \$_AND_  _1457_ (
    .A(_0377_),
    .B(inst_alu[4]),
    .Y(_0650_)
  );
  \$_AND_  _1458_ (
    .A(_0327_),
    .B(_0057_),
    .Y(_0651_)
  );
  \$_AND_  _1459_ (
    .A(op_src[0]),
    .B(inst_so[1]),
    .Y(_0652_)
  );
  \$_AND_  _1460_ (
    .A(op_src[9]),
    .B(inst_alu[10]),
    .Y(_0653_)
  );
  \$_OR_  _1461_ (
    .A(_0653_),
    .B(_0330_),
    .Y(_0654_)
  );
  \$_OR_  _1462_ (
    .A(_0654_),
    .B(_0652_),
    .Y(_0655_)
  );
  \$_OR_  _1463_ (
    .A(_0655_),
    .B(_0651_),
    .Y(_0656_)
  );
  \$_OR_  _1464_ (
    .A(_0656_),
    .B(_0650_),
    .Y(_0657_)
  );
  \$_INV_  _1465_ (
    .A(_0657_),
    .Y(_0658_)
  );
  \$_AND_  _1466_ (
    .A(_0658_),
    .B(_0649_),
    .Y(_0659_)
  );
  \$_AND_  _1467_ (
    .A(_0659_),
    .B(_0647_),
    .Y(_0660_)
  );
  \$_MUX_  _1468_ (
    .A(_0660_),
    .B(_0645_),
    .S(inst_alu[7]),
    .Y(_0661_)
  );
  \$_MUX_  _1469_ (
    .A(_0661_),
    .B(_0644_),
    .S(_0218_),
    .Y(_0662_)
  );
  \$_AND_  _1470_ (
    .A(_0598_),
    .B(_0308_),
    .Y(_0663_)
  );
  \$_AND_  _1471_ (
    .A(_0663_),
    .B(_0662_),
    .Y(_0664_)
  );
  \$_INV_  _1472_ (
    .A(_0664_),
    .Y(_0665_)
  );
  \$_OR_  _1473_ (
    .A(_0665_),
    .B(alu_out[11]),
    .Y(_0666_)
  );
  \$_XOR_  _1474_ (
    .A(_0342_),
    .B(_0138_),
    .Y(_0667_)
  );
  \$_INV_  _1475_ (
    .A(_0399_),
    .Y(_0668_)
  );
  \$_XOR_  _1476_ (
    .A(_0401_),
    .B(_0399_),
    .Y(_0669_)
  );
  \$_MUX_  _1477_ (
    .A(_0669_),
    .B(_0668_),
    .S(_0624_),
    .Y(_0670_)
  );
  \$_AND_  _1478_ (
    .A(_0373_),
    .B(inst_alu[6]),
    .Y(_0671_)
  );
  \$_INV_  _1479_ (
    .A(_0671_),
    .Y(_0672_)
  );
  \$_AND_  _1480_ (
    .A(_0041_),
    .B(_0036_),
    .Y(_0673_)
  );
  \$_OR_  _1481_ (
    .A(_0673_),
    .B(_0315_),
    .Y(_0674_)
  );
  \$_AND_  _1482_ (
    .A(_0371_),
    .B(inst_alu[4]),
    .Y(_0675_)
  );
  \$_AND_  _1483_ (
    .A(_0327_),
    .B(_0037_),
    .Y(_0676_)
  );
  \$_AND_  _1484_ (
    .A(inst_so[1]),
    .B(op_src[2]),
    .Y(_0677_)
  );
  \$_AND_  _1485_ (
    .A(op_src[11]),
    .B(inst_alu[10]),
    .Y(_0678_)
  );
  \$_OR_  _1486_ (
    .A(_0678_),
    .B(_0330_),
    .Y(_0679_)
  );
  \$_OR_  _1487_ (
    .A(_0679_),
    .B(_0677_),
    .Y(_0680_)
  );
  \$_OR_  _1488_ (
    .A(_0680_),
    .B(_0676_),
    .Y(_0681_)
  );
  \$_OR_  _1489_ (
    .A(_0681_),
    .B(_0675_),
    .Y(_0682_)
  );
  \$_INV_  _1490_ (
    .A(_0682_),
    .Y(_0683_)
  );
  \$_AND_  _1491_ (
    .A(_0683_),
    .B(_0674_),
    .Y(_0684_)
  );
  \$_AND_  _1492_ (
    .A(_0684_),
    .B(_0672_),
    .Y(_0685_)
  );
  \$_MUX_  _1493_ (
    .A(_0685_),
    .B(_0670_),
    .S(inst_alu[7]),
    .Y(_0686_)
  );
  \$_MUX_  _1494_ (
    .A(_0686_),
    .B(_0667_),
    .S(_0218_),
    .Y(_0687_)
  );
  \$_XOR_  _1495_ (
    .A(_0341_),
    .B(_0216_),
    .Y(_0688_)
  );
  \$_XOR_  _1496_ (
    .A(_0624_),
    .B(_0401_),
    .Y(_0689_)
  );
  \$_AND_  _1497_ (
    .A(_0376_),
    .B(inst_alu[6]),
    .Y(_0690_)
  );
  \$_INV_  _1498_ (
    .A(_0690_),
    .Y(_0691_)
  );
  \$_AND_  _1499_ (
    .A(_0052_),
    .B(_0046_),
    .Y(_0692_)
  );
  \$_OR_  _1500_ (
    .A(_0692_),
    .B(_0315_),
    .Y(_0693_)
  );
  \$_AND_  _1501_ (
    .A(_0374_),
    .B(inst_alu[4]),
    .Y(_0694_)
  );
  \$_AND_  _1502_ (
    .A(_0327_),
    .B(_0047_),
    .Y(_0695_)
  );
  \$_AND_  _1503_ (
    .A(inst_so[1]),
    .B(op_src[1]),
    .Y(_0696_)
  );
  \$_AND_  _1504_ (
    .A(op_src[10]),
    .B(inst_alu[10]),
    .Y(_0697_)
  );
  \$_OR_  _1505_ (
    .A(_0697_),
    .B(_0330_),
    .Y(_0698_)
  );
  \$_OR_  _1506_ (
    .A(_0698_),
    .B(_0696_),
    .Y(_0699_)
  );
  \$_OR_  _1507_ (
    .A(_0699_),
    .B(_0695_),
    .Y(_0700_)
  );
  \$_OR_  _1508_ (
    .A(_0700_),
    .B(_0694_),
    .Y(_0701_)
  );
  \$_INV_  _1509_ (
    .A(_0701_),
    .Y(_0702_)
  );
  \$_AND_  _1510_ (
    .A(_0702_),
    .B(_0693_),
    .Y(_0703_)
  );
  \$_AND_  _1511_ (
    .A(_0703_),
    .B(_0691_),
    .Y(_0704_)
  );
  \$_MUX_  _1512_ (
    .A(_0704_),
    .B(_0689_),
    .S(inst_alu[7]),
    .Y(_0705_)
  );
  \$_MUX_  _1513_ (
    .A(_0705_),
    .B(_0688_),
    .S(_0218_),
    .Y(_0706_)
  );
  \$_AND_  _1514_ (
    .A(_0706_),
    .B(_0687_),
    .Y(_0707_)
  );
  \$_INV_  _1515_ (
    .A(_0707_),
    .Y(_0708_)
  );
  \$_OR_  _1516_ (
    .A(_0708_),
    .B(_0666_),
    .Y(_0709_)
  );
  \$_OR_  _1517_ (
    .A(_0709_),
    .B(alu_out[12]),
    .Y(_0710_)
  );
  \$_OR_  _1518_ (
    .A(_0710_),
    .B(alu_out[15]),
    .Y(_0711_)
  );
  \$_XOR_  _1519_ (
    .A(_0346_),
    .B(alu_add[14]),
    .Y(_0712_)
  );
  \$_INV_  _1520_ (
    .A(_0418_),
    .Y(_0713_)
  );
  \$_XOR_  _1521_ (
    .A(_0419_),
    .B(_0418_),
    .Y(_0714_)
  );
  \$_INV_  _1522_ (
    .A(_0714_),
    .Y(_0715_)
  );
  \$_MUX_  _1523_ (
    .A(_0715_),
    .B(_0713_),
    .S(_0422_),
    .Y(_0716_)
  );
  \$_AND_  _1524_ (
    .A(_0352_),
    .B(inst_alu[6]),
    .Y(_0717_)
  );
  \$_INV_  _1525_ (
    .A(_0717_),
    .Y(_0718_)
  );
  \$_AND_  _1526_ (
    .A(_0181_),
    .B(_0177_),
    .Y(_0719_)
  );
  \$_OR_  _1527_ (
    .A(_0719_),
    .B(_0315_),
    .Y(_0720_)
  );
  \$_AND_  _1528_ (
    .A(_0350_),
    .B(inst_alu[4]),
    .Y(_0721_)
  );
  \$_AND_  _1529_ (
    .A(_0327_),
    .B(_0178_),
    .Y(_0722_)
  );
  \$_AND_  _1530_ (
    .A(inst_so[1]),
    .B(op_src[6]),
    .Y(_0723_)
  );
  \$_AND_  _1531_ (
    .A(op_src[15]),
    .B(inst_alu[10]),
    .Y(_0724_)
  );
  \$_OR_  _1532_ (
    .A(_0724_),
    .B(_0330_),
    .Y(_0725_)
  );
  \$_OR_  _1533_ (
    .A(_0725_),
    .B(_0723_),
    .Y(_0726_)
  );
  \$_OR_  _1534_ (
    .A(_0726_),
    .B(_0722_),
    .Y(_0727_)
  );
  \$_OR_  _1535_ (
    .A(_0727_),
    .B(_0721_),
    .Y(_0728_)
  );
  \$_INV_  _1536_ (
    .A(_0728_),
    .Y(_0729_)
  );
  \$_AND_  _1537_ (
    .A(_0729_),
    .B(_0720_),
    .Y(_0730_)
  );
  \$_AND_  _1538_ (
    .A(_0730_),
    .B(_0718_),
    .Y(_0731_)
  );
  \$_INV_  _1539_ (
    .A(_0731_),
    .Y(_0732_)
  );
  \$_MUX_  _1540_ (
    .A(_0732_),
    .B(_0716_),
    .S(inst_alu[7]),
    .Y(_0733_)
  );
  \$_MUX_  _1541_ (
    .A(_0733_),
    .B(_0712_),
    .S(_0218_),
    .Y(alu_out[14])
  );
  \$_XOR_  _1542_ (
    .A(_0345_),
    .B(alu_add[13]),
    .Y(_0734_)
  );
  \$_XOR_  _1543_ (
    .A(_0422_),
    .B(_0419_),
    .Y(_0735_)
  );
  \$_AND_  _1544_ (
    .A(_0355_),
    .B(inst_alu[6]),
    .Y(_0736_)
  );
  \$_INV_  _1545_ (
    .A(_0736_),
    .Y(_0737_)
  );
  \$_AND_  _1546_ (
    .A(_0169_),
    .B(_0165_),
    .Y(_0738_)
  );
  \$_OR_  _1547_ (
    .A(_0738_),
    .B(_0315_),
    .Y(_0739_)
  );
  \$_AND_  _1548_ (
    .A(_0353_),
    .B(inst_alu[4]),
    .Y(_0740_)
  );
  \$_AND_  _1549_ (
    .A(_0327_),
    .B(_0166_),
    .Y(_0741_)
  );
  \$_AND_  _1550_ (
    .A(inst_so[1]),
    .B(op_src[5]),
    .Y(_0742_)
  );
  \$_AND_  _1551_ (
    .A(op_src[14]),
    .B(inst_alu[10]),
    .Y(_0743_)
  );
  \$_OR_  _1552_ (
    .A(_0743_),
    .B(_0330_),
    .Y(_0744_)
  );
  \$_OR_  _1553_ (
    .A(_0744_),
    .B(_0742_),
    .Y(_0745_)
  );
  \$_OR_  _1554_ (
    .A(_0745_),
    .B(_0741_),
    .Y(_0746_)
  );
  \$_OR_  _1555_ (
    .A(_0746_),
    .B(_0740_),
    .Y(_0747_)
  );
  \$_INV_  _1556_ (
    .A(_0747_),
    .Y(_0748_)
  );
  \$_AND_  _1557_ (
    .A(_0748_),
    .B(_0739_),
    .Y(_0749_)
  );
  \$_AND_  _1558_ (
    .A(_0749_),
    .B(_0737_),
    .Y(_0750_)
  );
  \$_INV_  _1559_ (
    .A(_0750_),
    .Y(_0751_)
  );
  \$_MUX_  _1560_ (
    .A(_0751_),
    .B(_0735_),
    .S(inst_alu[7]),
    .Y(_0752_)
  );
  \$_MUX_  _1561_ (
    .A(_0752_),
    .B(_0734_),
    .S(_0218_),
    .Y(alu_out[13])
  );
  \$_OR_  _1562_ (
    .A(alu_out[13]),
    .B(alu_out[14]),
    .Y(_0753_)
  );
  \$_OR_  _1563_ (
    .A(_0753_),
    .B(_0711_),
    .Y(_0754_)
  );
  \$_AND_  _1564_ (
    .A(_0754_),
    .B(_0600_),
    .Y(_0755_)
  );
  \$_INV_  _1565_ (
    .A(_0755_),
    .Y(Z)
  );
  \$_INV_  _1566_ (
    .A(_0507_),
    .Y(alu_out[0])
  );
  \$_INV_  _1567_ (
    .A(_0550_),
    .Y(alu_out[1])
  );
  \$_INV_  _1568_ (
    .A(_0529_),
    .Y(alu_out[2])
  );
  \$_INV_  _1569_ (
    .A(_0487_),
    .Y(alu_out[3])
  );
  \$_INV_  _1570_ (
    .A(_0463_),
    .Y(alu_out[4])
  );
  \$_INV_  _1571_ (
    .A(_0596_),
    .Y(alu_out[5])
  );
  \$_INV_  _1572_ (
    .A(_0576_),
    .Y(alu_out[6])
  );
  \$_INV_  _1573_ (
    .A(_0687_),
    .Y(alu_out[10])
  );
  \$_INV_  _1574_ (
    .A(_0662_),
    .Y(alu_out[8])
  );
  \$_INV_  _1575_ (
    .A(_0706_),
    .Y(alu_out[9])
  );
  \$_MUX_  _1576_ (
    .A(alu_out[15]),
    .B(alu_out[7]),
    .S(inst_bw),
    .Y(N)
  );
  \$_INV_  _1577_ (
    .A(_0191_),
    .Y(_0756_)
  );
  \$_OR_  _1578_ (
    .A(_0193_),
    .B(_0756_),
    .Y(_0757_)
  );
  \$_OR_  _1579_ (
    .A(_0198_),
    .B(_0194_),
    .Y(_0758_)
  );
  \$_AND_  _1580_ (
    .A(_0758_),
    .B(_0757_),
    .Y(_0759_)
  );
  \$_INV_  _1581_ (
    .A(_0194_),
    .Y(_0760_)
  );
  \$_XOR_  _1582_ (
    .A(_0198_),
    .B(_0760_),
    .Y(_0761_)
  );
  \$_INV_  _1583_ (
    .A(alu_add[14]),
    .Y(_0762_)
  );
  \$_INV_  _1584_ (
    .A(_0346_),
    .Y(_0763_)
  );
  \$_OR_  _1585_ (
    .A(_0763_),
    .B(_0762_),
    .Y(_0764_)
  );
  \$_OR_  _1586_ (
    .A(_0764_),
    .B(_0761_),
    .Y(_0765_)
  );
  \$_XOR_  _1587_ (
    .A(_0765_),
    .B(_0759_),
    .Y(_0766_)
  );
  \$_AND_  _1588_ (
    .A(_0766_),
    .B(_0218_),
    .Y(_0767_)
  );
  \$_XOR_  _1589_ (
    .A(_0421_),
    .B(_0417_),
    .Y(_0768_)
  );
  \$_INV_  _1590_ (
    .A(_0218_),
    .Y(_0769_)
  );
  \$_AND_  _1591_ (
    .A(_0769_),
    .B(inst_alu[7]),
    .Y(_0770_)
  );
  \$_AND_  _1592_ (
    .A(_0770_),
    .B(_0768_),
    .Y(_0771_)
  );
  \$_OR_  _1593_ (
    .A(_0771_),
    .B(_0767_),
    .Y(_0772_)
  );
  \$_MUX_  _1594_ (
    .A(_0772_),
    .B(alu_out[8]),
    .S(inst_bw),
    .Y(_0773_)
  );
  \$_MUX_  _1595_ (
    .A(_0773_),
    .B(_0755_),
    .S(inst_alu[6]),
    .Y(_0774_)
  );
  \$_MUX_  _1596_ (
    .A(_0774_),
    .B(_0755_),
    .S(inst_alu[8]),
    .Y(_0775_)
  );
  \$_MUX_  _1597_ (
    .A(_0775_),
    .B(_0784_),
    .S(inst_alu[10]),
    .Y(alu_stat[0])
  );
  \$_MUX_  _1598_ (
    .A(_0410_),
    .B(_0291_),
    .S(inst_bw),
    .Y(_0776_)
  );
  \$_MUX_  _1599_ (
    .A(_0316_),
    .B(_0291_),
    .S(_0339_),
    .Y(_0777_)
  );
  \$_MUX_  _1600_ (
    .A(_0410_),
    .B(_0437_),
    .S(alu_out[15]),
    .Y(_0778_)
  );
  \$_MUX_  _1601_ (
    .A(_0778_),
    .B(_0777_),
    .S(inst_bw),
    .Y(_0779_)
  );
  \$_MUX_  _1602_ (
    .A(_0779_),
    .B(_0776_),
    .S(inst_alu[6]),
    .Y(_0780_)
  );
  \$_INV_  _1603_ (
    .A(inst_alu[8]),
    .Y(_0781_)
  );
  \$_AND_  _1604_ (
    .A(_0781_),
    .B(_0307_),
    .Y(_0782_)
  );
  \$_AND_  _1605_ (
    .A(_0782_),
    .B(_0780_),
    .Y(alu_stat[3])
  );
  \$_AND_  _1606_ (
    .A(inst_alu[9]),
    .B(exec_cycle),
    .Y(alu_stat_wr[3])
  );
  assign alu_out_add = alu_add[15:0];
  assign alu_out_nxt[15:0] = alu_out;
  assign { alu_shift[16], alu_shift[14:8], alu_shift[6:0] } = { 1'b0, op_src[15:9], op_src[7:1] };
  assign alu_stat[2:1] = { N, Z };
  assign alu_stat_wr[2:0] = { alu_stat_wr[3], alu_stat_wr[3], alu_stat_wr[3] };
  assign alu_swpb = { 1'b0, op_src[7:0], op_src[15:8] };
  assign alu_sxt = { 1'b0, op_src[7], op_src[7], op_src[7], op_src[7], op_src[7], op_src[7], op_src[7], op_src[7], op_src[7:0] };
  assign { op_dst_in[16], op_dst_in[7:0] } = { 1'b0, op_dst[7:0] };
endmodule

module omsp_clock_module(aclk, aclk_en, cpu_en_s, dbg_clk, dbg_en_s, dbg_rst, dco_enable, dco_wkup, lfxt_enable, lfxt_wkup, mclk, per_dout, por, puc_pnd_set, puc_rst, smclk, smclk_en, cpu_en, cpuoff, dbg_cpu_reset, dbg_en, dco_clk, lfxt_clk, mclk_enable, mclk_wkup, oscoff, per_addr, per_din, per_en, per_we, reset_n, scan_enable, scan_mode, scg0, scg1, wdt_reset);
  wire [2:0] _000_;
  wire _001_;
  wire [7:0] _002_;
  wire [7:0] _003_;
  wire [2:0] _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  output aclk;
  wire [2:0] aclk_div;
  output aclk_en;
  wire [7:0] bcsctl1;
  wire [7:0] bcsctl1_nxt;
  wire [15:0] bcsctl1_rd;
  wire [7:0] bcsctl2;
  wire [7:0] bcsctl2_nxt;
  wire [15:0] bcsctl2_rd;
  input cpu_en;
  wire cpu_en_aux_s;
  output cpu_en_s;
  input cpuoff;
  output dbg_clk;
  input dbg_cpu_reset;
  input dbg_en;
  output dbg_en_s;
  output dbg_rst;
  wire dbg_rst_noscan;
  wire dbg_rst_nxt;
  input dco_clk;
  output dco_enable;
  output dco_wkup;
  input lfxt_clk;
  wire lfxt_clk_dly;
  wire lfxt_clk_s;
  output lfxt_enable;
  output lfxt_wkup;
  output mclk;
  input mclk_enable;
  input mclk_wkup;
  wire nodiv_mclk;
  wire nodiv_smclk;
  input oscoff;
  input [13:0] per_addr;
  input [15:0] per_din;
  output [15:0] per_dout;
  input per_en;
  input [1:0] per_we;
  output por;
  wire por_a;
  wire por_noscan;
  wire puc_a;
  wire puc_a_scan;
  wire puc_noscan_n;
  output puc_pnd_set;
  output puc_rst;
  wire [3:0] reg_addr;
  input reset_n;
  input scan_enable;
  input scan_mode;
  input scg0;
  input scg1;
  output smclk;
  wire [2:0] smclk_div;
  output smclk_en;
  input wdt_reset;
  \$_INV_  _109_ (
    .A(puc_noscan_n),
    .Y(puc_pnd_set)
  );
  \$_INV_  _110_ (
    .A(per_addr[2]),
    .Y(_006_)
  );
  \$_AND_  _111_ (
    .A(per_addr[0]),
    .B(_006_),
    .Y(_007_)
  );
  \$_AND_  _112_ (
    .A(_007_),
    .B(per_addr[1]),
    .Y(_008_)
  );
  \$_OR_  _113_ (
    .A(per_addr[12]),
    .B(per_addr[11]),
    .Y(_009_)
  );
  \$_INV_  _114_ (
    .A(_009_),
    .Y(_010_)
  );
  \$_AND_  _115_ (
    .A(per_addr[5]),
    .B(per_addr[3]),
    .Y(_011_)
  );
  \$_AND_  _116_ (
    .A(_011_),
    .B(_010_),
    .Y(_012_)
  );
  \$_INV_  _117_ (
    .A(per_addr[7]),
    .Y(_013_)
  );
  \$_INV_  _118_ (
    .A(per_addr[8]),
    .Y(_014_)
  );
  \$_AND_  _119_ (
    .A(_014_),
    .B(_013_),
    .Y(_015_)
  );
  \$_INV_  _120_ (
    .A(per_addr[9]),
    .Y(_016_)
  );
  \$_INV_  _121_ (
    .A(per_addr[10]),
    .Y(_017_)
  );
  \$_AND_  _122_ (
    .A(_017_),
    .B(_016_),
    .Y(_018_)
  );
  \$_AND_  _123_ (
    .A(_018_),
    .B(_015_),
    .Y(_019_)
  );
  \$_INV_  _124_ (
    .A(per_addr[13]),
    .Y(_020_)
  );
  \$_AND_  _125_ (
    .A(_020_),
    .B(per_en),
    .Y(_021_)
  );
  \$_INV_  _126_ (
    .A(per_addr[4]),
    .Y(_022_)
  );
  \$_INV_  _127_ (
    .A(per_addr[6]),
    .Y(_023_)
  );
  \$_AND_  _128_ (
    .A(_023_),
    .B(_022_),
    .Y(_024_)
  );
  \$_AND_  _129_ (
    .A(_024_),
    .B(_021_),
    .Y(_025_)
  );
  \$_AND_  _130_ (
    .A(_025_),
    .B(_019_),
    .Y(_026_)
  );
  \$_AND_  _131_ (
    .A(_026_),
    .B(_012_),
    .Y(_027_)
  );
  \$_INV_  _132_ (
    .A(per_we[0]),
    .Y(_028_)
  );
  \$_INV_  _133_ (
    .A(per_we[1]),
    .Y(_029_)
  );
  \$_AND_  _134_ (
    .A(_029_),
    .B(_028_),
    .Y(_030_)
  );
  \$_AND_  _135_ (
    .A(_030_),
    .B(_027_),
    .Y(_031_)
  );
  \$_AND_  _136_ (
    .A(_031_),
    .B(_008_),
    .Y(_032_)
  );
  \$_AND_  _137_ (
    .A(_032_),
    .B(bcsctl1[0]),
    .Y(bcsctl1_rd[8])
  );
  \$_AND_  _138_ (
    .A(_032_),
    .B(bcsctl1[1]),
    .Y(bcsctl1_rd[9])
  );
  \$_AND_  _139_ (
    .A(_032_),
    .B(bcsctl1[2]),
    .Y(bcsctl1_rd[10])
  );
  \$_AND_  _140_ (
    .A(_032_),
    .B(bcsctl1[3]),
    .Y(bcsctl1_rd[11])
  );
  \$_AND_  _141_ (
    .A(_032_),
    .B(bcsctl1[4]),
    .Y(bcsctl1_rd[12])
  );
  \$_AND_  _142_ (
    .A(_032_),
    .B(bcsctl1[5]),
    .Y(bcsctl1_rd[13])
  );
  \$_AND_  _143_ (
    .A(_032_),
    .B(bcsctl1[6]),
    .Y(bcsctl1_rd[14])
  );
  \$_AND_  _144_ (
    .A(_032_),
    .B(bcsctl1[7]),
    .Y(bcsctl1_rd[15])
  );
  \$_OR_  _145_ (
    .A(per_addr[0]),
    .B(_006_),
    .Y(_033_)
  );
  \$_OR_  _146_ (
    .A(_033_),
    .B(per_addr[1]),
    .Y(_034_)
  );
  \$_INV_  _147_ (
    .A(_034_),
    .Y(_035_)
  );
  \$_AND_  _148_ (
    .A(_035_),
    .B(_031_),
    .Y(_036_)
  );
  \$_AND_  _149_ (
    .A(_036_),
    .B(bcsctl2[0]),
    .Y(bcsctl2_rd[0])
  );
  \$_AND_  _150_ (
    .A(_036_),
    .B(bcsctl2[1]),
    .Y(bcsctl2_rd[1])
  );
  \$_AND_  _151_ (
    .A(_036_),
    .B(bcsctl2[2]),
    .Y(bcsctl2_rd[2])
  );
  \$_AND_  _152_ (
    .A(_036_),
    .B(bcsctl2[3]),
    .Y(bcsctl2_rd[3])
  );
  \$_AND_  _153_ (
    .A(_036_),
    .B(bcsctl2[4]),
    .Y(bcsctl2_rd[4])
  );
  \$_AND_  _154_ (
    .A(_036_),
    .B(bcsctl2[5]),
    .Y(bcsctl2_rd[5])
  );
  \$_AND_  _155_ (
    .A(_036_),
    .B(bcsctl2[6]),
    .Y(bcsctl2_rd[6])
  );
  \$_AND_  _156_ (
    .A(_036_),
    .B(bcsctl2[7]),
    .Y(bcsctl2_rd[7])
  );
  \$_OR_  _157_ (
    .A(bcsctl1[5]),
    .B(bcsctl1[4]),
    .Y(_037_)
  );
  \$_INV_  _158_ (
    .A(_037_),
    .Y(_038_)
  );
  \$_INV_  _159_ (
    .A(bcsctl1[5]),
    .Y(_039_)
  );
  \$_AND_  _160_ (
    .A(_039_),
    .B(bcsctl1[4]),
    .Y(_040_)
  );
  \$_INV_  _161_ (
    .A(bcsctl1[4]),
    .Y(_041_)
  );
  \$_AND_  _162_ (
    .A(bcsctl1[5]),
    .B(_041_),
    .Y(_042_)
  );
  \$_AND_  _163_ (
    .A(aclk_div[1]),
    .B(aclk_div[0]),
    .Y(_043_)
  );
  \$_AND_  _164_ (
    .A(_043_),
    .B(_042_),
    .Y(_044_)
  );
  \$_OR_  _165_ (
    .A(_039_),
    .B(bcsctl1[4]),
    .Y(_045_)
  );
  \$_AND_  _166_ (
    .A(_045_),
    .B(aclk_div[2]),
    .Y(_046_)
  );
  \$_AND_  _167_ (
    .A(_046_),
    .B(_043_),
    .Y(_047_)
  );
  \$_OR_  _168_ (
    .A(_047_),
    .B(_044_),
    .Y(_048_)
  );
  \$_MUX_  _169_ (
    .A(_048_),
    .B(aclk_div[0]),
    .S(_040_),
    .Y(_049_)
  );
  \$_OR_  _170_ (
    .A(_049_),
    .B(_038_),
    .Y(_050_)
  );
  \$_INV_  _171_ (
    .A(oscoff),
    .Y(_051_)
  );
  \$_OR_  _172_ (
    .A(_051_),
    .B(bcsctl2[3]),
    .Y(_052_)
  );
  \$_INV_  _173_ (
    .A(lfxt_clk_dly),
    .Y(_053_)
  );
  \$_AND_  _174_ (
    .A(_053_),
    .B(lfxt_clk_s),
    .Y(_054_)
  );
  \$_AND_  _175_ (
    .A(_054_),
    .B(_052_),
    .Y(_055_)
  );
  \$_AND_  _176_ (
    .A(_055_),
    .B(cpu_en),
    .Y(_056_)
  );
  \$_AND_  _177_ (
    .A(_056_),
    .B(_050_),
    .Y(_001_)
  );
  \$_OR_  _178_ (
    .A(bcsctl2[2]),
    .B(bcsctl2[1]),
    .Y(_057_)
  );
  \$_INV_  _179_ (
    .A(_057_),
    .Y(_058_)
  );
  \$_INV_  _180_ (
    .A(bcsctl2[2]),
    .Y(_059_)
  );
  \$_AND_  _181_ (
    .A(_059_),
    .B(bcsctl2[1]),
    .Y(_060_)
  );
  \$_INV_  _182_ (
    .A(bcsctl2[1]),
    .Y(_061_)
  );
  \$_AND_  _183_ (
    .A(bcsctl2[2]),
    .B(_061_),
    .Y(_062_)
  );
  \$_AND_  _184_ (
    .A(smclk_div[1]),
    .B(smclk_div[0]),
    .Y(_063_)
  );
  \$_AND_  _185_ (
    .A(_063_),
    .B(_062_),
    .Y(_064_)
  );
  \$_OR_  _186_ (
    .A(_059_),
    .B(bcsctl2[1]),
    .Y(_065_)
  );
  \$_AND_  _187_ (
    .A(_065_),
    .B(smclk_div[2]),
    .Y(_066_)
  );
  \$_AND_  _188_ (
    .A(_066_),
    .B(_063_),
    .Y(_067_)
  );
  \$_OR_  _189_ (
    .A(_067_),
    .B(_064_),
    .Y(_068_)
  );
  \$_MUX_  _190_ (
    .A(_068_),
    .B(smclk_div[0]),
    .S(_060_),
    .Y(_069_)
  );
  \$_OR_  _191_ (
    .A(_069_),
    .B(_058_),
    .Y(_070_)
  );
  \$_INV_  _192_ (
    .A(scg1),
    .Y(_071_)
  );
  \$_INV_  _193_ (
    .A(bcsctl2[3]),
    .Y(_072_)
  );
  \$_OR_  _194_ (
    .A(_055_),
    .B(_072_),
    .Y(_073_)
  );
  \$_AND_  _195_ (
    .A(_073_),
    .B(_071_),
    .Y(_074_)
  );
  \$_AND_  _196_ (
    .A(_074_),
    .B(cpu_en),
    .Y(_075_)
  );
  \$_AND_  _197_ (
    .A(_075_),
    .B(_070_),
    .Y(_005_)
  );
  \$_INV_  _198_ (
    .A(reset_n),
    .Y(por_a)
  );
  \$_INV_  _199_ (
    .A(dbg_cpu_reset),
    .Y(_076_)
  );
  \$_INV_  _200_ (
    .A(dbg_rst),
    .Y(_077_)
  );
  \$_INV_  _201_ (
    .A(dbg_en),
    .Y(dbg_rst_nxt)
  );
  \$_OR_  _202_ (
    .A(dbg_rst_nxt),
    .B(_077_),
    .Y(_078_)
  );
  \$_OR_  _203_ (
    .A(_078_),
    .B(puc_noscan_n),
    .Y(_079_)
  );
  \$_AND_  _204_ (
    .A(_079_),
    .B(_076_),
    .Y(_108_)
  );
  \$_OR_  _205_ (
    .A(por),
    .B(wdt_reset),
    .Y(puc_a)
  );
  \$_INV_  _206_ (
    .A(_012_),
    .Y(_080_)
  );
  \$_OR_  _207_ (
    .A(per_addr[8]),
    .B(per_addr[7]),
    .Y(_081_)
  );
  \$_OR_  _208_ (
    .A(per_addr[10]),
    .B(per_addr[9]),
    .Y(_082_)
  );
  \$_OR_  _209_ (
    .A(_082_),
    .B(_081_),
    .Y(_083_)
  );
  \$_INV_  _210_ (
    .A(per_en),
    .Y(_084_)
  );
  \$_OR_  _211_ (
    .A(per_addr[13]),
    .B(_084_),
    .Y(_085_)
  );
  \$_OR_  _212_ (
    .A(per_addr[6]),
    .B(per_addr[4]),
    .Y(_086_)
  );
  \$_OR_  _213_ (
    .A(_086_),
    .B(_085_),
    .Y(_087_)
  );
  \$_OR_  _214_ (
    .A(_087_),
    .B(_083_),
    .Y(_088_)
  );
  \$_OR_  _215_ (
    .A(_088_),
    .B(_080_),
    .Y(_089_)
  );
  \$_INV_  _216_ (
    .A(_008_),
    .Y(_090_)
  );
  \$_OR_  _217_ (
    .A(_090_),
    .B(_029_),
    .Y(_091_)
  );
  \$_OR_  _218_ (
    .A(_091_),
    .B(_089_),
    .Y(_092_)
  );
  \$_AND_  _219_ (
    .A(_092_),
    .B(bcsctl1[0]),
    .Y(_002_[0])
  );
  \$_AND_  _220_ (
    .A(_092_),
    .B(bcsctl1[1]),
    .Y(_002_[1])
  );
  \$_AND_  _221_ (
    .A(_092_),
    .B(bcsctl1[2]),
    .Y(_002_[2])
  );
  \$_AND_  _222_ (
    .A(_092_),
    .B(bcsctl1[3]),
    .Y(_002_[3])
  );
  \$_MUX_  _223_ (
    .A(per_din[12]),
    .B(bcsctl1[4]),
    .S(_092_),
    .Y(_002_[4])
  );
  \$_MUX_  _224_ (
    .A(per_din[13]),
    .B(bcsctl1[5]),
    .S(_092_),
    .Y(_002_[5])
  );
  \$_AND_  _225_ (
    .A(_092_),
    .B(bcsctl1[6]),
    .Y(_002_[6])
  );
  \$_AND_  _226_ (
    .A(_092_),
    .B(bcsctl1[7]),
    .Y(_002_[7])
  );
  \$_OR_  _227_ (
    .A(_034_),
    .B(_028_),
    .Y(_093_)
  );
  \$_OR_  _228_ (
    .A(_093_),
    .B(_089_),
    .Y(_094_)
  );
  \$_AND_  _229_ (
    .A(_094_),
    .B(bcsctl2[0]),
    .Y(_003_[0])
  );
  \$_MUX_  _230_ (
    .A(per_din[1]),
    .B(bcsctl2[1]),
    .S(_094_),
    .Y(_003_[1])
  );
  \$_MUX_  _231_ (
    .A(per_din[2]),
    .B(bcsctl2[2]),
    .S(_094_),
    .Y(_003_[2])
  );
  \$_MUX_  _232_ (
    .A(per_din[3]),
    .B(bcsctl2[3]),
    .S(_094_),
    .Y(_003_[3])
  );
  \$_AND_  _233_ (
    .A(_094_),
    .B(bcsctl2[4]),
    .Y(_003_[4])
  );
  \$_AND_  _234_ (
    .A(_094_),
    .B(bcsctl2[5]),
    .Y(_003_[5])
  );
  \$_AND_  _235_ (
    .A(_094_),
    .B(bcsctl2[6]),
    .Y(_003_[6])
  );
  \$_AND_  _236_ (
    .A(_094_),
    .B(bcsctl2[7]),
    .Y(_003_[7])
  );
  \$_AND_  _237_ (
    .A(_055_),
    .B(_037_),
    .Y(_095_)
  );
  \$_XOR_  _238_ (
    .A(_095_),
    .B(aclk_div[0]),
    .Y(_000_[0])
  );
  \$_XOR_  _239_ (
    .A(aclk_div[1]),
    .B(aclk_div[0]),
    .Y(_096_)
  );
  \$_MUX_  _240_ (
    .A(aclk_div[1]),
    .B(_096_),
    .S(_095_),
    .Y(_000_[1])
  );
  \$_XOR_  _241_ (
    .A(_043_),
    .B(aclk_div[2]),
    .Y(_097_)
  );
  \$_MUX_  _242_ (
    .A(aclk_div[2]),
    .B(_097_),
    .S(_095_),
    .Y(_000_[2])
  );
  \$_AND_  _243_ (
    .A(_074_),
    .B(_057_),
    .Y(_098_)
  );
  \$_XOR_  _244_ (
    .A(_098_),
    .B(smclk_div[0]),
    .Y(_004_[0])
  );
  \$_AND_  _245_ (
    .A(oscoff),
    .B(_072_),
    .Y(_099_)
  );
  \$_INV_  _246_ (
    .A(lfxt_clk_s),
    .Y(_100_)
  );
  \$_OR_  _247_ (
    .A(lfxt_clk_dly),
    .B(_100_),
    .Y(_101_)
  );
  \$_OR_  _248_ (
    .A(_101_),
    .B(_099_),
    .Y(_102_)
  );
  \$_AND_  _249_ (
    .A(_102_),
    .B(bcsctl2[3]),
    .Y(_103_)
  );
  \$_OR_  _250_ (
    .A(_103_),
    .B(scg1),
    .Y(_104_)
  );
  \$_OR_  _251_ (
    .A(_104_),
    .B(_058_),
    .Y(_105_)
  );
  \$_XOR_  _252_ (
    .A(smclk_div[1]),
    .B(smclk_div[0]),
    .Y(_106_)
  );
  \$_MUX_  _253_ (
    .A(_106_),
    .B(smclk_div[1]),
    .S(_105_),
    .Y(_004_[1])
  );
  \$_XOR_  _254_ (
    .A(_063_),
    .B(smclk_div[2]),
    .Y(_107_)
  );
  \$_MUX_  _255_ (
    .A(_107_),
    .B(smclk_div[2]),
    .S(_105_),
    .Y(_004_[2])
  );
  \$_DFF_PP0_  \bcsctl1_reg[0]  /* _256_ */ (
    .C(dco_clk),
    .D(_002_[0]),
    .Q(bcsctl1[0]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[1]  /* _257_ */ (
    .C(dco_clk),
    .D(_002_[1]),
    .Q(bcsctl1[1]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[2]  /* _258_ */ (
    .C(dco_clk),
    .D(_002_[2]),
    .Q(bcsctl1[2]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[3]  /* _259_ */ (
    .C(dco_clk),
    .D(_002_[3]),
    .Q(bcsctl1[3]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[4]  /* _260_ */ (
    .C(dco_clk),
    .D(_002_[4]),
    .Q(bcsctl1[4]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[5]  /* _261_ */ (
    .C(dco_clk),
    .D(_002_[5]),
    .Q(bcsctl1[5]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[6]  /* _262_ */ (
    .C(dco_clk),
    .D(_002_[6]),
    .Q(bcsctl1[6]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl1_reg[7]  /* _263_ */ (
    .C(dco_clk),
    .D(_002_[7]),
    .Q(bcsctl1[7]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[0]  /* _264_ */ (
    .C(dco_clk),
    .D(_003_[0]),
    .Q(bcsctl2[0]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[1]  /* _265_ */ (
    .C(dco_clk),
    .D(_003_[1]),
    .Q(bcsctl2[1]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[2]  /* _266_ */ (
    .C(dco_clk),
    .D(_003_[2]),
    .Q(bcsctl2[2]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[3]  /* _267_ */ (
    .C(dco_clk),
    .D(_003_[3]),
    .Q(bcsctl2[3]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[4]  /* _268_ */ (
    .C(dco_clk),
    .D(_003_[4]),
    .Q(bcsctl2[4]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[5]  /* _269_ */ (
    .C(dco_clk),
    .D(_003_[5]),
    .Q(bcsctl2[5]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[6]  /* _270_ */ (
    .C(dco_clk),
    .D(_003_[6]),
    .Q(bcsctl2[6]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \bcsctl2_reg[7]  /* _271_ */ (
    .C(dco_clk),
    .D(_003_[7]),
    .Q(bcsctl2[7]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  lfxt_clk_dly_reg /* _272_ */ (
    .C(dco_clk),
    .D(lfxt_clk_s),
    .Q(lfxt_clk_dly),
    .R(por)
  );
  \$_DFF_PP0_  \aclk_div_reg[0]  /* _273_ */ (
    .C(dco_clk),
    .D(_000_[0]),
    .Q(aclk_div[0]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \aclk_div_reg[1]  /* _274_ */ (
    .C(dco_clk),
    .D(_000_[1]),
    .Q(aclk_div[1]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \aclk_div_reg[2]  /* _275_ */ (
    .C(dco_clk),
    .D(_000_[2]),
    .Q(aclk_div[2]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  aclk_en_reg /* _276_ */ (
    .C(dco_clk),
    .D(_001_),
    .Q(aclk_en),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  smclk_en_reg /* _277_ */ (
    .C(dco_clk),
    .D(_005_),
    .Q(smclk_en),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \smclk_div_reg[0]  /* _278_ */ (
    .C(dco_clk),
    .D(_004_[0]),
    .Q(smclk_div[0]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \smclk_div_reg[1]  /* _279_ */ (
    .C(dco_clk),
    .D(_004_[1]),
    .Q(smclk_div[1]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP0_  \smclk_div_reg[2]  /* _280_ */ (
    .C(dco_clk),
    .D(_004_[2]),
    .Q(smclk_div[2]),
    .R(puc_pnd_set)
  );
  \$_DFF_PP1_  dbg_rst_reg /* _281_ */ (
    .C(dco_clk),
    .D(dbg_rst_nxt),
    .Q(dbg_rst),
    .R(por)
  );
  omsp_sync_cell sync_cell_lfxt_clk (
    .clk(dco_clk),
    .data_in(lfxt_clk),
    .data_out(lfxt_clk_s),
    .rst(por)
  );
  omsp_sync_cell sync_cell_puc (
    .clk(dco_clk),
    .data_in(_108_),
    .data_out(puc_noscan_n),
    .rst(puc_a)
  );
  omsp_sync_reset sync_reset_por (
    .clk(dco_clk),
    .rst_a(por_a),
    .rst_s(por)
  );
  assign aclk = dco_clk;
  assign bcsctl1_nxt = per_din[15:8];
  assign bcsctl1_rd[7:0] = 8'b00000000;
  assign bcsctl2_nxt = per_din[7:0];
  assign bcsctl2_rd[15:8] = 8'b00000000;
  assign cpu_en_aux_s = cpu_en;
  assign cpu_en_s = cpu_en;
  assign dbg_clk = dco_clk;
  assign dbg_en_s = dbg_en;
  assign dbg_rst_noscan = dbg_rst;
  assign dco_enable = 1'b1;
  assign dco_wkup = 1'b1;
  assign lfxt_enable = 1'b1;
  assign lfxt_wkup = 1'b0;
  assign mclk = dco_clk;
  assign nodiv_mclk = dco_clk;
  assign nodiv_smclk = dco_clk;
  assign per_dout = { bcsctl1_rd[15:8], bcsctl2_rd[7:0] };
  assign por_noscan = por;
  assign puc_a_scan = puc_a;
  assign puc_rst = puc_pnd_set;
  assign reg_addr = { 1'b0, per_addr[2:0] };
  assign smclk = dco_clk;
endmodule

module omsp_dbg(dbg_freeze, dbg_halt_cmd, dbg_mem_addr, dbg_mem_dout, dbg_mem_en, dbg_mem_wr, dbg_reg_wr, dbg_cpu_reset, dbg_uart_txd, cpu_en_s, cpu_id, dbg_clk, dbg_en_s, dbg_halt_st, dbg_mem_din, dbg_reg_din, dbg_rst, dbg_uart_rxd, decode_noirq, eu_mab, eu_mb_en, eu_mb_wr, eu_mdb_in, eu_mdb_out, exec_done, fe_mb_en, fe_mdb_in, pc, puc_pnd_set);
  wire [3:0] _0000_;
  wire [1:0] _0001_;
  wire _0002_;
  wire _0003_;
  wire [1:0] _0004_;
  wire [15:0] _0005_;
  wire _0006_;
  wire [15:0] _0007_;
  wire [2:0] _0008_;
  wire [15:0] _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire [6:3] cpu_ctl;
  wire [7:0] cpu_ctl_full;
  input cpu_en_s;
  input [31:0] cpu_id;
  wire [3:2] cpu_stat;
  wire [7:0] cpu_stat_full;
  wire [3:2] cpu_stat_set;
  wire [5:0] dbg_addr;
  input dbg_clk;
  output dbg_cpu_reset;
  wire [15:0] dbg_din;
  wire [15:0] dbg_dout;
  input dbg_en_s;
  output dbg_freeze;
  output dbg_halt_cmd;
  input dbg_halt_st;
  output [15:0] dbg_mem_addr;
  input [15:0] dbg_mem_din;
  output [15:0] dbg_mem_dout;
  output dbg_mem_en;
  wire dbg_mem_rd;
  wire dbg_mem_rd_dly;
  output [1:0] dbg_mem_wr;
  wire dbg_rd;
  wire dbg_rd_rdy;
  input [15:0] dbg_reg_din;
  output dbg_reg_wr;
  input dbg_rst;
  input dbg_uart_rxd;
  output dbg_uart_txd;
  wire dbg_wr;
  input decode_noirq;
  input [15:0] eu_mab;
  input eu_mb_en;
  input [1:0] eu_mb_wr;
  input [15:0] eu_mdb_in;
  input [15:0] eu_mdb_out;
  input exec_done;
  input fe_mb_en;
  input [15:0] fe_mdb_in;
  wire halt_flag;
  wire [1:0] inc_step;
  wire [15:0] mem_addr;
  wire mem_burst;
  wire mem_burst_end;
  wire mem_burst_rd;
  wire mem_burst_wr;
  wire mem_bw;
  wire [15:0] mem_cnt;
  wire [3:1] mem_ctl;
  wire [7:0] mem_ctl_full;
  wire [15:0] mem_data;
  wire mem_start;
  wire mem_startb;
  wire [2:0] mem_state;
  input [15:0] pc;
  input puc_pnd_set;
  wire reg_write;
  \$_OR_  _0539_ (
    .A(dbg_addr[1]),
    .B(mem_burst),
    .Y(_0012_)
  );
  \$_INV_  _0540_ (
    .A(_0012_),
    .Y(_0013_)
  );
  \$_INV_  _0541_ (
    .A(mem_burst),
    .Y(_0014_)
  );
  \$_AND_  _0542_ (
    .A(dbg_addr[0]),
    .B(_0014_),
    .Y(_0015_)
  );
  \$_INV_  _0543_ (
    .A(_0015_),
    .Y(_0016_)
  );
  \$_AND_  _0544_ (
    .A(_0016_),
    .B(_0013_),
    .Y(_0017_)
  );
  \$_OR_  _0545_ (
    .A(dbg_addr[2]),
    .B(mem_burst),
    .Y(_0018_)
  );
  \$_AND_  _0546_ (
    .A(dbg_addr[3]),
    .B(_0014_),
    .Y(_0019_)
  );
  \$_AND_  _0547_ (
    .A(dbg_addr[5]),
    .B(_0014_),
    .Y(_0020_)
  );
  \$_AND_  _0548_ (
    .A(dbg_addr[4]),
    .B(_0014_),
    .Y(_0021_)
  );
  \$_OR_  _0549_ (
    .A(_0021_),
    .B(_0020_),
    .Y(_0022_)
  );
  \$_OR_  _0550_ (
    .A(_0022_),
    .B(_0019_),
    .Y(_0023_)
  );
  \$_INV_  _0551_ (
    .A(_0023_),
    .Y(_0024_)
  );
  \$_AND_  _0552_ (
    .A(_0024_),
    .B(_0018_),
    .Y(_0025_)
  );
  \$_AND_  _0553_ (
    .A(_0025_),
    .B(_0017_),
    .Y(_0026_)
  );
  \$_OR_  _0554_ (
    .A(_0023_),
    .B(_0018_),
    .Y(_0027_)
  );
  \$_INV_  _0555_ (
    .A(_0027_),
    .Y(_0028_)
  );
  \$_AND_  _0556_ (
    .A(_0015_),
    .B(_0012_),
    .Y(_0029_)
  );
  \$_AND_  _0557_ (
    .A(_0029_),
    .B(_0028_),
    .Y(_0030_)
  );
  \$_AND_  _0558_ (
    .A(_0015_),
    .B(_0013_),
    .Y(_0031_)
  );
  \$_AND_  _0559_ (
    .A(_0031_),
    .B(_0025_),
    .Y(_0032_)
  );
  \$_AND_  _0560_ (
    .A(_0016_),
    .B(_0012_),
    .Y(_0033_)
  );
  \$_AND_  _0561_ (
    .A(_0033_),
    .B(_0025_),
    .Y(_0034_)
  );
  \$_AND_  _0562_ (
    .A(_0029_),
    .B(_0025_),
    .Y(_0035_)
  );
  \$_AND_  _0563_ (
    .A(_0028_),
    .B(_0017_),
    .Y(_0036_)
  );
  \$_AND_  _0564_ (
    .A(_0031_),
    .B(_0028_),
    .Y(_0037_)
  );
  \$_AND_  _0565_ (
    .A(_0033_),
    .B(_0028_),
    .Y(_0038_)
  );
  \$_AND_  _0566_ (
    .A(_0026_),
    .B(dbg_wr),
    .Y(_0039_)
  );
  \$_AND_  _0567_ (
    .A(_0039_),
    .B(dbg_din[0]),
    .Y(_0010_)
  );
  \$_INV_  _0568_ (
    .A(cpu_en_s),
    .Y(_0040_)
  );
  \$_OR_  _0569_ (
    .A(_0040_),
    .B(cpu_ctl[4]),
    .Y(_0041_)
  );
  \$_AND_  _0570_ (
    .A(_0041_),
    .B(dbg_halt_st),
    .Y(dbg_freeze)
  );
  \$_INV_  _0571_ (
    .A(inc_step[1]),
    .Y(_0042_)
  );
  \$_AND_  _0572_ (
    .A(_0038_),
    .B(dbg_wr),
    .Y(_0043_)
  );
  \$_INV_  _0573_ (
    .A(dbg_halt_st),
    .Y(_0044_)
  );
  \$_AND_  _0574_ (
    .A(_0044_),
    .B(dbg_din[0]),
    .Y(_0045_)
  );
  \$_AND_  _0575_ (
    .A(_0045_),
    .B(_0043_),
    .Y(_0046_)
  );
  \$_OR_  _0576_ (
    .A(mem_cnt[14]),
    .B(mem_cnt[13]),
    .Y(_0047_)
  );
  \$_OR_  _0577_ (
    .A(mem_cnt[1]),
    .B(mem_cnt[15]),
    .Y(_0048_)
  );
  \$_OR_  _0578_ (
    .A(_0048_),
    .B(_0047_),
    .Y(_0049_)
  );
  \$_OR_  _0579_ (
    .A(mem_cnt[10]),
    .B(mem_cnt[0]),
    .Y(_0050_)
  );
  \$_OR_  _0580_ (
    .A(mem_cnt[12]),
    .B(mem_cnt[11]),
    .Y(_0051_)
  );
  \$_OR_  _0581_ (
    .A(_0051_),
    .B(_0050_),
    .Y(_0052_)
  );
  \$_OR_  _0582_ (
    .A(_0052_),
    .B(_0049_),
    .Y(_0053_)
  );
  \$_OR_  _0583_ (
    .A(mem_cnt[7]),
    .B(mem_cnt[6]),
    .Y(_0054_)
  );
  \$_OR_  _0584_ (
    .A(mem_cnt[9]),
    .B(mem_cnt[8]),
    .Y(_0055_)
  );
  \$_OR_  _0585_ (
    .A(_0055_),
    .B(_0054_),
    .Y(_0056_)
  );
  \$_OR_  _0586_ (
    .A(mem_cnt[3]),
    .B(mem_cnt[2]),
    .Y(_0057_)
  );
  \$_OR_  _0587_ (
    .A(mem_cnt[5]),
    .B(mem_cnt[4]),
    .Y(_0058_)
  );
  \$_OR_  _0588_ (
    .A(_0058_),
    .B(_0057_),
    .Y(_0059_)
  );
  \$_OR_  _0589_ (
    .A(_0059_),
    .B(_0056_),
    .Y(_0060_)
  );
  \$_OR_  _0590_ (
    .A(_0060_),
    .B(_0053_),
    .Y(_0061_)
  );
  \$_INV_  _0591_ (
    .A(_0061_),
    .Y(_0062_)
  );
  \$_AND_  _0592_ (
    .A(_0062_),
    .B(mem_start),
    .Y(_0063_)
  );
  \$_OR_  _0593_ (
    .A(_0063_),
    .B(mem_startb),
    .Y(_0064_)
  );
  \$_INV_  _0594_ (
    .A(mem_state[2]),
    .Y(_0065_)
  );
  \$_INV_  _0595_ (
    .A(mem_state[0]),
    .Y(_0066_)
  );
  \$_INV_  _0596_ (
    .A(mem_state[1]),
    .Y(_0067_)
  );
  \$_AND_  _0597_ (
    .A(_0067_),
    .B(_0066_),
    .Y(_0068_)
  );
  \$_AND_  _0598_ (
    .A(_0068_),
    .B(_0065_),
    .Y(_0069_)
  );
  \$_AND_  _0599_ (
    .A(_0069_),
    .B(dbg_halt_st),
    .Y(_0070_)
  );
  \$_AND_  _0600_ (
    .A(_0070_),
    .B(_0064_),
    .Y(_0537_)
  );
  \$_AND_  _0601_ (
    .A(mem_state[1]),
    .B(_0044_),
    .Y(_0071_)
  );
  \$_AND_  _0602_ (
    .A(_0069_),
    .B(_0044_),
    .Y(_0072_)
  );
  \$_AND_  _0603_ (
    .A(_0072_),
    .B(_0064_),
    .Y(_0073_)
  );
  \$_OR_  _0604_ (
    .A(_0073_),
    .B(_0071_),
    .Y(_0538_)
  );
  \$_OR_  _0605_ (
    .A(_0538_),
    .B(_0537_),
    .Y(_0074_)
  );
  \$_AND_  _0606_ (
    .A(mem_state[1]),
    .B(dbg_halt_st),
    .Y(_0536_)
  );
  \$_OR_  _0607_ (
    .A(_0536_),
    .B(_0537_),
    .Y(_0075_)
  );
  \$_AND_  _0608_ (
    .A(dbg_en_s),
    .B(cpu_ctl[5]),
    .Y(_0076_)
  );
  \$_AND_  _0609_ (
    .A(_0076_),
    .B(puc_pnd_set),
    .Y(_0077_)
  );
  \$_AND_  _0610_ (
    .A(decode_noirq),
    .B(cpu_ctl[3]),
    .Y(_0078_)
  );
  \$_INV_  _0611_ (
    .A(fe_mdb_in[10]),
    .Y(_0079_)
  );
  \$_INV_  _0612_ (
    .A(fe_mdb_in[11]),
    .Y(_0080_)
  );
  \$_AND_  _0613_ (
    .A(_0080_),
    .B(_0079_),
    .Y(_0081_)
  );
  \$_INV_  _0614_ (
    .A(fe_mdb_in[12]),
    .Y(_0082_)
  );
  \$_INV_  _0615_ (
    .A(fe_mdb_in[13]),
    .Y(_0083_)
  );
  \$_AND_  _0616_ (
    .A(_0083_),
    .B(_0082_),
    .Y(_0084_)
  );
  \$_AND_  _0617_ (
    .A(_0084_),
    .B(_0081_),
    .Y(_0085_)
  );
  \$_AND_  _0618_ (
    .A(_0085_),
    .B(_0078_),
    .Y(_0086_)
  );
  \$_AND_  _0619_ (
    .A(fe_mdb_in[6]),
    .B(fe_mdb_in[1]),
    .Y(_0087_)
  );
  \$_AND_  _0620_ (
    .A(fe_mdb_in[9]),
    .B(fe_mdb_in[8]),
    .Y(_0088_)
  );
  \$_AND_  _0621_ (
    .A(_0088_),
    .B(_0087_),
    .Y(_0089_)
  );
  \$_INV_  _0622_ (
    .A(fe_mdb_in[5]),
    .Y(_0090_)
  );
  \$_INV_  _0623_ (
    .A(fe_mdb_in[7]),
    .Y(_0091_)
  );
  \$_AND_  _0624_ (
    .A(_0091_),
    .B(_0090_),
    .Y(_0092_)
  );
  \$_AND_  _0625_ (
    .A(fe_mdb_in[14]),
    .B(fe_mdb_in[0]),
    .Y(_0093_)
  );
  \$_AND_  _0626_ (
    .A(_0093_),
    .B(_0092_),
    .Y(_0094_)
  );
  \$_INV_  _0627_ (
    .A(fe_mdb_in[15]),
    .Y(_0095_)
  );
  \$_INV_  _0628_ (
    .A(fe_mdb_in[2]),
    .Y(_0096_)
  );
  \$_AND_  _0629_ (
    .A(_0096_),
    .B(_0095_),
    .Y(_0097_)
  );
  \$_INV_  _0630_ (
    .A(fe_mdb_in[3]),
    .Y(_0098_)
  );
  \$_INV_  _0631_ (
    .A(fe_mdb_in[4]),
    .Y(_0099_)
  );
  \$_AND_  _0632_ (
    .A(_0099_),
    .B(_0098_),
    .Y(_0100_)
  );
  \$_AND_  _0633_ (
    .A(_0100_),
    .B(_0097_),
    .Y(_0101_)
  );
  \$_AND_  _0634_ (
    .A(_0101_),
    .B(_0094_),
    .Y(_0102_)
  );
  \$_AND_  _0635_ (
    .A(_0102_),
    .B(_0089_),
    .Y(_0103_)
  );
  \$_AND_  _0636_ (
    .A(_0103_),
    .B(_0086_),
    .Y(_0104_)
  );
  \$_OR_  _0637_ (
    .A(_0104_),
    .B(_0077_),
    .Y(_0105_)
  );
  \$_OR_  _0638_ (
    .A(_0105_),
    .B(_0073_),
    .Y(_0106_)
  );
  \$_OR_  _0639_ (
    .A(_0106_),
    .B(_0046_),
    .Y(_0107_)
  );
  \$_OR_  _0640_ (
    .A(_0107_),
    .B(halt_flag),
    .Y(_0108_)
  );
  \$_AND_  _0641_ (
    .A(_0108_),
    .B(_0042_),
    .Y(dbg_halt_cmd)
  );
  \$_INV_  _0642_ (
    .A(dbg_wr),
    .Y(_0109_)
  );
  \$_INV_  _0643_ (
    .A(dbg_rd_rdy),
    .Y(_0110_)
  );
  \$_AND_  _0644_ (
    .A(_0110_),
    .B(_0109_),
    .Y(_0111_)
  );
  \$_OR_  _0645_ (
    .A(_0111_),
    .B(_0061_),
    .Y(_0112_)
  );
  \$_INV_  _0646_ (
    .A(_0112_),
    .Y(mem_burst_end)
  );
  \$_INV_  _0647_ (
    .A(mem_ctl[1]),
    .Y(_0113_)
  );
  \$_AND_  _0648_ (
    .A(_0061_),
    .B(mem_start),
    .Y(_0114_)
  );
  \$_AND_  _0649_ (
    .A(_0114_),
    .B(_0113_),
    .Y(mem_burst_rd)
  );
  \$_AND_  _0650_ (
    .A(_0114_),
    .B(mem_ctl[1]),
    .Y(mem_burst_wr)
  );
  \$_OR_  _0651_ (
    .A(mem_state[2]),
    .B(mem_state[0]),
    .Y(_0115_)
  );
  \$_AND_  _0652_ (
    .A(mem_ctl[1]),
    .B(mem_ctl[2]),
    .Y(_0116_)
  );
  \$_AND_  _0653_ (
    .A(_0116_),
    .B(_0115_),
    .Y(dbg_reg_wr)
  );
  \$_INV_  _0654_ (
    .A(mem_ctl[2]),
    .Y(_0117_)
  );
  \$_AND_  _0655_ (
    .A(_0115_),
    .B(_0117_),
    .Y(dbg_mem_en)
  );
  \$_AND_  _0656_ (
    .A(dbg_mem_en),
    .B(_0113_),
    .Y(dbg_mem_rd)
  );
  \$_AND_  _0657_ (
    .A(dbg_mem_en),
    .B(mem_ctl[1]),
    .Y(_0118_)
  );
  \$_INV_  _0658_ (
    .A(dbg_mem_addr[0]),
    .Y(_0119_)
  );
  \$_INV_  _0659_ (
    .A(mem_bw),
    .Y(_0120_)
  );
  \$_OR_  _0660_ (
    .A(_0120_),
    .B(_0119_),
    .Y(_0121_)
  );
  \$_AND_  _0661_ (
    .A(_0121_),
    .B(_0118_),
    .Y(dbg_mem_wr[0])
  );
  \$_OR_  _0662_ (
    .A(_0120_),
    .B(dbg_mem_addr[0]),
    .Y(_0122_)
  );
  \$_AND_  _0663_ (
    .A(_0122_),
    .B(_0118_),
    .Y(dbg_mem_wr[1])
  );
  \$_AND_  _0664_ (
    .A(_0036_),
    .B(cpu_id[0]),
    .Y(_0123_)
  );
  \$_AND_  _0665_ (
    .A(_0037_),
    .B(cpu_id[16]),
    .Y(_0124_)
  );
  \$_OR_  _0666_ (
    .A(_0124_),
    .B(_0123_),
    .Y(_0125_)
  );
  \$_AND_  _0667_ (
    .A(_0030_),
    .B(dbg_halt_st),
    .Y(_0126_)
  );
  \$_AND_  _0668_ (
    .A(_0034_),
    .B(mem_data[0]),
    .Y(_0127_)
  );
  \$_OR_  _0669_ (
    .A(_0127_),
    .B(_0126_),
    .Y(_0128_)
  );
  \$_AND_  _0670_ (
    .A(_0032_),
    .B(dbg_mem_addr[0]),
    .Y(_0129_)
  );
  \$_AND_  _0671_ (
    .A(_0035_),
    .B(mem_cnt[0]),
    .Y(_0130_)
  );
  \$_OR_  _0672_ (
    .A(_0130_),
    .B(_0129_),
    .Y(_0131_)
  );
  \$_OR_  _0673_ (
    .A(_0131_),
    .B(_0128_),
    .Y(_0132_)
  );
  \$_OR_  _0674_ (
    .A(_0132_),
    .B(_0125_),
    .Y(dbg_dout[0])
  );
  \$_AND_  _0675_ (
    .A(_0036_),
    .B(cpu_id[10]),
    .Y(_0133_)
  );
  \$_AND_  _0676_ (
    .A(_0037_),
    .B(cpu_id[26]),
    .Y(_0134_)
  );
  \$_OR_  _0677_ (
    .A(_0134_),
    .B(_0133_),
    .Y(_0135_)
  );
  \$_AND_  _0678_ (
    .A(_0035_),
    .B(mem_cnt[10]),
    .Y(_0136_)
  );
  \$_AND_  _0679_ (
    .A(_0034_),
    .B(mem_data[10]),
    .Y(_0137_)
  );
  \$_AND_  _0680_ (
    .A(_0032_),
    .B(dbg_mem_addr[10]),
    .Y(_0138_)
  );
  \$_OR_  _0681_ (
    .A(_0138_),
    .B(_0137_),
    .Y(_0139_)
  );
  \$_OR_  _0682_ (
    .A(_0139_),
    .B(_0136_),
    .Y(_0140_)
  );
  \$_OR_  _0683_ (
    .A(_0140_),
    .B(_0135_),
    .Y(dbg_dout[10])
  );
  \$_AND_  _0684_ (
    .A(_0036_),
    .B(cpu_id[11]),
    .Y(_0141_)
  );
  \$_AND_  _0685_ (
    .A(_0037_),
    .B(cpu_id[27]),
    .Y(_0142_)
  );
  \$_OR_  _0686_ (
    .A(_0142_),
    .B(_0141_),
    .Y(_0143_)
  );
  \$_AND_  _0687_ (
    .A(_0035_),
    .B(mem_cnt[11]),
    .Y(_0144_)
  );
  \$_AND_  _0688_ (
    .A(_0034_),
    .B(mem_data[11]),
    .Y(_0145_)
  );
  \$_AND_  _0689_ (
    .A(_0032_),
    .B(dbg_mem_addr[11]),
    .Y(_0146_)
  );
  \$_OR_  _0690_ (
    .A(_0146_),
    .B(_0145_),
    .Y(_0147_)
  );
  \$_OR_  _0691_ (
    .A(_0147_),
    .B(_0144_),
    .Y(_0148_)
  );
  \$_OR_  _0692_ (
    .A(_0148_),
    .B(_0143_),
    .Y(dbg_dout[11])
  );
  \$_AND_  _0693_ (
    .A(_0036_),
    .B(cpu_id[12]),
    .Y(_0149_)
  );
  \$_AND_  _0694_ (
    .A(_0037_),
    .B(cpu_id[28]),
    .Y(_0150_)
  );
  \$_OR_  _0695_ (
    .A(_0150_),
    .B(_0149_),
    .Y(_0151_)
  );
  \$_AND_  _0696_ (
    .A(_0035_),
    .B(mem_cnt[12]),
    .Y(_0152_)
  );
  \$_AND_  _0697_ (
    .A(_0034_),
    .B(mem_data[12]),
    .Y(_0153_)
  );
  \$_AND_  _0698_ (
    .A(_0032_),
    .B(dbg_mem_addr[12]),
    .Y(_0154_)
  );
  \$_OR_  _0699_ (
    .A(_0154_),
    .B(_0153_),
    .Y(_0155_)
  );
  \$_OR_  _0700_ (
    .A(_0155_),
    .B(_0152_),
    .Y(_0156_)
  );
  \$_OR_  _0701_ (
    .A(_0156_),
    .B(_0151_),
    .Y(dbg_dout[12])
  );
  \$_AND_  _0702_ (
    .A(_0036_),
    .B(cpu_id[13]),
    .Y(_0157_)
  );
  \$_AND_  _0703_ (
    .A(_0037_),
    .B(cpu_id[29]),
    .Y(_0158_)
  );
  \$_OR_  _0704_ (
    .A(_0158_),
    .B(_0157_),
    .Y(_0159_)
  );
  \$_AND_  _0705_ (
    .A(_0035_),
    .B(mem_cnt[13]),
    .Y(_0160_)
  );
  \$_AND_  _0706_ (
    .A(_0034_),
    .B(mem_data[13]),
    .Y(_0161_)
  );
  \$_AND_  _0707_ (
    .A(_0032_),
    .B(dbg_mem_addr[13]),
    .Y(_0162_)
  );
  \$_OR_  _0708_ (
    .A(_0162_),
    .B(_0161_),
    .Y(_0163_)
  );
  \$_OR_  _0709_ (
    .A(_0163_),
    .B(_0160_),
    .Y(_0164_)
  );
  \$_OR_  _0710_ (
    .A(_0164_),
    .B(_0159_),
    .Y(dbg_dout[13])
  );
  \$_AND_  _0711_ (
    .A(_0036_),
    .B(cpu_id[14]),
    .Y(_0165_)
  );
  \$_AND_  _0712_ (
    .A(_0037_),
    .B(cpu_id[30]),
    .Y(_0166_)
  );
  \$_OR_  _0713_ (
    .A(_0166_),
    .B(_0165_),
    .Y(_0167_)
  );
  \$_AND_  _0714_ (
    .A(_0035_),
    .B(mem_cnt[14]),
    .Y(_0168_)
  );
  \$_AND_  _0715_ (
    .A(_0034_),
    .B(mem_data[14]),
    .Y(_0169_)
  );
  \$_AND_  _0716_ (
    .A(_0032_),
    .B(dbg_mem_addr[14]),
    .Y(_0170_)
  );
  \$_OR_  _0717_ (
    .A(_0170_),
    .B(_0169_),
    .Y(_0171_)
  );
  \$_OR_  _0718_ (
    .A(_0171_),
    .B(_0168_),
    .Y(_0172_)
  );
  \$_OR_  _0719_ (
    .A(_0172_),
    .B(_0167_),
    .Y(dbg_dout[14])
  );
  \$_AND_  _0720_ (
    .A(_0036_),
    .B(cpu_id[15]),
    .Y(_0173_)
  );
  \$_AND_  _0721_ (
    .A(_0037_),
    .B(cpu_id[31]),
    .Y(_0174_)
  );
  \$_OR_  _0722_ (
    .A(_0174_),
    .B(_0173_),
    .Y(_0175_)
  );
  \$_AND_  _0723_ (
    .A(_0035_),
    .B(mem_cnt[15]),
    .Y(_0176_)
  );
  \$_AND_  _0724_ (
    .A(_0034_),
    .B(mem_data[15]),
    .Y(_0177_)
  );
  \$_AND_  _0725_ (
    .A(_0032_),
    .B(dbg_mem_addr[15]),
    .Y(_0178_)
  );
  \$_OR_  _0726_ (
    .A(_0178_),
    .B(_0177_),
    .Y(_0179_)
  );
  \$_OR_  _0727_ (
    .A(_0179_),
    .B(_0176_),
    .Y(_0180_)
  );
  \$_OR_  _0728_ (
    .A(_0180_),
    .B(_0175_),
    .Y(dbg_dout[15])
  );
  \$_AND_  _0729_ (
    .A(_0036_),
    .B(cpu_id[1]),
    .Y(_0181_)
  );
  \$_AND_  _0730_ (
    .A(_0037_),
    .B(cpu_id[17]),
    .Y(_0182_)
  );
  \$_OR_  _0731_ (
    .A(_0182_),
    .B(_0181_),
    .Y(_0183_)
  );
  \$_AND_  _0732_ (
    .A(_0026_),
    .B(mem_ctl[1]),
    .Y(_0184_)
  );
  \$_AND_  _0733_ (
    .A(_0034_),
    .B(mem_data[1]),
    .Y(_0185_)
  );
  \$_OR_  _0734_ (
    .A(_0185_),
    .B(_0184_),
    .Y(_0186_)
  );
  \$_AND_  _0735_ (
    .A(_0032_),
    .B(dbg_mem_addr[1]),
    .Y(_0187_)
  );
  \$_AND_  _0736_ (
    .A(_0035_),
    .B(mem_cnt[1]),
    .Y(_0188_)
  );
  \$_OR_  _0737_ (
    .A(_0188_),
    .B(_0187_),
    .Y(_0189_)
  );
  \$_OR_  _0738_ (
    .A(_0189_),
    .B(_0186_),
    .Y(_0190_)
  );
  \$_OR_  _0739_ (
    .A(_0190_),
    .B(_0183_),
    .Y(dbg_dout[1])
  );
  \$_AND_  _0740_ (
    .A(_0035_),
    .B(mem_cnt[2]),
    .Y(_0191_)
  );
  \$_AND_  _0741_ (
    .A(_0034_),
    .B(mem_data[2]),
    .Y(_0192_)
  );
  \$_AND_  _0742_ (
    .A(_0032_),
    .B(dbg_mem_addr[2]),
    .Y(_0193_)
  );
  \$_OR_  _0743_ (
    .A(_0193_),
    .B(_0192_),
    .Y(_0194_)
  );
  \$_OR_  _0744_ (
    .A(_0194_),
    .B(_0191_),
    .Y(_0195_)
  );
  \$_AND_  _0745_ (
    .A(_0036_),
    .B(cpu_id[2]),
    .Y(_0196_)
  );
  \$_AND_  _0746_ (
    .A(_0037_),
    .B(cpu_id[18]),
    .Y(_0197_)
  );
  \$_OR_  _0747_ (
    .A(_0197_),
    .B(_0196_),
    .Y(_0198_)
  );
  \$_AND_  _0748_ (
    .A(_0030_),
    .B(cpu_stat[2]),
    .Y(_0199_)
  );
  \$_AND_  _0749_ (
    .A(_0026_),
    .B(mem_ctl[2]),
    .Y(_0200_)
  );
  \$_OR_  _0750_ (
    .A(_0200_),
    .B(_0199_),
    .Y(_0201_)
  );
  \$_OR_  _0751_ (
    .A(_0201_),
    .B(_0198_),
    .Y(_0202_)
  );
  \$_OR_  _0752_ (
    .A(_0202_),
    .B(_0195_),
    .Y(dbg_dout[2])
  );
  \$_AND_  _0753_ (
    .A(_0026_),
    .B(mem_bw),
    .Y(_0203_)
  );
  \$_AND_  _0754_ (
    .A(_0034_),
    .B(mem_data[3]),
    .Y(_0204_)
  );
  \$_OR_  _0755_ (
    .A(_0204_),
    .B(_0203_),
    .Y(_0205_)
  );
  \$_AND_  _0756_ (
    .A(_0032_),
    .B(dbg_mem_addr[3]),
    .Y(_0206_)
  );
  \$_AND_  _0757_ (
    .A(_0035_),
    .B(mem_cnt[3]),
    .Y(_0207_)
  );
  \$_OR_  _0758_ (
    .A(_0207_),
    .B(_0206_),
    .Y(_0208_)
  );
  \$_OR_  _0759_ (
    .A(_0208_),
    .B(_0205_),
    .Y(_0209_)
  );
  \$_AND_  _0760_ (
    .A(_0036_),
    .B(cpu_id[3]),
    .Y(_0210_)
  );
  \$_AND_  _0761_ (
    .A(_0037_),
    .B(cpu_id[19]),
    .Y(_0211_)
  );
  \$_OR_  _0762_ (
    .A(_0211_),
    .B(_0210_),
    .Y(_0212_)
  );
  \$_AND_  _0763_ (
    .A(_0038_),
    .B(cpu_ctl[3]),
    .Y(_0213_)
  );
  \$_AND_  _0764_ (
    .A(_0030_),
    .B(cpu_stat[3]),
    .Y(_0214_)
  );
  \$_OR_  _0765_ (
    .A(_0214_),
    .B(_0213_),
    .Y(_0215_)
  );
  \$_OR_  _0766_ (
    .A(_0215_),
    .B(_0212_),
    .Y(_0216_)
  );
  \$_OR_  _0767_ (
    .A(_0216_),
    .B(_0209_),
    .Y(dbg_dout[3])
  );
  \$_AND_  _0768_ (
    .A(_0036_),
    .B(cpu_id[4]),
    .Y(_0217_)
  );
  \$_AND_  _0769_ (
    .A(_0037_),
    .B(cpu_id[20]),
    .Y(_0218_)
  );
  \$_OR_  _0770_ (
    .A(_0218_),
    .B(_0217_),
    .Y(_0219_)
  );
  \$_AND_  _0771_ (
    .A(_0038_),
    .B(cpu_ctl[4]),
    .Y(_0220_)
  );
  \$_AND_  _0772_ (
    .A(_0034_),
    .B(mem_data[4]),
    .Y(_0221_)
  );
  \$_OR_  _0773_ (
    .A(_0221_),
    .B(_0220_),
    .Y(_0222_)
  );
  \$_AND_  _0774_ (
    .A(_0032_),
    .B(dbg_mem_addr[4]),
    .Y(_0223_)
  );
  \$_AND_  _0775_ (
    .A(_0035_),
    .B(mem_cnt[4]),
    .Y(_0224_)
  );
  \$_OR_  _0776_ (
    .A(_0224_),
    .B(_0223_),
    .Y(_0225_)
  );
  \$_OR_  _0777_ (
    .A(_0225_),
    .B(_0222_),
    .Y(_0226_)
  );
  \$_OR_  _0778_ (
    .A(_0226_),
    .B(_0219_),
    .Y(dbg_dout[4])
  );
  \$_AND_  _0779_ (
    .A(_0036_),
    .B(cpu_id[5]),
    .Y(_0227_)
  );
  \$_AND_  _0780_ (
    .A(_0037_),
    .B(cpu_id[21]),
    .Y(_0228_)
  );
  \$_OR_  _0781_ (
    .A(_0228_),
    .B(_0227_),
    .Y(_0229_)
  );
  \$_AND_  _0782_ (
    .A(_0038_),
    .B(cpu_ctl[5]),
    .Y(_0230_)
  );
  \$_AND_  _0783_ (
    .A(_0034_),
    .B(mem_data[5]),
    .Y(_0231_)
  );
  \$_OR_  _0784_ (
    .A(_0231_),
    .B(_0230_),
    .Y(_0232_)
  );
  \$_AND_  _0785_ (
    .A(_0032_),
    .B(dbg_mem_addr[5]),
    .Y(_0233_)
  );
  \$_AND_  _0786_ (
    .A(_0035_),
    .B(mem_cnt[5]),
    .Y(_0234_)
  );
  \$_OR_  _0787_ (
    .A(_0234_),
    .B(_0233_),
    .Y(_0235_)
  );
  \$_OR_  _0788_ (
    .A(_0235_),
    .B(_0232_),
    .Y(_0236_)
  );
  \$_OR_  _0789_ (
    .A(_0236_),
    .B(_0229_),
    .Y(dbg_dout[5])
  );
  \$_AND_  _0790_ (
    .A(_0036_),
    .B(cpu_id[6]),
    .Y(_0237_)
  );
  \$_AND_  _0791_ (
    .A(_0037_),
    .B(cpu_id[22]),
    .Y(_0238_)
  );
  \$_OR_  _0792_ (
    .A(_0238_),
    .B(_0237_),
    .Y(_0239_)
  );
  \$_AND_  _0793_ (
    .A(_0038_),
    .B(cpu_ctl[6]),
    .Y(_0240_)
  );
  \$_AND_  _0794_ (
    .A(_0034_),
    .B(mem_data[6]),
    .Y(_0241_)
  );
  \$_OR_  _0795_ (
    .A(_0241_),
    .B(_0240_),
    .Y(_0242_)
  );
  \$_AND_  _0796_ (
    .A(_0032_),
    .B(dbg_mem_addr[6]),
    .Y(_0243_)
  );
  \$_AND_  _0797_ (
    .A(_0035_),
    .B(mem_cnt[6]),
    .Y(_0244_)
  );
  \$_OR_  _0798_ (
    .A(_0244_),
    .B(_0243_),
    .Y(_0245_)
  );
  \$_OR_  _0799_ (
    .A(_0245_),
    .B(_0242_),
    .Y(_0246_)
  );
  \$_OR_  _0800_ (
    .A(_0246_),
    .B(_0239_),
    .Y(dbg_dout[6])
  );
  \$_AND_  _0801_ (
    .A(_0036_),
    .B(cpu_id[7]),
    .Y(_0247_)
  );
  \$_AND_  _0802_ (
    .A(_0037_),
    .B(cpu_id[23]),
    .Y(_0248_)
  );
  \$_OR_  _0803_ (
    .A(_0248_),
    .B(_0247_),
    .Y(_0249_)
  );
  \$_AND_  _0804_ (
    .A(_0035_),
    .B(mem_cnt[7]),
    .Y(_0250_)
  );
  \$_AND_  _0805_ (
    .A(_0034_),
    .B(mem_data[7]),
    .Y(_0251_)
  );
  \$_AND_  _0806_ (
    .A(_0032_),
    .B(dbg_mem_addr[7]),
    .Y(_0252_)
  );
  \$_OR_  _0807_ (
    .A(_0252_),
    .B(_0251_),
    .Y(_0253_)
  );
  \$_OR_  _0808_ (
    .A(_0253_),
    .B(_0250_),
    .Y(_0254_)
  );
  \$_OR_  _0809_ (
    .A(_0254_),
    .B(_0249_),
    .Y(dbg_dout[7])
  );
  \$_AND_  _0810_ (
    .A(_0036_),
    .B(cpu_id[8]),
    .Y(_0255_)
  );
  \$_AND_  _0811_ (
    .A(_0037_),
    .B(cpu_id[24]),
    .Y(_0256_)
  );
  \$_OR_  _0812_ (
    .A(_0256_),
    .B(_0255_),
    .Y(_0257_)
  );
  \$_AND_  _0813_ (
    .A(_0035_),
    .B(mem_cnt[8]),
    .Y(_0258_)
  );
  \$_AND_  _0814_ (
    .A(_0034_),
    .B(mem_data[8]),
    .Y(_0259_)
  );
  \$_AND_  _0815_ (
    .A(_0032_),
    .B(dbg_mem_addr[8]),
    .Y(_0260_)
  );
  \$_OR_  _0816_ (
    .A(_0260_),
    .B(_0259_),
    .Y(_0261_)
  );
  \$_OR_  _0817_ (
    .A(_0261_),
    .B(_0258_),
    .Y(_0262_)
  );
  \$_OR_  _0818_ (
    .A(_0262_),
    .B(_0257_),
    .Y(dbg_dout[8])
  );
  \$_AND_  _0819_ (
    .A(_0036_),
    .B(cpu_id[9]),
    .Y(_0263_)
  );
  \$_AND_  _0820_ (
    .A(_0037_),
    .B(cpu_id[25]),
    .Y(_0264_)
  );
  \$_OR_  _0821_ (
    .A(_0264_),
    .B(_0263_),
    .Y(_0265_)
  );
  \$_AND_  _0822_ (
    .A(_0035_),
    .B(mem_cnt[9]),
    .Y(_0266_)
  );
  \$_AND_  _0823_ (
    .A(_0034_),
    .B(mem_data[9]),
    .Y(_0267_)
  );
  \$_AND_  _0824_ (
    .A(_0032_),
    .B(dbg_mem_addr[9]),
    .Y(_0268_)
  );
  \$_OR_  _0825_ (
    .A(_0268_),
    .B(_0267_),
    .Y(_0269_)
  );
  \$_OR_  _0826_ (
    .A(_0269_),
    .B(_0266_),
    .Y(_0270_)
  );
  \$_OR_  _0827_ (
    .A(_0270_),
    .B(_0265_),
    .Y(dbg_dout[9])
  );
  \$_OR_  _0828_ (
    .A(dbg_rd),
    .B(dbg_wr),
    .Y(_0271_)
  );
  \$_AND_  _0829_ (
    .A(_0271_),
    .B(mem_burst),
    .Y(_0272_)
  );
  \$_OR_  _0830_ (
    .A(_0272_),
    .B(mem_burst_rd),
    .Y(_0011_)
  );
  \$_MUX_  _0831_ (
    .A(cpu_ctl[3]),
    .B(dbg_din[3]),
    .S(_0043_),
    .Y(_0000_[0])
  );
  \$_MUX_  _0832_ (
    .A(cpu_ctl[4]),
    .B(dbg_din[4]),
    .S(_0043_),
    .Y(_0000_[1])
  );
  \$_MUX_  _0833_ (
    .A(cpu_ctl[5]),
    .B(dbg_din[5]),
    .S(_0043_),
    .Y(_0000_[2])
  );
  \$_MUX_  _0834_ (
    .A(cpu_ctl[6]),
    .B(dbg_din[6]),
    .S(_0043_),
    .Y(_0000_[3])
  );
  \$_INV_  _0835_ (
    .A(_0030_),
    .Y(_0273_)
  );
  \$_OR_  _0836_ (
    .A(_0273_),
    .B(_0109_),
    .Y(_0274_)
  );
  \$_OR_  _0837_ (
    .A(puc_pnd_set),
    .B(cpu_stat[2]),
    .Y(_0275_)
  );
  \$_INV_  _0838_ (
    .A(dbg_din[2]),
    .Y(_0276_)
  );
  \$_AND_  _0839_ (
    .A(cpu_stat[2]),
    .B(_0276_),
    .Y(_0277_)
  );
  \$_OR_  _0840_ (
    .A(_0277_),
    .B(puc_pnd_set),
    .Y(_0278_)
  );
  \$_MUX_  _0841_ (
    .A(_0278_),
    .B(_0275_),
    .S(_0274_),
    .Y(_0001_[0])
  );
  \$_OR_  _0842_ (
    .A(_0104_),
    .B(cpu_stat[3]),
    .Y(_0279_)
  );
  \$_INV_  _0843_ (
    .A(dbg_din[3]),
    .Y(_0280_)
  );
  \$_AND_  _0844_ (
    .A(_0280_),
    .B(cpu_stat[3]),
    .Y(_0281_)
  );
  \$_OR_  _0845_ (
    .A(_0281_),
    .B(_0104_),
    .Y(_0282_)
  );
  \$_MUX_  _0846_ (
    .A(_0282_),
    .B(_0279_),
    .S(_0274_),
    .Y(_0001_[1])
  );
  \$_MUX_  _0847_ (
    .A(mem_ctl[1]),
    .B(dbg_din[1]),
    .S(_0039_),
    .Y(_0008_[0])
  );
  \$_MUX_  _0848_ (
    .A(mem_ctl[2]),
    .B(dbg_din[2]),
    .S(_0039_),
    .Y(_0008_[1])
  );
  \$_MUX_  _0849_ (
    .A(mem_bw),
    .B(dbg_din[3]),
    .S(_0039_),
    .Y(_0008_[2])
  );
  \$_AND_  _0850_ (
    .A(_0034_),
    .B(dbg_wr),
    .Y(_0283_)
  );
  \$_AND_  _0851_ (
    .A(_0113_),
    .B(mem_ctl[2]),
    .Y(_0284_)
  );
  \$_AND_  _0852_ (
    .A(_0284_),
    .B(_0115_),
    .Y(_0285_)
  );
  \$_INV_  _0853_ (
    .A(dbg_mem_rd_dly),
    .Y(_0286_)
  );
  \$_MUX_  _0854_ (
    .A(dbg_mem_din[0]),
    .B(dbg_mem_din[8]),
    .S(dbg_mem_addr[0]),
    .Y(_0287_)
  );
  \$_MUX_  _0855_ (
    .A(_0287_),
    .B(dbg_mem_din[0]),
    .S(_0120_),
    .Y(_0288_)
  );
  \$_MUX_  _0856_ (
    .A(_0288_),
    .B(mem_data[0]),
    .S(_0286_),
    .Y(_0289_)
  );
  \$_MUX_  _0857_ (
    .A(_0289_),
    .B(dbg_reg_din[0]),
    .S(_0285_),
    .Y(_0290_)
  );
  \$_MUX_  _0858_ (
    .A(_0290_),
    .B(dbg_din[0]),
    .S(_0283_),
    .Y(_0009_[0])
  );
  \$_AND_  _0859_ (
    .A(_0286_),
    .B(mem_data[10]),
    .Y(_0291_)
  );
  \$_AND_  _0860_ (
    .A(dbg_mem_rd_dly),
    .B(_0120_),
    .Y(_0292_)
  );
  \$_AND_  _0861_ (
    .A(_0292_),
    .B(dbg_mem_din[10]),
    .Y(_0293_)
  );
  \$_OR_  _0862_ (
    .A(_0293_),
    .B(_0291_),
    .Y(_0294_)
  );
  \$_MUX_  _0863_ (
    .A(_0294_),
    .B(dbg_reg_din[10]),
    .S(_0285_),
    .Y(_0295_)
  );
  \$_MUX_  _0864_ (
    .A(_0295_),
    .B(dbg_din[10]),
    .S(_0283_),
    .Y(_0009_[10])
  );
  \$_AND_  _0865_ (
    .A(_0286_),
    .B(mem_data[11]),
    .Y(_0296_)
  );
  \$_AND_  _0866_ (
    .A(_0292_),
    .B(dbg_mem_din[11]),
    .Y(_0297_)
  );
  \$_OR_  _0867_ (
    .A(_0297_),
    .B(_0296_),
    .Y(_0298_)
  );
  \$_MUX_  _0868_ (
    .A(_0298_),
    .B(dbg_reg_din[11]),
    .S(_0285_),
    .Y(_0299_)
  );
  \$_MUX_  _0869_ (
    .A(_0299_),
    .B(dbg_din[11]),
    .S(_0283_),
    .Y(_0009_[11])
  );
  \$_AND_  _0870_ (
    .A(_0286_),
    .B(mem_data[12]),
    .Y(_0300_)
  );
  \$_AND_  _0871_ (
    .A(_0292_),
    .B(dbg_mem_din[12]),
    .Y(_0301_)
  );
  \$_OR_  _0872_ (
    .A(_0301_),
    .B(_0300_),
    .Y(_0302_)
  );
  \$_MUX_  _0873_ (
    .A(_0302_),
    .B(dbg_reg_din[12]),
    .S(_0285_),
    .Y(_0303_)
  );
  \$_MUX_  _0874_ (
    .A(_0303_),
    .B(dbg_din[12]),
    .S(_0283_),
    .Y(_0009_[12])
  );
  \$_AND_  _0875_ (
    .A(_0286_),
    .B(mem_data[13]),
    .Y(_0304_)
  );
  \$_AND_  _0876_ (
    .A(_0292_),
    .B(dbg_mem_din[13]),
    .Y(_0305_)
  );
  \$_OR_  _0877_ (
    .A(_0305_),
    .B(_0304_),
    .Y(_0306_)
  );
  \$_MUX_  _0878_ (
    .A(_0306_),
    .B(dbg_reg_din[13]),
    .S(_0285_),
    .Y(_0307_)
  );
  \$_MUX_  _0879_ (
    .A(_0307_),
    .B(dbg_din[13]),
    .S(_0283_),
    .Y(_0009_[13])
  );
  \$_AND_  _0880_ (
    .A(_0286_),
    .B(mem_data[14]),
    .Y(_0308_)
  );
  \$_AND_  _0881_ (
    .A(_0292_),
    .B(dbg_mem_din[14]),
    .Y(_0309_)
  );
  \$_OR_  _0882_ (
    .A(_0309_),
    .B(_0308_),
    .Y(_0310_)
  );
  \$_MUX_  _0883_ (
    .A(_0310_),
    .B(dbg_reg_din[14]),
    .S(_0285_),
    .Y(_0311_)
  );
  \$_MUX_  _0884_ (
    .A(_0311_),
    .B(dbg_din[14]),
    .S(_0283_),
    .Y(_0009_[14])
  );
  \$_AND_  _0885_ (
    .A(_0286_),
    .B(mem_data[15]),
    .Y(_0312_)
  );
  \$_AND_  _0886_ (
    .A(_0292_),
    .B(dbg_mem_din[15]),
    .Y(_0313_)
  );
  \$_OR_  _0887_ (
    .A(_0313_),
    .B(_0312_),
    .Y(_0314_)
  );
  \$_MUX_  _0888_ (
    .A(_0314_),
    .B(dbg_reg_din[15]),
    .S(_0285_),
    .Y(_0315_)
  );
  \$_MUX_  _0889_ (
    .A(_0315_),
    .B(dbg_din[15]),
    .S(_0283_),
    .Y(_0009_[15])
  );
  \$_MUX_  _0890_ (
    .A(dbg_mem_din[1]),
    .B(dbg_mem_din[9]),
    .S(dbg_mem_addr[0]),
    .Y(_0316_)
  );
  \$_MUX_  _0891_ (
    .A(_0316_),
    .B(dbg_mem_din[1]),
    .S(_0120_),
    .Y(_0317_)
  );
  \$_MUX_  _0892_ (
    .A(_0317_),
    .B(mem_data[1]),
    .S(_0286_),
    .Y(_0318_)
  );
  \$_MUX_  _0893_ (
    .A(_0318_),
    .B(dbg_reg_din[1]),
    .S(_0285_),
    .Y(_0319_)
  );
  \$_MUX_  _0894_ (
    .A(_0319_),
    .B(dbg_din[1]),
    .S(_0283_),
    .Y(_0009_[1])
  );
  \$_MUX_  _0895_ (
    .A(dbg_mem_din[2]),
    .B(dbg_mem_din[10]),
    .S(dbg_mem_addr[0]),
    .Y(_0320_)
  );
  \$_MUX_  _0896_ (
    .A(_0320_),
    .B(dbg_mem_din[2]),
    .S(_0120_),
    .Y(_0321_)
  );
  \$_MUX_  _0897_ (
    .A(_0321_),
    .B(mem_data[2]),
    .S(_0286_),
    .Y(_0322_)
  );
  \$_MUX_  _0898_ (
    .A(_0322_),
    .B(dbg_reg_din[2]),
    .S(_0285_),
    .Y(_0323_)
  );
  \$_MUX_  _0899_ (
    .A(_0323_),
    .B(dbg_din[2]),
    .S(_0283_),
    .Y(_0009_[2])
  );
  \$_MUX_  _0900_ (
    .A(dbg_mem_din[3]),
    .B(dbg_mem_din[11]),
    .S(dbg_mem_addr[0]),
    .Y(_0324_)
  );
  \$_MUX_  _0901_ (
    .A(_0324_),
    .B(dbg_mem_din[3]),
    .S(_0120_),
    .Y(_0325_)
  );
  \$_MUX_  _0902_ (
    .A(_0325_),
    .B(mem_data[3]),
    .S(_0286_),
    .Y(_0326_)
  );
  \$_MUX_  _0903_ (
    .A(_0326_),
    .B(dbg_reg_din[3]),
    .S(_0285_),
    .Y(_0327_)
  );
  \$_MUX_  _0904_ (
    .A(_0327_),
    .B(dbg_din[3]),
    .S(_0283_),
    .Y(_0009_[3])
  );
  \$_MUX_  _0905_ (
    .A(dbg_mem_din[4]),
    .B(dbg_mem_din[12]),
    .S(dbg_mem_addr[0]),
    .Y(_0328_)
  );
  \$_MUX_  _0906_ (
    .A(_0328_),
    .B(dbg_mem_din[4]),
    .S(_0120_),
    .Y(_0329_)
  );
  \$_MUX_  _0907_ (
    .A(_0329_),
    .B(mem_data[4]),
    .S(_0286_),
    .Y(_0330_)
  );
  \$_MUX_  _0908_ (
    .A(_0330_),
    .B(dbg_reg_din[4]),
    .S(_0285_),
    .Y(_0331_)
  );
  \$_MUX_  _0909_ (
    .A(_0331_),
    .B(dbg_din[4]),
    .S(_0283_),
    .Y(_0009_[4])
  );
  \$_MUX_  _0910_ (
    .A(dbg_mem_din[5]),
    .B(dbg_mem_din[13]),
    .S(dbg_mem_addr[0]),
    .Y(_0332_)
  );
  \$_MUX_  _0911_ (
    .A(_0332_),
    .B(dbg_mem_din[5]),
    .S(_0120_),
    .Y(_0333_)
  );
  \$_MUX_  _0912_ (
    .A(_0333_),
    .B(mem_data[5]),
    .S(_0286_),
    .Y(_0334_)
  );
  \$_MUX_  _0913_ (
    .A(_0334_),
    .B(dbg_reg_din[5]),
    .S(_0285_),
    .Y(_0335_)
  );
  \$_MUX_  _0914_ (
    .A(_0335_),
    .B(dbg_din[5]),
    .S(_0283_),
    .Y(_0009_[5])
  );
  \$_MUX_  _0915_ (
    .A(dbg_mem_din[6]),
    .B(dbg_mem_din[14]),
    .S(dbg_mem_addr[0]),
    .Y(_0336_)
  );
  \$_MUX_  _0916_ (
    .A(_0336_),
    .B(dbg_mem_din[6]),
    .S(_0120_),
    .Y(_0337_)
  );
  \$_MUX_  _0917_ (
    .A(_0337_),
    .B(mem_data[6]),
    .S(_0286_),
    .Y(_0338_)
  );
  \$_MUX_  _0918_ (
    .A(_0338_),
    .B(dbg_reg_din[6]),
    .S(_0285_),
    .Y(_0339_)
  );
  \$_MUX_  _0919_ (
    .A(_0339_),
    .B(dbg_din[6]),
    .S(_0283_),
    .Y(_0009_[6])
  );
  \$_MUX_  _0920_ (
    .A(dbg_mem_din[7]),
    .B(dbg_mem_din[15]),
    .S(dbg_mem_addr[0]),
    .Y(_0340_)
  );
  \$_MUX_  _0921_ (
    .A(_0340_),
    .B(dbg_mem_din[7]),
    .S(_0120_),
    .Y(_0341_)
  );
  \$_MUX_  _0922_ (
    .A(_0341_),
    .B(mem_data[7]),
    .S(_0286_),
    .Y(_0342_)
  );
  \$_MUX_  _0923_ (
    .A(_0342_),
    .B(dbg_reg_din[7]),
    .S(_0285_),
    .Y(_0343_)
  );
  \$_MUX_  _0924_ (
    .A(_0343_),
    .B(dbg_din[7]),
    .S(_0283_),
    .Y(_0009_[7])
  );
  \$_AND_  _0925_ (
    .A(_0286_),
    .B(mem_data[8]),
    .Y(_0344_)
  );
  \$_AND_  _0926_ (
    .A(_0292_),
    .B(dbg_mem_din[8]),
    .Y(_0345_)
  );
  \$_OR_  _0927_ (
    .A(_0345_),
    .B(_0344_),
    .Y(_0346_)
  );
  \$_MUX_  _0928_ (
    .A(_0346_),
    .B(dbg_reg_din[8]),
    .S(_0285_),
    .Y(_0347_)
  );
  \$_MUX_  _0929_ (
    .A(_0347_),
    .B(dbg_din[8]),
    .S(_0283_),
    .Y(_0009_[8])
  );
  \$_AND_  _0930_ (
    .A(_0286_),
    .B(mem_data[9]),
    .Y(_0348_)
  );
  \$_AND_  _0931_ (
    .A(_0292_),
    .B(dbg_mem_din[9]),
    .Y(_0349_)
  );
  \$_OR_  _0932_ (
    .A(_0349_),
    .B(_0348_),
    .Y(_0350_)
  );
  \$_MUX_  _0933_ (
    .A(_0350_),
    .B(dbg_reg_din[9]),
    .S(_0285_),
    .Y(_0351_)
  );
  \$_MUX_  _0934_ (
    .A(_0351_),
    .B(dbg_din[9]),
    .S(_0283_),
    .Y(_0009_[9])
  );
  \$_AND_  _0935_ (
    .A(_0032_),
    .B(dbg_wr),
    .Y(_0352_)
  );
  \$_AND_  _0936_ (
    .A(_0117_),
    .B(dbg_rd_rdy),
    .Y(_0353_)
  );
  \$_OR_  _0937_ (
    .A(_0353_),
    .B(dbg_mem_wr[0]),
    .Y(_0354_)
  );
  \$_OR_  _0938_ (
    .A(_0354_),
    .B(dbg_mem_wr[1]),
    .Y(_0355_)
  );
  \$_AND_  _0939_ (
    .A(mem_ctl[2]),
    .B(dbg_rd_rdy),
    .Y(_0356_)
  );
  \$_OR_  _0940_ (
    .A(_0356_),
    .B(dbg_reg_wr),
    .Y(_0357_)
  );
  \$_OR_  _0941_ (
    .A(_0357_),
    .B(_0355_),
    .Y(_0358_)
  );
  \$_INV_  _0942_ (
    .A(_0358_),
    .Y(_0359_)
  );
  \$_AND_  _0943_ (
    .A(_0355_),
    .B(_0120_),
    .Y(_0360_)
  );
  \$_OR_  _0944_ (
    .A(_0360_),
    .B(_0062_),
    .Y(_0361_)
  );
  \$_OR_  _0945_ (
    .A(_0361_),
    .B(_0359_),
    .Y(_0362_)
  );
  \$_XOR_  _0946_ (
    .A(_0362_),
    .B(_0119_),
    .Y(_0363_)
  );
  \$_MUX_  _0947_ (
    .A(_0363_),
    .B(dbg_din[0]),
    .S(_0352_),
    .Y(_0005_[0])
  );
  \$_INV_  _0948_ (
    .A(dbg_mem_addr[10]),
    .Y(_0364_)
  );
  \$_INV_  _0949_ (
    .A(dbg_mem_addr[9]),
    .Y(_0365_)
  );
  \$_INV_  _0950_ (
    .A(dbg_mem_addr[8]),
    .Y(_0366_)
  );
  \$_INV_  _0951_ (
    .A(dbg_mem_addr[7]),
    .Y(_0367_)
  );
  \$_INV_  _0952_ (
    .A(dbg_mem_addr[6]),
    .Y(_0368_)
  );
  \$_INV_  _0953_ (
    .A(dbg_mem_addr[5]),
    .Y(_0369_)
  );
  \$_INV_  _0954_ (
    .A(dbg_mem_addr[4]),
    .Y(_0370_)
  );
  \$_INV_  _0955_ (
    .A(dbg_mem_addr[3]),
    .Y(_0371_)
  );
  \$_INV_  _0956_ (
    .A(dbg_mem_addr[2]),
    .Y(_0372_)
  );
  \$_INV_  _0957_ (
    .A(dbg_mem_addr[1]),
    .Y(_0373_)
  );
  \$_AND_  _0958_ (
    .A(_0360_),
    .B(_0061_),
    .Y(_0374_)
  );
  \$_INV_  _0959_ (
    .A(_0374_),
    .Y(_0375_)
  );
  \$_OR_  _0960_ (
    .A(_0375_),
    .B(_0373_),
    .Y(_0376_)
  );
  \$_XOR_  _0961_ (
    .A(_0374_),
    .B(_0373_),
    .Y(_0377_)
  );
  \$_OR_  _0962_ (
    .A(_0362_),
    .B(_0119_),
    .Y(_0378_)
  );
  \$_OR_  _0963_ (
    .A(_0378_),
    .B(_0377_),
    .Y(_0379_)
  );
  \$_AND_  _0964_ (
    .A(_0379_),
    .B(_0376_),
    .Y(_0380_)
  );
  \$_OR_  _0965_ (
    .A(_0380_),
    .B(_0372_),
    .Y(_0381_)
  );
  \$_OR_  _0966_ (
    .A(_0381_),
    .B(_0371_),
    .Y(_0382_)
  );
  \$_OR_  _0967_ (
    .A(_0382_),
    .B(_0370_),
    .Y(_0383_)
  );
  \$_OR_  _0968_ (
    .A(_0383_),
    .B(_0369_),
    .Y(_0384_)
  );
  \$_OR_  _0969_ (
    .A(_0384_),
    .B(_0368_),
    .Y(_0385_)
  );
  \$_OR_  _0970_ (
    .A(_0385_),
    .B(_0367_),
    .Y(_0386_)
  );
  \$_OR_  _0971_ (
    .A(_0386_),
    .B(_0366_),
    .Y(_0387_)
  );
  \$_OR_  _0972_ (
    .A(_0387_),
    .B(_0365_),
    .Y(_0388_)
  );
  \$_XOR_  _0973_ (
    .A(_0388_),
    .B(_0364_),
    .Y(_0389_)
  );
  \$_MUX_  _0974_ (
    .A(_0389_),
    .B(dbg_din[10]),
    .S(_0352_),
    .Y(_0005_[10])
  );
  \$_INV_  _0975_ (
    .A(dbg_mem_addr[11]),
    .Y(_0390_)
  );
  \$_OR_  _0976_ (
    .A(_0388_),
    .B(_0364_),
    .Y(_0391_)
  );
  \$_XOR_  _0977_ (
    .A(_0391_),
    .B(_0390_),
    .Y(_0392_)
  );
  \$_MUX_  _0978_ (
    .A(_0392_),
    .B(dbg_din[11]),
    .S(_0352_),
    .Y(_0005_[11])
  );
  \$_INV_  _0979_ (
    .A(dbg_mem_addr[12]),
    .Y(_0393_)
  );
  \$_OR_  _0980_ (
    .A(_0391_),
    .B(_0390_),
    .Y(_0394_)
  );
  \$_XOR_  _0981_ (
    .A(_0394_),
    .B(_0393_),
    .Y(_0395_)
  );
  \$_MUX_  _0982_ (
    .A(_0395_),
    .B(dbg_din[12]),
    .S(_0352_),
    .Y(_0005_[12])
  );
  \$_INV_  _0983_ (
    .A(dbg_mem_addr[13]),
    .Y(_0396_)
  );
  \$_OR_  _0984_ (
    .A(_0394_),
    .B(_0393_),
    .Y(_0397_)
  );
  \$_XOR_  _0985_ (
    .A(_0397_),
    .B(_0396_),
    .Y(_0398_)
  );
  \$_MUX_  _0986_ (
    .A(_0398_),
    .B(dbg_din[13]),
    .S(_0352_),
    .Y(_0005_[13])
  );
  \$_INV_  _0987_ (
    .A(dbg_mem_addr[14]),
    .Y(_0399_)
  );
  \$_OR_  _0988_ (
    .A(_0397_),
    .B(_0396_),
    .Y(_0400_)
  );
  \$_XOR_  _0989_ (
    .A(_0400_),
    .B(_0399_),
    .Y(_0401_)
  );
  \$_MUX_  _0990_ (
    .A(_0401_),
    .B(dbg_din[14]),
    .S(_0352_),
    .Y(_0005_[14])
  );
  \$_INV_  _0991_ (
    .A(dbg_mem_addr[15]),
    .Y(_0402_)
  );
  \$_OR_  _0992_ (
    .A(_0400_),
    .B(_0399_),
    .Y(_0403_)
  );
  \$_XOR_  _0993_ (
    .A(_0403_),
    .B(_0402_),
    .Y(_0404_)
  );
  \$_MUX_  _0994_ (
    .A(_0404_),
    .B(dbg_din[15]),
    .S(_0352_),
    .Y(_0005_[15])
  );
  \$_XOR_  _0995_ (
    .A(_0378_),
    .B(_0377_),
    .Y(_0405_)
  );
  \$_MUX_  _0996_ (
    .A(_0405_),
    .B(dbg_din[1]),
    .S(_0352_),
    .Y(_0005_[1])
  );
  \$_XOR_  _0997_ (
    .A(_0380_),
    .B(_0372_),
    .Y(_0406_)
  );
  \$_MUX_  _0998_ (
    .A(_0406_),
    .B(dbg_din[2]),
    .S(_0352_),
    .Y(_0005_[2])
  );
  \$_XOR_  _0999_ (
    .A(_0381_),
    .B(_0371_),
    .Y(_0407_)
  );
  \$_MUX_  _1000_ (
    .A(_0407_),
    .B(dbg_din[3]),
    .S(_0352_),
    .Y(_0005_[3])
  );
  \$_XOR_  _1001_ (
    .A(_0382_),
    .B(_0370_),
    .Y(_0408_)
  );
  \$_MUX_  _1002_ (
    .A(_0408_),
    .B(dbg_din[4]),
    .S(_0352_),
    .Y(_0005_[4])
  );
  \$_XOR_  _1003_ (
    .A(_0383_),
    .B(_0369_),
    .Y(_0409_)
  );
  \$_MUX_  _1004_ (
    .A(_0409_),
    .B(dbg_din[5]),
    .S(_0352_),
    .Y(_0005_[5])
  );
  \$_XOR_  _1005_ (
    .A(_0384_),
    .B(_0368_),
    .Y(_0410_)
  );
  \$_MUX_  _1006_ (
    .A(_0410_),
    .B(dbg_din[6]),
    .S(_0352_),
    .Y(_0005_[6])
  );
  \$_XOR_  _1007_ (
    .A(_0385_),
    .B(_0367_),
    .Y(_0411_)
  );
  \$_MUX_  _1008_ (
    .A(_0411_),
    .B(dbg_din[7]),
    .S(_0352_),
    .Y(_0005_[7])
  );
  \$_XOR_  _1009_ (
    .A(_0386_),
    .B(_0366_),
    .Y(_0412_)
  );
  \$_MUX_  _1010_ (
    .A(_0412_),
    .B(dbg_din[8]),
    .S(_0352_),
    .Y(_0005_[8])
  );
  \$_XOR_  _1011_ (
    .A(_0387_),
    .B(_0365_),
    .Y(_0413_)
  );
  \$_MUX_  _1012_ (
    .A(_0413_),
    .B(dbg_din[9]),
    .S(_0352_),
    .Y(_0005_[9])
  );
  \$_AND_  _1013_ (
    .A(_0035_),
    .B(dbg_wr),
    .Y(_0414_)
  );
  \$_AND_  _1014_ (
    .A(_0061_),
    .B(mem_burst),
    .Y(_0415_)
  );
  \$_AND_  _1015_ (
    .A(_0415_),
    .B(_0358_),
    .Y(_0416_)
  );
  \$_XOR_  _1016_ (
    .A(_0416_),
    .B(mem_cnt[0]),
    .Y(_0417_)
  );
  \$_MUX_  _1017_ (
    .A(_0417_),
    .B(dbg_din[0]),
    .S(_0414_),
    .Y(_0007_[0])
  );
  \$_XOR_  _1018_ (
    .A(_0416_),
    .B(mem_cnt[10]),
    .Y(_0418_)
  );
  \$_AND_  _1019_ (
    .A(_0416_),
    .B(mem_cnt[9]),
    .Y(_0419_)
  );
  \$_XOR_  _1020_ (
    .A(_0416_),
    .B(mem_cnt[9]),
    .Y(_0420_)
  );
  \$_AND_  _1021_ (
    .A(_0416_),
    .B(mem_cnt[8]),
    .Y(_0421_)
  );
  \$_XOR_  _1022_ (
    .A(_0416_),
    .B(mem_cnt[8]),
    .Y(_0422_)
  );
  \$_AND_  _1023_ (
    .A(_0416_),
    .B(mem_cnt[7]),
    .Y(_0423_)
  );
  \$_XOR_  _1024_ (
    .A(_0416_),
    .B(mem_cnt[7]),
    .Y(_0424_)
  );
  \$_AND_  _1025_ (
    .A(_0416_),
    .B(mem_cnt[6]),
    .Y(_0425_)
  );
  \$_XOR_  _1026_ (
    .A(_0416_),
    .B(mem_cnt[6]),
    .Y(_0426_)
  );
  \$_AND_  _1027_ (
    .A(_0416_),
    .B(mem_cnt[5]),
    .Y(_0427_)
  );
  \$_XOR_  _1028_ (
    .A(_0416_),
    .B(mem_cnt[5]),
    .Y(_0428_)
  );
  \$_AND_  _1029_ (
    .A(_0416_),
    .B(mem_cnt[4]),
    .Y(_0429_)
  );
  \$_XOR_  _1030_ (
    .A(_0416_),
    .B(mem_cnt[4]),
    .Y(_0430_)
  );
  \$_AND_  _1031_ (
    .A(_0416_),
    .B(mem_cnt[3]),
    .Y(_0431_)
  );
  \$_XOR_  _1032_ (
    .A(_0416_),
    .B(mem_cnt[3]),
    .Y(_0432_)
  );
  \$_AND_  _1033_ (
    .A(_0416_),
    .B(mem_cnt[2]),
    .Y(_0433_)
  );
  \$_XOR_  _1034_ (
    .A(_0416_),
    .B(mem_cnt[2]),
    .Y(_0434_)
  );
  \$_AND_  _1035_ (
    .A(_0416_),
    .B(mem_cnt[1]),
    .Y(_0435_)
  );
  \$_XOR_  _1036_ (
    .A(_0416_),
    .B(mem_cnt[1]),
    .Y(_0436_)
  );
  \$_AND_  _1037_ (
    .A(_0416_),
    .B(mem_cnt[0]),
    .Y(_0437_)
  );
  \$_AND_  _1038_ (
    .A(_0437_),
    .B(_0436_),
    .Y(_0438_)
  );
  \$_OR_  _1039_ (
    .A(_0438_),
    .B(_0435_),
    .Y(_0439_)
  );
  \$_AND_  _1040_ (
    .A(_0439_),
    .B(_0434_),
    .Y(_0440_)
  );
  \$_OR_  _1041_ (
    .A(_0440_),
    .B(_0433_),
    .Y(_0441_)
  );
  \$_AND_  _1042_ (
    .A(_0441_),
    .B(_0432_),
    .Y(_0442_)
  );
  \$_OR_  _1043_ (
    .A(_0442_),
    .B(_0431_),
    .Y(_0443_)
  );
  \$_AND_  _1044_ (
    .A(_0443_),
    .B(_0430_),
    .Y(_0444_)
  );
  \$_OR_  _1045_ (
    .A(_0444_),
    .B(_0429_),
    .Y(_0445_)
  );
  \$_AND_  _1046_ (
    .A(_0445_),
    .B(_0428_),
    .Y(_0446_)
  );
  \$_OR_  _1047_ (
    .A(_0446_),
    .B(_0427_),
    .Y(_0447_)
  );
  \$_AND_  _1048_ (
    .A(_0447_),
    .B(_0426_),
    .Y(_0448_)
  );
  \$_OR_  _1049_ (
    .A(_0448_),
    .B(_0425_),
    .Y(_0449_)
  );
  \$_AND_  _1050_ (
    .A(_0449_),
    .B(_0424_),
    .Y(_0450_)
  );
  \$_OR_  _1051_ (
    .A(_0450_),
    .B(_0423_),
    .Y(_0451_)
  );
  \$_AND_  _1052_ (
    .A(_0451_),
    .B(_0422_),
    .Y(_0452_)
  );
  \$_OR_  _1053_ (
    .A(_0452_),
    .B(_0421_),
    .Y(_0453_)
  );
  \$_AND_  _1054_ (
    .A(_0453_),
    .B(_0420_),
    .Y(_0454_)
  );
  \$_OR_  _1055_ (
    .A(_0454_),
    .B(_0419_),
    .Y(_0455_)
  );
  \$_XOR_  _1056_ (
    .A(_0455_),
    .B(_0418_),
    .Y(_0456_)
  );
  \$_MUX_  _1057_ (
    .A(_0456_),
    .B(dbg_din[10]),
    .S(_0414_),
    .Y(_0007_[10])
  );
  \$_XOR_  _1058_ (
    .A(_0416_),
    .B(mem_cnt[11]),
    .Y(_0457_)
  );
  \$_AND_  _1059_ (
    .A(_0416_),
    .B(mem_cnt[10]),
    .Y(_0458_)
  );
  \$_AND_  _1060_ (
    .A(_0455_),
    .B(_0418_),
    .Y(_0459_)
  );
  \$_OR_  _1061_ (
    .A(_0459_),
    .B(_0458_),
    .Y(_0460_)
  );
  \$_XOR_  _1062_ (
    .A(_0460_),
    .B(_0457_),
    .Y(_0461_)
  );
  \$_MUX_  _1063_ (
    .A(_0461_),
    .B(dbg_din[11]),
    .S(_0414_),
    .Y(_0007_[11])
  );
  \$_XOR_  _1064_ (
    .A(_0416_),
    .B(mem_cnt[12]),
    .Y(_0462_)
  );
  \$_AND_  _1065_ (
    .A(_0416_),
    .B(mem_cnt[11]),
    .Y(_0463_)
  );
  \$_AND_  _1066_ (
    .A(_0460_),
    .B(_0457_),
    .Y(_0464_)
  );
  \$_OR_  _1067_ (
    .A(_0464_),
    .B(_0463_),
    .Y(_0465_)
  );
  \$_XOR_  _1068_ (
    .A(_0465_),
    .B(_0462_),
    .Y(_0466_)
  );
  \$_MUX_  _1069_ (
    .A(_0466_),
    .B(dbg_din[12]),
    .S(_0414_),
    .Y(_0007_[12])
  );
  \$_XOR_  _1070_ (
    .A(_0416_),
    .B(mem_cnt[13]),
    .Y(_0467_)
  );
  \$_AND_  _1071_ (
    .A(_0416_),
    .B(mem_cnt[12]),
    .Y(_0468_)
  );
  \$_AND_  _1072_ (
    .A(_0465_),
    .B(_0462_),
    .Y(_0469_)
  );
  \$_OR_  _1073_ (
    .A(_0469_),
    .B(_0468_),
    .Y(_0470_)
  );
  \$_XOR_  _1074_ (
    .A(_0470_),
    .B(_0467_),
    .Y(_0471_)
  );
  \$_MUX_  _1075_ (
    .A(_0471_),
    .B(dbg_din[13]),
    .S(_0414_),
    .Y(_0007_[13])
  );
  \$_XOR_  _1076_ (
    .A(_0416_),
    .B(mem_cnt[14]),
    .Y(_0472_)
  );
  \$_AND_  _1077_ (
    .A(_0416_),
    .B(mem_cnt[13]),
    .Y(_0473_)
  );
  \$_AND_  _1078_ (
    .A(_0470_),
    .B(_0467_),
    .Y(_0474_)
  );
  \$_OR_  _1079_ (
    .A(_0474_),
    .B(_0473_),
    .Y(_0475_)
  );
  \$_XOR_  _1080_ (
    .A(_0475_),
    .B(_0472_),
    .Y(_0476_)
  );
  \$_MUX_  _1081_ (
    .A(_0476_),
    .B(dbg_din[14]),
    .S(_0414_),
    .Y(_0007_[14])
  );
  \$_XOR_  _1082_ (
    .A(_0416_),
    .B(mem_cnt[15]),
    .Y(_0477_)
  );
  \$_AND_  _1083_ (
    .A(_0416_),
    .B(mem_cnt[14]),
    .Y(_0478_)
  );
  \$_AND_  _1084_ (
    .A(_0475_),
    .B(_0472_),
    .Y(_0479_)
  );
  \$_OR_  _1085_ (
    .A(_0479_),
    .B(_0478_),
    .Y(_0480_)
  );
  \$_XOR_  _1086_ (
    .A(_0480_),
    .B(_0477_),
    .Y(_0481_)
  );
  \$_MUX_  _1087_ (
    .A(_0481_),
    .B(dbg_din[15]),
    .S(_0414_),
    .Y(_0007_[15])
  );
  \$_XOR_  _1088_ (
    .A(_0437_),
    .B(_0436_),
    .Y(_0482_)
  );
  \$_MUX_  _1089_ (
    .A(_0482_),
    .B(dbg_din[1]),
    .S(_0414_),
    .Y(_0007_[1])
  );
  \$_XOR_  _1090_ (
    .A(_0439_),
    .B(_0434_),
    .Y(_0483_)
  );
  \$_MUX_  _1091_ (
    .A(_0483_),
    .B(dbg_din[2]),
    .S(_0414_),
    .Y(_0007_[2])
  );
  \$_XOR_  _1092_ (
    .A(_0441_),
    .B(_0432_),
    .Y(_0484_)
  );
  \$_MUX_  _1093_ (
    .A(_0484_),
    .B(dbg_din[3]),
    .S(_0414_),
    .Y(_0007_[3])
  );
  \$_XOR_  _1094_ (
    .A(_0443_),
    .B(_0430_),
    .Y(_0485_)
  );
  \$_MUX_  _1095_ (
    .A(_0485_),
    .B(dbg_din[4]),
    .S(_0414_),
    .Y(_0007_[4])
  );
  \$_XOR_  _1096_ (
    .A(_0445_),
    .B(_0428_),
    .Y(_0486_)
  );
  \$_MUX_  _1097_ (
    .A(_0486_),
    .B(dbg_din[5]),
    .S(_0414_),
    .Y(_0007_[5])
  );
  \$_XOR_  _1098_ (
    .A(_0447_),
    .B(_0426_),
    .Y(_0487_)
  );
  \$_MUX_  _1099_ (
    .A(_0487_),
    .B(dbg_din[6]),
    .S(_0414_),
    .Y(_0007_[6])
  );
  \$_XOR_  _1100_ (
    .A(_0449_),
    .B(_0424_),
    .Y(_0488_)
  );
  \$_MUX_  _1101_ (
    .A(_0488_),
    .B(dbg_din[7]),
    .S(_0414_),
    .Y(_0007_[7])
  );
  \$_XOR_  _1102_ (
    .A(_0451_),
    .B(_0422_),
    .Y(_0489_)
  );
  \$_MUX_  _1103_ (
    .A(_0489_),
    .B(dbg_din[8]),
    .S(_0414_),
    .Y(_0007_[8])
  );
  \$_XOR_  _1104_ (
    .A(_0453_),
    .B(_0420_),
    .Y(_0490_)
  );
  \$_MUX_  _1105_ (
    .A(_0490_),
    .B(dbg_din[9]),
    .S(_0414_),
    .Y(_0007_[9])
  );
  \$_OR_  _1106_ (
    .A(mem_burst_rd),
    .B(mem_burst),
    .Y(_0491_)
  );
  \$_OR_  _1107_ (
    .A(_0285_),
    .B(dbg_mem_rd_dly),
    .Y(_0492_)
  );
  \$_MUX_  _1108_ (
    .A(dbg_rd),
    .B(_0492_),
    .S(_0491_),
    .Y(_0002_)
  );
  \$_AND_  _1109_ (
    .A(dbg_din[2]),
    .B(dbg_halt_st),
    .Y(_0493_)
  );
  \$_AND_  _1110_ (
    .A(_0493_),
    .B(_0043_),
    .Y(_0004_[0])
  );
  \$_OR_  _1111_ (
    .A(_0004_[0]),
    .B(inc_step[0]),
    .Y(_0004_[1])
  );
  \$_INV_  _1112_ (
    .A(_0043_),
    .Y(_0494_)
  );
  \$_INV_  _1113_ (
    .A(dbg_din[1]),
    .Y(_0495_)
  );
  \$_OR_  _1114_ (
    .A(_0044_),
    .B(_0495_),
    .Y(_0496_)
  );
  \$_OR_  _1115_ (
    .A(_0496_),
    .B(_0494_),
    .Y(_0497_)
  );
  \$_OR_  _1116_ (
    .A(_0075_),
    .B(_0066_),
    .Y(_0498_)
  );
  \$_OR_  _1117_ (
    .A(_0498_),
    .B(_0074_),
    .Y(_0499_)
  );
  \$_AND_  _1118_ (
    .A(_0499_),
    .B(_0497_),
    .Y(_0500_)
  );
  \$_AND_  _1119_ (
    .A(_0500_),
    .B(_0108_),
    .Y(_0003_)
  );
  \$_AND_  _1120_ (
    .A(_0112_),
    .B(mem_burst),
    .Y(_0501_)
  );
  \$_OR_  _1121_ (
    .A(_0501_),
    .B(_0114_),
    .Y(_0006_)
  );
  \$_AND_  _1122_ (
    .A(mem_bw),
    .B(_0119_),
    .Y(_0502_)
  );
  \$_AND_  _1123_ (
    .A(_0502_),
    .B(mem_data[0]),
    .Y(_0503_)
  );
  \$_AND_  _1124_ (
    .A(mem_data[0]),
    .B(_0120_),
    .Y(_0504_)
  );
  \$_OR_  _1125_ (
    .A(_0504_),
    .B(_0503_),
    .Y(dbg_mem_dout[0])
  );
  \$_AND_  _1126_ (
    .A(mem_bw),
    .B(dbg_mem_addr[0]),
    .Y(_0505_)
  );
  \$_AND_  _1127_ (
    .A(_0505_),
    .B(mem_data[2]),
    .Y(_0506_)
  );
  \$_AND_  _1128_ (
    .A(mem_data[10]),
    .B(_0120_),
    .Y(_0507_)
  );
  \$_OR_  _1129_ (
    .A(_0507_),
    .B(_0506_),
    .Y(dbg_mem_dout[10])
  );
  \$_AND_  _1130_ (
    .A(_0505_),
    .B(mem_data[3]),
    .Y(_0508_)
  );
  \$_AND_  _1131_ (
    .A(mem_data[11]),
    .B(_0120_),
    .Y(_0509_)
  );
  \$_OR_  _1132_ (
    .A(_0509_),
    .B(_0508_),
    .Y(dbg_mem_dout[11])
  );
  \$_AND_  _1133_ (
    .A(_0505_),
    .B(mem_data[4]),
    .Y(_0510_)
  );
  \$_AND_  _1134_ (
    .A(mem_data[12]),
    .B(_0120_),
    .Y(_0511_)
  );
  \$_OR_  _1135_ (
    .A(_0511_),
    .B(_0510_),
    .Y(dbg_mem_dout[12])
  );
  \$_AND_  _1136_ (
    .A(_0505_),
    .B(mem_data[5]),
    .Y(_0512_)
  );
  \$_AND_  _1137_ (
    .A(mem_data[13]),
    .B(_0120_),
    .Y(_0513_)
  );
  \$_OR_  _1138_ (
    .A(_0513_),
    .B(_0512_),
    .Y(dbg_mem_dout[13])
  );
  \$_AND_  _1139_ (
    .A(_0505_),
    .B(mem_data[6]),
    .Y(_0514_)
  );
  \$_AND_  _1140_ (
    .A(mem_data[14]),
    .B(_0120_),
    .Y(_0515_)
  );
  \$_OR_  _1141_ (
    .A(_0515_),
    .B(_0514_),
    .Y(dbg_mem_dout[14])
  );
  \$_AND_  _1142_ (
    .A(_0505_),
    .B(mem_data[7]),
    .Y(_0516_)
  );
  \$_AND_  _1143_ (
    .A(mem_data[15]),
    .B(_0120_),
    .Y(_0517_)
  );
  \$_OR_  _1144_ (
    .A(_0517_),
    .B(_0516_),
    .Y(dbg_mem_dout[15])
  );
  \$_AND_  _1145_ (
    .A(_0502_),
    .B(mem_data[1]),
    .Y(_0518_)
  );
  \$_AND_  _1146_ (
    .A(mem_data[1]),
    .B(_0120_),
    .Y(_0519_)
  );
  \$_OR_  _1147_ (
    .A(_0519_),
    .B(_0518_),
    .Y(dbg_mem_dout[1])
  );
  \$_AND_  _1148_ (
    .A(_0502_),
    .B(mem_data[2]),
    .Y(_0520_)
  );
  \$_AND_  _1149_ (
    .A(mem_data[2]),
    .B(_0120_),
    .Y(_0521_)
  );
  \$_OR_  _1150_ (
    .A(_0521_),
    .B(_0520_),
    .Y(dbg_mem_dout[2])
  );
  \$_AND_  _1151_ (
    .A(_0502_),
    .B(mem_data[3]),
    .Y(_0522_)
  );
  \$_AND_  _1152_ (
    .A(mem_data[3]),
    .B(_0120_),
    .Y(_0523_)
  );
  \$_OR_  _1153_ (
    .A(_0523_),
    .B(_0522_),
    .Y(dbg_mem_dout[3])
  );
  \$_AND_  _1154_ (
    .A(_0502_),
    .B(mem_data[4]),
    .Y(_0524_)
  );
  \$_AND_  _1155_ (
    .A(mem_data[4]),
    .B(_0120_),
    .Y(_0525_)
  );
  \$_OR_  _1156_ (
    .A(_0525_),
    .B(_0524_),
    .Y(dbg_mem_dout[4])
  );
  \$_AND_  _1157_ (
    .A(_0502_),
    .B(mem_data[5]),
    .Y(_0526_)
  );
  \$_AND_  _1158_ (
    .A(mem_data[5]),
    .B(_0120_),
    .Y(_0527_)
  );
  \$_OR_  _1159_ (
    .A(_0527_),
    .B(_0526_),
    .Y(dbg_mem_dout[5])
  );
  \$_AND_  _1160_ (
    .A(_0502_),
    .B(mem_data[6]),
    .Y(_0528_)
  );
  \$_AND_  _1161_ (
    .A(mem_data[6]),
    .B(_0120_),
    .Y(_0529_)
  );
  \$_OR_  _1162_ (
    .A(_0529_),
    .B(_0528_),
    .Y(dbg_mem_dout[6])
  );
  \$_AND_  _1163_ (
    .A(_0502_),
    .B(mem_data[7]),
    .Y(_0530_)
  );
  \$_AND_  _1164_ (
    .A(mem_data[7]),
    .B(_0120_),
    .Y(_0531_)
  );
  \$_OR_  _1165_ (
    .A(_0531_),
    .B(_0530_),
    .Y(dbg_mem_dout[7])
  );
  \$_AND_  _1166_ (
    .A(_0505_),
    .B(mem_data[0]),
    .Y(_0532_)
  );
  \$_AND_  _1167_ (
    .A(mem_data[8]),
    .B(_0120_),
    .Y(_0533_)
  );
  \$_OR_  _1168_ (
    .A(_0533_),
    .B(_0532_),
    .Y(dbg_mem_dout[8])
  );
  \$_AND_  _1169_ (
    .A(_0505_),
    .B(mem_data[1]),
    .Y(_0534_)
  );
  \$_AND_  _1170_ (
    .A(mem_data[9]),
    .B(_0120_),
    .Y(_0535_)
  );
  \$_OR_  _1171_ (
    .A(_0535_),
    .B(_0534_),
    .Y(dbg_mem_dout[9])
  );
  \$_DFF_PP0_  \mem_state_reg[0]  /* _1172_ */ (
    .C(dbg_clk),
    .D(_0536_),
    .Q(mem_state[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_state_reg[1]  /* _1173_ */ (
    .C(dbg_clk),
    .D(_0538_),
    .Q(mem_state[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_state_reg[2]  /* _1174_ */ (
    .C(dbg_clk),
    .D(_0537_),
    .Q(mem_state[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \cpu_ctl_reg[3]  /* _1175_ */ (
    .C(dbg_clk),
    .D(_0000_[0]),
    .Q(cpu_ctl[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \cpu_ctl_reg[4]  /* _1176_ */ (
    .C(dbg_clk),
    .D(_0000_[1]),
    .Q(cpu_ctl[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \cpu_ctl_reg[5]  /* _1177_ */ (
    .C(dbg_clk),
    .D(_0000_[2]),
    .Q(cpu_ctl[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \cpu_ctl_reg[6]  /* _1178_ */ (
    .C(dbg_clk),
    .D(_0000_[3]),
    .Q(cpu_ctl[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \cpu_stat_reg[2]  /* _1179_ */ (
    .C(dbg_clk),
    .D(_0001_[0]),
    .Q(cpu_stat[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \cpu_stat_reg[3]  /* _1180_ */ (
    .C(dbg_clk),
    .D(_0001_[1]),
    .Q(cpu_stat[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_ctl_reg[1]  /* _1181_ */ (
    .C(dbg_clk),
    .D(_0008_[0]),
    .Q(mem_ctl[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_ctl_reg[2]  /* _1182_ */ (
    .C(dbg_clk),
    .D(_0008_[1]),
    .Q(mem_ctl[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  mem_bw_reg /* _1183_ */ (
    .C(dbg_clk),
    .D(_0008_[2]),
    .Q(mem_bw),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  mem_start_reg /* _1184_ */ (
    .C(dbg_clk),
    .D(_0010_),
    .Q(mem_start),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[0]  /* _1185_ */ (
    .C(dbg_clk),
    .D(_0009_[0]),
    .Q(mem_data[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[10]  /* _1186_ */ (
    .C(dbg_clk),
    .D(_0009_[10]),
    .Q(mem_data[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[11]  /* _1187_ */ (
    .C(dbg_clk),
    .D(_0009_[11]),
    .Q(mem_data[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[12]  /* _1188_ */ (
    .C(dbg_clk),
    .D(_0009_[12]),
    .Q(mem_data[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[13]  /* _1189_ */ (
    .C(dbg_clk),
    .D(_0009_[13]),
    .Q(mem_data[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[14]  /* _1190_ */ (
    .C(dbg_clk),
    .D(_0009_[14]),
    .Q(mem_data[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[15]  /* _1191_ */ (
    .C(dbg_clk),
    .D(_0009_[15]),
    .Q(mem_data[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[1]  /* _1192_ */ (
    .C(dbg_clk),
    .D(_0009_[1]),
    .Q(mem_data[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[2]  /* _1193_ */ (
    .C(dbg_clk),
    .D(_0009_[2]),
    .Q(mem_data[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[3]  /* _1194_ */ (
    .C(dbg_clk),
    .D(_0009_[3]),
    .Q(mem_data[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[4]  /* _1195_ */ (
    .C(dbg_clk),
    .D(_0009_[4]),
    .Q(mem_data[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[5]  /* _1196_ */ (
    .C(dbg_clk),
    .D(_0009_[5]),
    .Q(mem_data[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[6]  /* _1197_ */ (
    .C(dbg_clk),
    .D(_0009_[6]),
    .Q(mem_data[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[7]  /* _1198_ */ (
    .C(dbg_clk),
    .D(_0009_[7]),
    .Q(mem_data[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[8]  /* _1199_ */ (
    .C(dbg_clk),
    .D(_0009_[8]),
    .Q(mem_data[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_data_reg[9]  /* _1200_ */ (
    .C(dbg_clk),
    .D(_0009_[9]),
    .Q(mem_data[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[0]  /* _1201_ */ (
    .C(dbg_clk),
    .D(_0005_[0]),
    .Q(dbg_mem_addr[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[10]  /* _1202_ */ (
    .C(dbg_clk),
    .D(_0005_[10]),
    .Q(dbg_mem_addr[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[11]  /* _1203_ */ (
    .C(dbg_clk),
    .D(_0005_[11]),
    .Q(dbg_mem_addr[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[12]  /* _1204_ */ (
    .C(dbg_clk),
    .D(_0005_[12]),
    .Q(dbg_mem_addr[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[13]  /* _1205_ */ (
    .C(dbg_clk),
    .D(_0005_[13]),
    .Q(dbg_mem_addr[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[14]  /* _1206_ */ (
    .C(dbg_clk),
    .D(_0005_[14]),
    .Q(dbg_mem_addr[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[15]  /* _1207_ */ (
    .C(dbg_clk),
    .D(_0005_[15]),
    .Q(dbg_mem_addr[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[1]  /* _1208_ */ (
    .C(dbg_clk),
    .D(_0005_[1]),
    .Q(dbg_mem_addr[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[2]  /* _1209_ */ (
    .C(dbg_clk),
    .D(_0005_[2]),
    .Q(dbg_mem_addr[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[3]  /* _1210_ */ (
    .C(dbg_clk),
    .D(_0005_[3]),
    .Q(dbg_mem_addr[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[4]  /* _1211_ */ (
    .C(dbg_clk),
    .D(_0005_[4]),
    .Q(dbg_mem_addr[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[5]  /* _1212_ */ (
    .C(dbg_clk),
    .D(_0005_[5]),
    .Q(dbg_mem_addr[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[6]  /* _1213_ */ (
    .C(dbg_clk),
    .D(_0005_[6]),
    .Q(dbg_mem_addr[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[7]  /* _1214_ */ (
    .C(dbg_clk),
    .D(_0005_[7]),
    .Q(dbg_mem_addr[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[8]  /* _1215_ */ (
    .C(dbg_clk),
    .D(_0005_[8]),
    .Q(dbg_mem_addr[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_mem_addr_reg[9]  /* _1216_ */ (
    .C(dbg_clk),
    .D(_0005_[9]),
    .Q(dbg_mem_addr[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[0]  /* _1217_ */ (
    .C(dbg_clk),
    .D(_0007_[0]),
    .Q(mem_cnt[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[10]  /* _1218_ */ (
    .C(dbg_clk),
    .D(_0007_[10]),
    .Q(mem_cnt[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[11]  /* _1219_ */ (
    .C(dbg_clk),
    .D(_0007_[11]),
    .Q(mem_cnt[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[12]  /* _1220_ */ (
    .C(dbg_clk),
    .D(_0007_[12]),
    .Q(mem_cnt[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[13]  /* _1221_ */ (
    .C(dbg_clk),
    .D(_0007_[13]),
    .Q(mem_cnt[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[14]  /* _1222_ */ (
    .C(dbg_clk),
    .D(_0007_[14]),
    .Q(mem_cnt[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[15]  /* _1223_ */ (
    .C(dbg_clk),
    .D(_0007_[15]),
    .Q(mem_cnt[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[1]  /* _1224_ */ (
    .C(dbg_clk),
    .D(_0007_[1]),
    .Q(mem_cnt[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[2]  /* _1225_ */ (
    .C(dbg_clk),
    .D(_0007_[2]),
    .Q(mem_cnt[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[3]  /* _1226_ */ (
    .C(dbg_clk),
    .D(_0007_[3]),
    .Q(mem_cnt[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[4]  /* _1227_ */ (
    .C(dbg_clk),
    .D(_0007_[4]),
    .Q(mem_cnt[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[5]  /* _1228_ */ (
    .C(dbg_clk),
    .D(_0007_[5]),
    .Q(mem_cnt[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[6]  /* _1229_ */ (
    .C(dbg_clk),
    .D(_0007_[6]),
    .Q(mem_cnt[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[7]  /* _1230_ */ (
    .C(dbg_clk),
    .D(_0007_[7]),
    .Q(mem_cnt[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[8]  /* _1231_ */ (
    .C(dbg_clk),
    .D(_0007_[8]),
    .Q(mem_cnt[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \mem_cnt_reg[9]  /* _1232_ */ (
    .C(dbg_clk),
    .D(_0007_[9]),
    .Q(mem_cnt[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  dbg_rd_rdy_reg /* _1233_ */ (
    .C(dbg_clk),
    .D(_0002_),
    .Q(dbg_rd_rdy),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \inc_step_reg[0]  /* _1234_ */ (
    .C(dbg_clk),
    .D(_0004_[0]),
    .Q(inc_step[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \inc_step_reg[1]  /* _1235_ */ (
    .C(dbg_clk),
    .D(_0004_[1]),
    .Q(inc_step[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  halt_flag_reg /* _1236_ */ (
    .C(dbg_clk),
    .D(_0003_),
    .Q(halt_flag),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  mem_burst_reg /* _1237_ */ (
    .C(dbg_clk),
    .D(_0006_),
    .Q(mem_burst),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  mem_startb_reg /* _1238_ */ (
    .C(dbg_clk),
    .D(_0011_),
    .Q(mem_startb),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  dbg_mem_rd_dly_reg /* _1239_ */ (
    .C(dbg_clk),
    .D(dbg_mem_rd),
    .Q(dbg_mem_rd_dly),
    .R(dbg_rst)
  );
  omsp_dbg_uart dbg_uart_0 (
    .dbg_addr(dbg_addr),
    .dbg_clk(dbg_clk),
    .dbg_din(dbg_din),
    .dbg_dout(dbg_dout),
    .dbg_rd(dbg_rd),
    .dbg_rd_rdy(dbg_rd_rdy),
    .dbg_rst(dbg_rst),
    .dbg_uart_rxd(dbg_uart_rxd),
    .dbg_uart_txd(dbg_uart_txd),
    .dbg_wr(dbg_wr),
    .mem_burst(mem_burst),
    .mem_burst_end(mem_burst_end),
    .mem_burst_rd(mem_burst_rd),
    .mem_burst_wr(mem_burst_wr),
    .mem_bw(mem_bw)
  );
  assign cpu_ctl_full = { 1'b0, cpu_ctl, 3'b000 };
  assign cpu_stat_full = { 4'b0000, cpu_stat, 1'b0, dbg_halt_st };
  assign cpu_stat_set[2] = puc_pnd_set;
  assign dbg_cpu_reset = cpu_ctl[6];
  assign mem_addr = dbg_mem_addr;
  assign mem_ctl[3] = mem_bw;
  assign mem_ctl_full = { 4'b0000, mem_bw, mem_ctl[2:1], 1'b0 };
  assign reg_write = dbg_wr;
endmodule

module omsp_dbg_uart(dbg_addr, dbg_din, dbg_rd, dbg_uart_txd, dbg_wr, dbg_clk, dbg_dout, dbg_rd_rdy, dbg_rst, dbg_uart_rxd, mem_burst, mem_burst_end, mem_burst_rd, mem_burst_wr, mem_bw);
  wire [5:0] _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire [18:0] _004_;
  wire [3:0] _005_;
  wire [19:0] _006_;
  wire [15:0] _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire [15:0] bit_cnt_max;
  output [5:0] dbg_addr;
  wire dbg_bw;
  input dbg_clk;
  output [15:0] dbg_din;
  input [15:0] dbg_dout;
  output dbg_rd;
  input dbg_rd_rdy;
  input dbg_rst;
  input dbg_uart_rxd;
  output dbg_uart_txd;
  output dbg_wr;
  input mem_burst;
  input mem_burst_end;
  input mem_burst_rd;
  input mem_burst_wr;
  input mem_bw;
  wire [1:0] rxd_buf;
  wire rxd_maj;
  wire rxd_maj_nxt;
  wire rxd_s;
  wire sync_busy;
  wire [18:0] sync_cnt;
  wire uart_rxd;
  wire uart_rxd_n;
  wire [4:0] uart_state;
  wire [3:0] xfer_bit;
  wire [19:0] xfer_buf;
  wire [19:0] xfer_buf_nxt;
  wire [15:0] xfer_cnt;
  \$_INV_  _286_ (
    .A(uart_rxd_n),
    .Y(uart_rxd)
  );
  \$_AND_  _287_ (
    .A(rxd_buf[1]),
    .B(rxd_buf[0]),
    .Y(_008_)
  );
  \$_AND_  _288_ (
    .A(uart_rxd),
    .B(rxd_buf[0]),
    .Y(_009_)
  );
  \$_AND_  _289_ (
    .A(uart_rxd),
    .B(rxd_buf[1]),
    .Y(_010_)
  );
  \$_OR_  _290_ (
    .A(_010_),
    .B(_009_),
    .Y(_011_)
  );
  \$_OR_  _291_ (
    .A(_011_),
    .B(_008_),
    .Y(rxd_maj_nxt)
  );
  \$_OR_  _292_ (
    .A(uart_state[4]),
    .B(uart_state[2]),
    .Y(_012_)
  );
  \$_OR_  _293_ (
    .A(_012_),
    .B(uart_state[1]),
    .Y(_013_)
  );
  \$_INV_  _294_ (
    .A(xfer_bit[0]),
    .Y(_014_)
  );
  \$_AND_  _295_ (
    .A(xfer_bit[1]),
    .B(_014_),
    .Y(_015_)
  );
  \$_INV_  _296_ (
    .A(xfer_bit[2]),
    .Y(_016_)
  );
  \$_AND_  _297_ (
    .A(xfer_bit[3]),
    .B(_016_),
    .Y(_017_)
  );
  \$_AND_  _298_ (
    .A(_017_),
    .B(_015_),
    .Y(_018_)
  );
  \$_AND_  _299_ (
    .A(_018_),
    .B(_013_),
    .Y(_019_)
  );
  \$_AND_  _300_ (
    .A(xfer_bit[1]),
    .B(xfer_bit[0]),
    .Y(_020_)
  );
  \$_AND_  _301_ (
    .A(_020_),
    .B(_016_),
    .Y(_021_)
  );
  \$_INV_  _302_ (
    .A(_013_),
    .Y(_022_)
  );
  \$_AND_  _303_ (
    .A(_022_),
    .B(xfer_bit[3]),
    .Y(_023_)
  );
  \$_AND_  _304_ (
    .A(_023_),
    .B(_021_),
    .Y(_024_)
  );
  \$_OR_  _305_ (
    .A(_024_),
    .B(_019_),
    .Y(_025_)
  );
  \$_AND_  _306_ (
    .A(_025_),
    .B(uart_state[4]),
    .Y(dbg_wr)
  );
  \$_INV_  _307_ (
    .A(mem_bw),
    .Y(_026_)
  );
  \$_OR_  _308_ (
    .A(uart_state[3]),
    .B(uart_state[0]),
    .Y(_027_)
  );
  \$_INV_  _309_ (
    .A(_027_),
    .Y(_028_)
  );
  \$_AND_  _310_ (
    .A(_028_),
    .B(_022_),
    .Y(_029_)
  );
  \$_INV_  _311_ (
    .A(rxd_maj),
    .Y(_030_)
  );
  \$_AND_  _312_ (
    .A(rxd_maj_nxt),
    .B(_030_),
    .Y(_031_)
  );
  \$_AND_  _313_ (
    .A(_031_),
    .B(_029_),
    .Y(_032_)
  );
  \$_AND_  _314_ (
    .A(_032_),
    .B(sync_busy),
    .Y(_033_)
  );
  \$_INV_  _315_ (
    .A(_033_),
    .Y(_034_)
  );
  \$_INV_  _316_ (
    .A(_025_),
    .Y(_035_)
  );
  \$_OR_  _317_ (
    .A(mem_burst_rd),
    .B(mem_burst_wr),
    .Y(_036_)
  );
  \$_INV_  _318_ (
    .A(_036_),
    .Y(_037_)
  );
  \$_AND_  _319_ (
    .A(_037_),
    .B(_035_),
    .Y(_038_)
  );
  \$_AND_  _320_ (
    .A(_038_),
    .B(_034_),
    .Y(_039_)
  );
  \$_INV_  _321_ (
    .A(_039_),
    .Y(_040_)
  );
  \$_INV_  _322_ (
    .A(mem_burst),
    .Y(_041_)
  );
  \$_OR_  _323_ (
    .A(mem_burst_end),
    .B(_041_),
    .Y(_042_)
  );
  \$_INV_  _324_ (
    .A(_042_),
    .Y(_043_)
  );
  \$_AND_  _325_ (
    .A(_043_),
    .B(_040_),
    .Y(_044_)
  );
  \$_AND_  _326_ (
    .A(_044_),
    .B(_026_),
    .Y(_045_)
  );
  \$_AND_  _327_ (
    .A(_045_),
    .B(uart_state[3]),
    .Y(_046_)
  );
  \$_INV_  _328_ (
    .A(xfer_buf[19]),
    .Y(_047_)
  );
  \$_AND_  _329_ (
    .A(_040_),
    .B(_037_),
    .Y(_048_)
  );
  \$_AND_  _330_ (
    .A(_048_),
    .B(_047_),
    .Y(_049_)
  );
  \$_INV_  _331_ (
    .A(xfer_buf[18]),
    .Y(_050_)
  );
  \$_AND_  _332_ (
    .A(_050_),
    .B(uart_state[2]),
    .Y(_051_)
  );
  \$_AND_  _333_ (
    .A(_051_),
    .B(_049_),
    .Y(_052_)
  );
  \$_AND_  _334_ (
    .A(_040_),
    .B(_026_),
    .Y(_053_)
  );
  \$_INV_  _335_ (
    .A(mem_burst_wr),
    .Y(_054_)
  );
  \$_AND_  _336_ (
    .A(_054_),
    .B(uart_state[2]),
    .Y(_055_)
  );
  \$_AND_  _337_ (
    .A(_055_),
    .B(mem_burst_rd),
    .Y(_056_)
  );
  \$_AND_  _338_ (
    .A(_056_),
    .B(_053_),
    .Y(_057_)
  );
  \$_AND_  _339_ (
    .A(_039_),
    .B(uart_state[0]),
    .Y(_058_)
  );
  \$_OR_  _340_ (
    .A(_058_),
    .B(_057_),
    .Y(_059_)
  );
  \$_OR_  _341_ (
    .A(_059_),
    .B(_052_),
    .Y(_060_)
  );
  \$_OR_  _342_ (
    .A(_060_),
    .B(_046_),
    .Y(_280_)
  );
  \$_AND_  _343_ (
    .A(_045_),
    .B(uart_state[4]),
    .Y(_061_)
  );
  \$_AND_  _344_ (
    .A(_048_),
    .B(xfer_buf[19]),
    .Y(_062_)
  );
  \$_AND_  _345_ (
    .A(_062_),
    .B(_051_),
    .Y(_063_)
  );
  \$_AND_  _346_ (
    .A(mem_burst_wr),
    .B(uart_state[2]),
    .Y(_064_)
  );
  \$_AND_  _347_ (
    .A(_064_),
    .B(_053_),
    .Y(_065_)
  );
  \$_AND_  _348_ (
    .A(_039_),
    .B(uart_state[1]),
    .Y(_066_)
  );
  \$_OR_  _349_ (
    .A(_066_),
    .B(_065_),
    .Y(_067_)
  );
  \$_OR_  _350_ (
    .A(_067_),
    .B(_063_),
    .Y(_068_)
  );
  \$_OR_  _351_ (
    .A(_068_),
    .B(_061_),
    .Y(_281_)
  );
  \$_AND_  _352_ (
    .A(_039_),
    .B(uart_state[2]),
    .Y(_069_)
  );
  \$_AND_  _353_ (
    .A(_040_),
    .B(_029_),
    .Y(_070_)
  );
  \$_OR_  _354_ (
    .A(uart_state[3]),
    .B(uart_state[4]),
    .Y(_071_)
  );
  \$_AND_  _355_ (
    .A(_071_),
    .B(_042_),
    .Y(_072_)
  );
  \$_AND_  _356_ (
    .A(_072_),
    .B(_040_),
    .Y(_073_)
  );
  \$_OR_  _357_ (
    .A(_073_),
    .B(_070_),
    .Y(_074_)
  );
  \$_OR_  _358_ (
    .A(_074_),
    .B(_069_),
    .Y(_282_)
  );
  \$_AND_  _359_ (
    .A(_044_),
    .B(mem_bw),
    .Y(_075_)
  );
  \$_AND_  _360_ (
    .A(_075_),
    .B(uart_state[3]),
    .Y(_076_)
  );
  \$_AND_  _361_ (
    .A(xfer_buf[18]),
    .B(uart_state[2]),
    .Y(_077_)
  );
  \$_AND_  _362_ (
    .A(_077_),
    .B(_049_),
    .Y(_078_)
  );
  \$_AND_  _363_ (
    .A(_040_),
    .B(mem_bw),
    .Y(_079_)
  );
  \$_AND_  _364_ (
    .A(_079_),
    .B(_056_),
    .Y(_080_)
  );
  \$_MUX_  _365_ (
    .A(uart_state[0]),
    .B(uart_state[3]),
    .S(_039_),
    .Y(_081_)
  );
  \$_OR_  _366_ (
    .A(_081_),
    .B(_080_),
    .Y(_082_)
  );
  \$_OR_  _367_ (
    .A(_082_),
    .B(_078_),
    .Y(_083_)
  );
  \$_OR_  _368_ (
    .A(_083_),
    .B(_076_),
    .Y(_283_)
  );
  \$_AND_  _369_ (
    .A(_075_),
    .B(uart_state[4]),
    .Y(_084_)
  );
  \$_AND_  _370_ (
    .A(_077_),
    .B(_062_),
    .Y(_085_)
  );
  \$_AND_  _371_ (
    .A(_079_),
    .B(_064_),
    .Y(_086_)
  );
  \$_MUX_  _372_ (
    .A(uart_state[1]),
    .B(uart_state[4]),
    .S(_039_),
    .Y(_087_)
  );
  \$_OR_  _373_ (
    .A(_087_),
    .B(_086_),
    .Y(_088_)
  );
  \$_OR_  _374_ (
    .A(_088_),
    .B(_085_),
    .Y(_089_)
  );
  \$_OR_  _375_ (
    .A(_089_),
    .B(_084_),
    .Y(_284_)
  );
  \$_INV_  _376_ (
    .A(dbg_uart_rxd),
    .Y(_285_)
  );
  \$_INV_  _377_ (
    .A(rxd_maj_nxt),
    .Y(_090_)
  );
  \$_AND_  _378_ (
    .A(_090_),
    .B(rxd_maj),
    .Y(_091_)
  );
  \$_AND_  _379_ (
    .A(_091_),
    .B(_029_),
    .Y(_092_)
  );
  \$_INV_  _380_ (
    .A(_032_),
    .Y(_093_)
  );
  \$_AND_  _381_ (
    .A(_093_),
    .B(sync_busy),
    .Y(_094_)
  );
  \$_OR_  _382_ (
    .A(_094_),
    .B(_092_),
    .Y(_003_)
  );
  \$_OR_  _383_ (
    .A(sync_busy),
    .B(sync_cnt[2]),
    .Y(_095_)
  );
  \$_XOR_  _384_ (
    .A(_095_),
    .B(sync_cnt[0]),
    .Y(_004_[0])
  );
  \$_INV_  _385_ (
    .A(_095_),
    .Y(_096_)
  );
  \$_AND_  _386_ (
    .A(sync_cnt[1]),
    .B(sync_cnt[0]),
    .Y(_097_)
  );
  \$_AND_  _387_ (
    .A(_097_),
    .B(sync_cnt[2]),
    .Y(_098_)
  );
  \$_AND_  _388_ (
    .A(_098_),
    .B(bit_cnt_max[0]),
    .Y(_099_)
  );
  \$_AND_  _389_ (
    .A(_099_),
    .B(bit_cnt_max[1]),
    .Y(_100_)
  );
  \$_AND_  _390_ (
    .A(_100_),
    .B(bit_cnt_max[2]),
    .Y(_101_)
  );
  \$_AND_  _391_ (
    .A(_101_),
    .B(bit_cnt_max[3]),
    .Y(_102_)
  );
  \$_AND_  _392_ (
    .A(_102_),
    .B(bit_cnt_max[4]),
    .Y(_103_)
  );
  \$_AND_  _393_ (
    .A(_103_),
    .B(bit_cnt_max[5]),
    .Y(_104_)
  );
  \$_AND_  _394_ (
    .A(_104_),
    .B(bit_cnt_max[6]),
    .Y(_105_)
  );
  \$_XOR_  _395_ (
    .A(_105_),
    .B(bit_cnt_max[7]),
    .Y(_106_)
  );
  \$_MUX_  _396_ (
    .A(_106_),
    .B(bit_cnt_max[7]),
    .S(_096_),
    .Y(_004_[10])
  );
  \$_AND_  _397_ (
    .A(_105_),
    .B(bit_cnt_max[7]),
    .Y(_107_)
  );
  \$_XOR_  _398_ (
    .A(_107_),
    .B(bit_cnt_max[8]),
    .Y(_108_)
  );
  \$_MUX_  _399_ (
    .A(_108_),
    .B(bit_cnt_max[8]),
    .S(_096_),
    .Y(_004_[11])
  );
  \$_AND_  _400_ (
    .A(_107_),
    .B(bit_cnt_max[8]),
    .Y(_109_)
  );
  \$_XOR_  _401_ (
    .A(_109_),
    .B(bit_cnt_max[9]),
    .Y(_110_)
  );
  \$_MUX_  _402_ (
    .A(_110_),
    .B(bit_cnt_max[9]),
    .S(_096_),
    .Y(_004_[12])
  );
  \$_AND_  _403_ (
    .A(_109_),
    .B(bit_cnt_max[9]),
    .Y(_111_)
  );
  \$_XOR_  _404_ (
    .A(_111_),
    .B(bit_cnt_max[10]),
    .Y(_112_)
  );
  \$_MUX_  _405_ (
    .A(_112_),
    .B(bit_cnt_max[10]),
    .S(_096_),
    .Y(_004_[13])
  );
  \$_AND_  _406_ (
    .A(_111_),
    .B(bit_cnt_max[10]),
    .Y(_113_)
  );
  \$_XOR_  _407_ (
    .A(_113_),
    .B(bit_cnt_max[11]),
    .Y(_114_)
  );
  \$_MUX_  _408_ (
    .A(_114_),
    .B(bit_cnt_max[11]),
    .S(_096_),
    .Y(_004_[14])
  );
  \$_AND_  _409_ (
    .A(_113_),
    .B(bit_cnt_max[11]),
    .Y(_115_)
  );
  \$_XOR_  _410_ (
    .A(_115_),
    .B(bit_cnt_max[12]),
    .Y(_116_)
  );
  \$_MUX_  _411_ (
    .A(_116_),
    .B(bit_cnt_max[12]),
    .S(_096_),
    .Y(_004_[15])
  );
  \$_AND_  _412_ (
    .A(_115_),
    .B(bit_cnt_max[12]),
    .Y(_117_)
  );
  \$_XOR_  _413_ (
    .A(_117_),
    .B(bit_cnt_max[13]),
    .Y(_118_)
  );
  \$_MUX_  _414_ (
    .A(_118_),
    .B(bit_cnt_max[13]),
    .S(_096_),
    .Y(_004_[16])
  );
  \$_AND_  _415_ (
    .A(_117_),
    .B(bit_cnt_max[13]),
    .Y(_119_)
  );
  \$_XOR_  _416_ (
    .A(_119_),
    .B(bit_cnt_max[14]),
    .Y(_120_)
  );
  \$_MUX_  _417_ (
    .A(_120_),
    .B(bit_cnt_max[14]),
    .S(_096_),
    .Y(_004_[17])
  );
  \$_AND_  _418_ (
    .A(_119_),
    .B(bit_cnt_max[14]),
    .Y(_121_)
  );
  \$_XOR_  _419_ (
    .A(_121_),
    .B(bit_cnt_max[15]),
    .Y(_122_)
  );
  \$_MUX_  _420_ (
    .A(_122_),
    .B(bit_cnt_max[15]),
    .S(_096_),
    .Y(_004_[18])
  );
  \$_XOR_  _421_ (
    .A(sync_cnt[1]),
    .B(sync_cnt[0]),
    .Y(_123_)
  );
  \$_MUX_  _422_ (
    .A(sync_cnt[1]),
    .B(_123_),
    .S(_095_),
    .Y(_004_[1])
  );
  \$_XOR_  _423_ (
    .A(_097_),
    .B(sync_cnt[2]),
    .Y(_124_)
  );
  \$_MUX_  _424_ (
    .A(_124_),
    .B(sync_cnt[2]),
    .S(_096_),
    .Y(_004_[2])
  );
  \$_XOR_  _425_ (
    .A(_098_),
    .B(bit_cnt_max[0]),
    .Y(_125_)
  );
  \$_MUX_  _426_ (
    .A(_125_),
    .B(bit_cnt_max[0]),
    .S(_096_),
    .Y(_004_[3])
  );
  \$_XOR_  _427_ (
    .A(_099_),
    .B(bit_cnt_max[1]),
    .Y(_126_)
  );
  \$_MUX_  _428_ (
    .A(_126_),
    .B(bit_cnt_max[1]),
    .S(_096_),
    .Y(_004_[4])
  );
  \$_XOR_  _429_ (
    .A(_100_),
    .B(bit_cnt_max[2]),
    .Y(_127_)
  );
  \$_MUX_  _430_ (
    .A(_127_),
    .B(bit_cnt_max[2]),
    .S(_096_),
    .Y(_004_[5])
  );
  \$_XOR_  _431_ (
    .A(_101_),
    .B(bit_cnt_max[3]),
    .Y(_128_)
  );
  \$_MUX_  _432_ (
    .A(_128_),
    .B(bit_cnt_max[3]),
    .S(_096_),
    .Y(_004_[6])
  );
  \$_XOR_  _433_ (
    .A(_102_),
    .B(bit_cnt_max[4]),
    .Y(_129_)
  );
  \$_MUX_  _434_ (
    .A(_129_),
    .B(bit_cnt_max[4]),
    .S(_096_),
    .Y(_004_[7])
  );
  \$_XOR_  _435_ (
    .A(_103_),
    .B(bit_cnt_max[5]),
    .Y(_130_)
  );
  \$_MUX_  _436_ (
    .A(_130_),
    .B(bit_cnt_max[5]),
    .S(_096_),
    .Y(_004_[8])
  );
  \$_XOR_  _437_ (
    .A(_104_),
    .B(bit_cnt_max[6]),
    .Y(_131_)
  );
  \$_MUX_  _438_ (
    .A(_131_),
    .B(bit_cnt_max[6]),
    .S(_096_),
    .Y(_004_[9])
  );
  \$_AND_  _439_ (
    .A(_025_),
    .B(uart_state[0]),
    .Y(_132_)
  );
  \$_OR_  _440_ (
    .A(_132_),
    .B(dbg_rd_rdy),
    .Y(_133_)
  );
  \$_OR_  _441_ (
    .A(xfer_bit[1]),
    .B(xfer_bit[0]),
    .Y(_134_)
  );
  \$_OR_  _442_ (
    .A(xfer_bit[3]),
    .B(xfer_bit[2]),
    .Y(_135_)
  );
  \$_OR_  _443_ (
    .A(_135_),
    .B(_134_),
    .Y(_136_)
  );
  \$_OR_  _444_ (
    .A(_136_),
    .B(_029_),
    .Y(_137_)
  );
  \$_INV_  _445_ (
    .A(_137_),
    .Y(_138_)
  );
  \$_AND_  _446_ (
    .A(_138_),
    .B(_091_),
    .Y(_139_)
  );
  \$_OR_  _447_ (
    .A(_139_),
    .B(_133_),
    .Y(_140_)
  );
  \$_INV_  _448_ (
    .A(xfer_cnt[12]),
    .Y(_141_)
  );
  \$_INV_  _449_ (
    .A(xfer_cnt[13]),
    .Y(_142_)
  );
  \$_AND_  _450_ (
    .A(_142_),
    .B(_141_),
    .Y(_143_)
  );
  \$_INV_  _451_ (
    .A(xfer_cnt[14]),
    .Y(_144_)
  );
  \$_INV_  _452_ (
    .A(xfer_cnt[15]),
    .Y(_145_)
  );
  \$_AND_  _453_ (
    .A(_145_),
    .B(_144_),
    .Y(_146_)
  );
  \$_AND_  _454_ (
    .A(_146_),
    .B(_143_),
    .Y(_147_)
  );
  \$_OR_  _455_ (
    .A(xfer_cnt[1]),
    .B(xfer_cnt[0]),
    .Y(_148_)
  );
  \$_INV_  _456_ (
    .A(_148_),
    .Y(_149_)
  );
  \$_INV_  _457_ (
    .A(xfer_cnt[10]),
    .Y(_150_)
  );
  \$_INV_  _458_ (
    .A(xfer_cnt[11]),
    .Y(_151_)
  );
  \$_AND_  _459_ (
    .A(_151_),
    .B(_150_),
    .Y(_152_)
  );
  \$_AND_  _460_ (
    .A(_152_),
    .B(_149_),
    .Y(_153_)
  );
  \$_AND_  _461_ (
    .A(_153_),
    .B(_147_),
    .Y(_154_)
  );
  \$_INV_  _462_ (
    .A(xfer_cnt[6]),
    .Y(_155_)
  );
  \$_INV_  _463_ (
    .A(xfer_cnt[7]),
    .Y(_156_)
  );
  \$_AND_  _464_ (
    .A(_156_),
    .B(_155_),
    .Y(_157_)
  );
  \$_INV_  _465_ (
    .A(xfer_cnt[8]),
    .Y(_158_)
  );
  \$_INV_  _466_ (
    .A(xfer_cnt[9]),
    .Y(_159_)
  );
  \$_AND_  _467_ (
    .A(_159_),
    .B(_158_),
    .Y(_160_)
  );
  \$_AND_  _468_ (
    .A(_160_),
    .B(_157_),
    .Y(_161_)
  );
  \$_INV_  _469_ (
    .A(xfer_cnt[2]),
    .Y(_162_)
  );
  \$_INV_  _470_ (
    .A(xfer_cnt[3]),
    .Y(_163_)
  );
  \$_AND_  _471_ (
    .A(_163_),
    .B(_162_),
    .Y(_164_)
  );
  \$_INV_  _472_ (
    .A(xfer_cnt[4]),
    .Y(_165_)
  );
  \$_INV_  _473_ (
    .A(xfer_cnt[5]),
    .Y(_166_)
  );
  \$_AND_  _474_ (
    .A(_166_),
    .B(_165_),
    .Y(_167_)
  );
  \$_AND_  _475_ (
    .A(_167_),
    .B(_164_),
    .Y(_168_)
  );
  \$_AND_  _476_ (
    .A(_168_),
    .B(_161_),
    .Y(_169_)
  );
  \$_AND_  _477_ (
    .A(_169_),
    .B(_154_),
    .Y(_170_)
  );
  \$_AND_  _478_ (
    .A(_170_),
    .B(_136_),
    .Y(_171_)
  );
  \$_XOR_  _479_ (
    .A(_171_),
    .B(xfer_bit[0]),
    .Y(_172_)
  );
  \$_AND_  _480_ (
    .A(_172_),
    .B(_035_),
    .Y(_173_)
  );
  \$_OR_  _481_ (
    .A(_173_),
    .B(_140_),
    .Y(_005_[0])
  );
  \$_INV_  _482_ (
    .A(_140_),
    .Y(_174_)
  );
  \$_XOR_  _483_ (
    .A(xfer_bit[1]),
    .B(xfer_bit[0]),
    .Y(_175_)
  );
  \$_MUX_  _484_ (
    .A(xfer_bit[1]),
    .B(_175_),
    .S(_171_),
    .Y(_176_)
  );
  \$_AND_  _485_ (
    .A(_176_),
    .B(_035_),
    .Y(_177_)
  );
  \$_AND_  _486_ (
    .A(_177_),
    .B(_174_),
    .Y(_005_[1])
  );
  \$_XOR_  _487_ (
    .A(_020_),
    .B(xfer_bit[2]),
    .Y(_178_)
  );
  \$_MUX_  _488_ (
    .A(xfer_bit[2]),
    .B(_178_),
    .S(_171_),
    .Y(_179_)
  );
  \$_AND_  _489_ (
    .A(_179_),
    .B(_035_),
    .Y(_180_)
  );
  \$_AND_  _490_ (
    .A(_180_),
    .B(_174_),
    .Y(_005_[2])
  );
  \$_AND_  _491_ (
    .A(_020_),
    .B(xfer_bit[2]),
    .Y(_181_)
  );
  \$_XOR_  _492_ (
    .A(_181_),
    .B(xfer_bit[3]),
    .Y(_182_)
  );
  \$_MUX_  _493_ (
    .A(xfer_bit[3]),
    .B(_182_),
    .S(_171_),
    .Y(_183_)
  );
  \$_AND_  _494_ (
    .A(_183_),
    .B(_035_),
    .Y(_184_)
  );
  \$_AND_  _495_ (
    .A(_184_),
    .B(_174_),
    .Y(_005_[3])
  );
  \$_XOR_  _496_ (
    .A(rxd_maj_nxt),
    .B(_030_),
    .Y(_185_)
  );
  \$_OR_  _497_ (
    .A(_185_),
    .B(_022_),
    .Y(_186_)
  );
  \$_INV_  _498_ (
    .A(_186_),
    .Y(_187_)
  );
  \$_OR_  _499_ (
    .A(_171_),
    .B(_133_),
    .Y(_188_)
  );
  \$_INV_  _500_ (
    .A(xfer_cnt[0]),
    .Y(_189_)
  );
  \$_XOR_  _501_ (
    .A(_170_),
    .B(_189_),
    .Y(_190_)
  );
  \$_MUX_  _502_ (
    .A(_190_),
    .B(bit_cnt_max[0]),
    .S(_188_),
    .Y(_191_)
  );
  \$_MUX_  _503_ (
    .A(_191_),
    .B(bit_cnt_max[1]),
    .S(_187_),
    .Y(_007_[0])
  );
  \$_OR_  _504_ (
    .A(_148_),
    .B(xfer_cnt[2]),
    .Y(_192_)
  );
  \$_OR_  _505_ (
    .A(_192_),
    .B(xfer_cnt[3]),
    .Y(_193_)
  );
  \$_OR_  _506_ (
    .A(_193_),
    .B(xfer_cnt[4]),
    .Y(_194_)
  );
  \$_OR_  _507_ (
    .A(_194_),
    .B(xfer_cnt[5]),
    .Y(_195_)
  );
  \$_OR_  _508_ (
    .A(_195_),
    .B(xfer_cnt[6]),
    .Y(_196_)
  );
  \$_OR_  _509_ (
    .A(_196_),
    .B(xfer_cnt[7]),
    .Y(_197_)
  );
  \$_OR_  _510_ (
    .A(_197_),
    .B(xfer_cnt[8]),
    .Y(_198_)
  );
  \$_OR_  _511_ (
    .A(_198_),
    .B(xfer_cnt[9]),
    .Y(_199_)
  );
  \$_XOR_  _512_ (
    .A(_199_),
    .B(_150_),
    .Y(_200_)
  );
  \$_MUX_  _513_ (
    .A(_200_),
    .B(xfer_cnt[10]),
    .S(_170_),
    .Y(_201_)
  );
  \$_MUX_  _514_ (
    .A(_201_),
    .B(bit_cnt_max[10]),
    .S(_188_),
    .Y(_202_)
  );
  \$_MUX_  _515_ (
    .A(_202_),
    .B(bit_cnt_max[11]),
    .S(_187_),
    .Y(_007_[10])
  );
  \$_OR_  _516_ (
    .A(_199_),
    .B(xfer_cnt[10]),
    .Y(_203_)
  );
  \$_XOR_  _517_ (
    .A(_203_),
    .B(_151_),
    .Y(_204_)
  );
  \$_MUX_  _518_ (
    .A(_204_),
    .B(xfer_cnt[11]),
    .S(_170_),
    .Y(_205_)
  );
  \$_MUX_  _519_ (
    .A(_205_),
    .B(bit_cnt_max[11]),
    .S(_188_),
    .Y(_206_)
  );
  \$_MUX_  _520_ (
    .A(_206_),
    .B(bit_cnt_max[12]),
    .S(_187_),
    .Y(_007_[11])
  );
  \$_OR_  _521_ (
    .A(_203_),
    .B(xfer_cnt[11]),
    .Y(_207_)
  );
  \$_XOR_  _522_ (
    .A(_207_),
    .B(_141_),
    .Y(_208_)
  );
  \$_MUX_  _523_ (
    .A(_208_),
    .B(xfer_cnt[12]),
    .S(_170_),
    .Y(_209_)
  );
  \$_MUX_  _524_ (
    .A(_209_),
    .B(bit_cnt_max[12]),
    .S(_188_),
    .Y(_210_)
  );
  \$_MUX_  _525_ (
    .A(_210_),
    .B(bit_cnt_max[13]),
    .S(_187_),
    .Y(_007_[12])
  );
  \$_OR_  _526_ (
    .A(_207_),
    .B(xfer_cnt[12]),
    .Y(_211_)
  );
  \$_XOR_  _527_ (
    .A(_211_),
    .B(_142_),
    .Y(_212_)
  );
  \$_MUX_  _528_ (
    .A(_212_),
    .B(xfer_cnt[13]),
    .S(_170_),
    .Y(_213_)
  );
  \$_MUX_  _529_ (
    .A(_213_),
    .B(bit_cnt_max[13]),
    .S(_188_),
    .Y(_214_)
  );
  \$_MUX_  _530_ (
    .A(_214_),
    .B(bit_cnt_max[14]),
    .S(_187_),
    .Y(_007_[13])
  );
  \$_OR_  _531_ (
    .A(_211_),
    .B(xfer_cnt[13]),
    .Y(_215_)
  );
  \$_XOR_  _532_ (
    .A(_215_),
    .B(_144_),
    .Y(_216_)
  );
  \$_MUX_  _533_ (
    .A(_216_),
    .B(xfer_cnt[14]),
    .S(_170_),
    .Y(_217_)
  );
  \$_MUX_  _534_ (
    .A(_217_),
    .B(bit_cnt_max[14]),
    .S(_188_),
    .Y(_218_)
  );
  \$_MUX_  _535_ (
    .A(_218_),
    .B(bit_cnt_max[15]),
    .S(_187_),
    .Y(_007_[14])
  );
  \$_OR_  _536_ (
    .A(_215_),
    .B(xfer_cnt[14]),
    .Y(_219_)
  );
  \$_XOR_  _537_ (
    .A(_219_),
    .B(_145_),
    .Y(_220_)
  );
  \$_MUX_  _538_ (
    .A(_220_),
    .B(xfer_cnt[15]),
    .S(_170_),
    .Y(_221_)
  );
  \$_MUX_  _539_ (
    .A(_221_),
    .B(bit_cnt_max[15]),
    .S(_188_),
    .Y(_222_)
  );
  \$_AND_  _540_ (
    .A(_222_),
    .B(_186_),
    .Y(_007_[15])
  );
  \$_XOR_  _541_ (
    .A(xfer_cnt[1]),
    .B(_189_),
    .Y(_223_)
  );
  \$_MUX_  _542_ (
    .A(_223_),
    .B(xfer_cnt[1]),
    .S(_170_),
    .Y(_224_)
  );
  \$_MUX_  _543_ (
    .A(_224_),
    .B(bit_cnt_max[1]),
    .S(_188_),
    .Y(_225_)
  );
  \$_MUX_  _544_ (
    .A(_225_),
    .B(bit_cnt_max[2]),
    .S(_187_),
    .Y(_007_[1])
  );
  \$_XOR_  _545_ (
    .A(_148_),
    .B(_162_),
    .Y(_226_)
  );
  \$_MUX_  _546_ (
    .A(_226_),
    .B(xfer_cnt[2]),
    .S(_170_),
    .Y(_227_)
  );
  \$_MUX_  _547_ (
    .A(_227_),
    .B(bit_cnt_max[2]),
    .S(_188_),
    .Y(_228_)
  );
  \$_MUX_  _548_ (
    .A(_228_),
    .B(bit_cnt_max[3]),
    .S(_187_),
    .Y(_007_[2])
  );
  \$_XOR_  _549_ (
    .A(_192_),
    .B(_163_),
    .Y(_229_)
  );
  \$_MUX_  _550_ (
    .A(_229_),
    .B(xfer_cnt[3]),
    .S(_170_),
    .Y(_230_)
  );
  \$_MUX_  _551_ (
    .A(_230_),
    .B(bit_cnt_max[3]),
    .S(_188_),
    .Y(_231_)
  );
  \$_MUX_  _552_ (
    .A(_231_),
    .B(bit_cnt_max[4]),
    .S(_187_),
    .Y(_007_[3])
  );
  \$_XOR_  _553_ (
    .A(_193_),
    .B(_165_),
    .Y(_232_)
  );
  \$_MUX_  _554_ (
    .A(_232_),
    .B(xfer_cnt[4]),
    .S(_170_),
    .Y(_233_)
  );
  \$_MUX_  _555_ (
    .A(_233_),
    .B(bit_cnt_max[4]),
    .S(_188_),
    .Y(_234_)
  );
  \$_MUX_  _556_ (
    .A(_234_),
    .B(bit_cnt_max[5]),
    .S(_187_),
    .Y(_007_[4])
  );
  \$_XOR_  _557_ (
    .A(_194_),
    .B(_166_),
    .Y(_235_)
  );
  \$_MUX_  _558_ (
    .A(_235_),
    .B(xfer_cnt[5]),
    .S(_170_),
    .Y(_236_)
  );
  \$_MUX_  _559_ (
    .A(_236_),
    .B(bit_cnt_max[5]),
    .S(_188_),
    .Y(_237_)
  );
  \$_MUX_  _560_ (
    .A(_237_),
    .B(bit_cnt_max[6]),
    .S(_187_),
    .Y(_007_[5])
  );
  \$_XOR_  _561_ (
    .A(_195_),
    .B(_155_),
    .Y(_238_)
  );
  \$_MUX_  _562_ (
    .A(_238_),
    .B(xfer_cnt[6]),
    .S(_170_),
    .Y(_239_)
  );
  \$_MUX_  _563_ (
    .A(_239_),
    .B(bit_cnt_max[6]),
    .S(_188_),
    .Y(_240_)
  );
  \$_MUX_  _564_ (
    .A(_240_),
    .B(bit_cnt_max[7]),
    .S(_187_),
    .Y(_007_[6])
  );
  \$_XOR_  _565_ (
    .A(_196_),
    .B(_156_),
    .Y(_241_)
  );
  \$_MUX_  _566_ (
    .A(_241_),
    .B(xfer_cnt[7]),
    .S(_170_),
    .Y(_242_)
  );
  \$_MUX_  _567_ (
    .A(_242_),
    .B(bit_cnt_max[7]),
    .S(_188_),
    .Y(_243_)
  );
  \$_MUX_  _568_ (
    .A(_243_),
    .B(bit_cnt_max[8]),
    .S(_187_),
    .Y(_007_[7])
  );
  \$_XOR_  _569_ (
    .A(_197_),
    .B(_158_),
    .Y(_244_)
  );
  \$_MUX_  _570_ (
    .A(_244_),
    .B(xfer_cnt[8]),
    .S(_170_),
    .Y(_245_)
  );
  \$_MUX_  _571_ (
    .A(_245_),
    .B(bit_cnt_max[8]),
    .S(_188_),
    .Y(_246_)
  );
  \$_MUX_  _572_ (
    .A(_246_),
    .B(bit_cnt_max[9]),
    .S(_187_),
    .Y(_007_[8])
  );
  \$_XOR_  _573_ (
    .A(_198_),
    .B(_159_),
    .Y(_247_)
  );
  \$_MUX_  _574_ (
    .A(_247_),
    .B(xfer_cnt[9]),
    .S(_170_),
    .Y(_248_)
  );
  \$_MUX_  _575_ (
    .A(_248_),
    .B(bit_cnt_max[9]),
    .S(_188_),
    .Y(_249_)
  );
  \$_MUX_  _576_ (
    .A(_249_),
    .B(bit_cnt_max[10]),
    .S(_187_),
    .Y(_007_[9])
  );
  \$_INV_  _577_ (
    .A(dbg_rd_rdy),
    .Y(_250_)
  );
  \$_MUX_  _578_ (
    .A(xfer_buf[0]),
    .B(xfer_buf[1]),
    .S(_171_),
    .Y(_251_)
  );
  \$_AND_  _579_ (
    .A(_251_),
    .B(_250_),
    .Y(_006_[0])
  );
  \$_MUX_  _580_ (
    .A(xfer_buf[10]),
    .B(xfer_buf[11]),
    .S(_171_),
    .Y(_252_)
  );
  \$_AND_  _581_ (
    .A(_252_),
    .B(_250_),
    .Y(_006_[10])
  );
  \$_MUX_  _582_ (
    .A(xfer_buf[11]),
    .B(xfer_buf[12]),
    .S(_171_),
    .Y(_253_)
  );
  \$_MUX_  _583_ (
    .A(_253_),
    .B(dbg_dout[8]),
    .S(dbg_rd_rdy),
    .Y(_006_[11])
  );
  \$_MUX_  _584_ (
    .A(xfer_buf[12]),
    .B(xfer_buf[13]),
    .S(_171_),
    .Y(_254_)
  );
  \$_MUX_  _585_ (
    .A(_254_),
    .B(dbg_dout[9]),
    .S(dbg_rd_rdy),
    .Y(_006_[12])
  );
  \$_MUX_  _586_ (
    .A(xfer_buf[13]),
    .B(xfer_buf[14]),
    .S(_171_),
    .Y(_255_)
  );
  \$_MUX_  _587_ (
    .A(_255_),
    .B(dbg_dout[10]),
    .S(dbg_rd_rdy),
    .Y(_006_[13])
  );
  \$_MUX_  _588_ (
    .A(xfer_buf[14]),
    .B(xfer_buf[15]),
    .S(_171_),
    .Y(_256_)
  );
  \$_MUX_  _589_ (
    .A(_256_),
    .B(dbg_dout[11]),
    .S(dbg_rd_rdy),
    .Y(_006_[14])
  );
  \$_MUX_  _590_ (
    .A(xfer_buf[15]),
    .B(xfer_buf[16]),
    .S(_171_),
    .Y(_257_)
  );
  \$_MUX_  _591_ (
    .A(_257_),
    .B(dbg_dout[12]),
    .S(dbg_rd_rdy),
    .Y(_006_[15])
  );
  \$_MUX_  _592_ (
    .A(xfer_buf[16]),
    .B(xfer_buf[17]),
    .S(_171_),
    .Y(_258_)
  );
  \$_MUX_  _593_ (
    .A(_258_),
    .B(dbg_dout[13]),
    .S(dbg_rd_rdy),
    .Y(_006_[16])
  );
  \$_MUX_  _594_ (
    .A(xfer_buf[17]),
    .B(xfer_buf[18]),
    .S(_171_),
    .Y(_259_)
  );
  \$_MUX_  _595_ (
    .A(_259_),
    .B(dbg_dout[14]),
    .S(dbg_rd_rdy),
    .Y(_006_[17])
  );
  \$_MUX_  _596_ (
    .A(xfer_buf[18]),
    .B(xfer_buf[19]),
    .S(_171_),
    .Y(_260_)
  );
  \$_MUX_  _597_ (
    .A(_260_),
    .B(dbg_dout[15]),
    .S(dbg_rd_rdy),
    .Y(_006_[18])
  );
  \$_MUX_  _598_ (
    .A(xfer_buf[19]),
    .B(rxd_maj),
    .S(_171_),
    .Y(_261_)
  );
  \$_OR_  _599_ (
    .A(_261_),
    .B(dbg_rd_rdy),
    .Y(_006_[19])
  );
  \$_MUX_  _600_ (
    .A(xfer_buf[1]),
    .B(xfer_buf[2]),
    .S(_171_),
    .Y(_262_)
  );
  \$_MUX_  _601_ (
    .A(_262_),
    .B(dbg_dout[0]),
    .S(dbg_rd_rdy),
    .Y(_006_[1])
  );
  \$_MUX_  _602_ (
    .A(xfer_buf[2]),
    .B(xfer_buf[3]),
    .S(_171_),
    .Y(_263_)
  );
  \$_MUX_  _603_ (
    .A(_263_),
    .B(dbg_dout[1]),
    .S(dbg_rd_rdy),
    .Y(_006_[2])
  );
  \$_MUX_  _604_ (
    .A(xfer_buf[3]),
    .B(xfer_buf[4]),
    .S(_171_),
    .Y(_264_)
  );
  \$_MUX_  _605_ (
    .A(_264_),
    .B(dbg_dout[2]),
    .S(dbg_rd_rdy),
    .Y(_006_[3])
  );
  \$_MUX_  _606_ (
    .A(xfer_buf[4]),
    .B(xfer_buf[5]),
    .S(_171_),
    .Y(_265_)
  );
  \$_MUX_  _607_ (
    .A(_265_),
    .B(dbg_dout[3]),
    .S(dbg_rd_rdy),
    .Y(_006_[4])
  );
  \$_MUX_  _608_ (
    .A(xfer_buf[5]),
    .B(xfer_buf[6]),
    .S(_171_),
    .Y(_266_)
  );
  \$_MUX_  _609_ (
    .A(_266_),
    .B(dbg_dout[4]),
    .S(dbg_rd_rdy),
    .Y(_006_[5])
  );
  \$_MUX_  _610_ (
    .A(xfer_buf[6]),
    .B(xfer_buf[7]),
    .S(_171_),
    .Y(_267_)
  );
  \$_MUX_  _611_ (
    .A(_267_),
    .B(dbg_dout[5]),
    .S(dbg_rd_rdy),
    .Y(_006_[6])
  );
  \$_MUX_  _612_ (
    .A(xfer_buf[7]),
    .B(xfer_buf[8]),
    .S(_171_),
    .Y(_268_)
  );
  \$_MUX_  _613_ (
    .A(_268_),
    .B(dbg_dout[6]),
    .S(dbg_rd_rdy),
    .Y(_006_[7])
  );
  \$_MUX_  _614_ (
    .A(xfer_buf[8]),
    .B(xfer_buf[9]),
    .S(_171_),
    .Y(_269_)
  );
  \$_MUX_  _615_ (
    .A(_269_),
    .B(dbg_dout[7]),
    .S(dbg_rd_rdy),
    .Y(_006_[8])
  );
  \$_MUX_  _616_ (
    .A(xfer_buf[9]),
    .B(xfer_buf[10]),
    .S(_171_),
    .Y(_270_)
  );
  \$_OR_  _617_ (
    .A(_270_),
    .B(dbg_rd_rdy),
    .Y(_006_[9])
  );
  \$_AND_  _618_ (
    .A(_171_),
    .B(_027_),
    .Y(_271_)
  );
  \$_MUX_  _619_ (
    .A(dbg_uart_txd),
    .B(xfer_buf[0]),
    .S(_271_),
    .Y(_002_)
  );
  \$_AND_  _620_ (
    .A(_025_),
    .B(uart_state[2]),
    .Y(_272_)
  );
  \$_MUX_  _621_ (
    .A(dbg_addr[0]),
    .B(xfer_buf[12]),
    .S(_272_),
    .Y(_000_[0])
  );
  \$_MUX_  _622_ (
    .A(dbg_addr[1]),
    .B(xfer_buf[13]),
    .S(_272_),
    .Y(_000_[1])
  );
  \$_MUX_  _623_ (
    .A(dbg_addr[2]),
    .B(xfer_buf[14]),
    .S(_272_),
    .Y(_000_[2])
  );
  \$_MUX_  _624_ (
    .A(dbg_addr[3]),
    .B(xfer_buf[15]),
    .S(_272_),
    .Y(_000_[3])
  );
  \$_MUX_  _625_ (
    .A(dbg_addr[4]),
    .B(xfer_buf[16]),
    .S(_272_),
    .Y(_000_[4])
  );
  \$_MUX_  _626_ (
    .A(dbg_addr[5]),
    .B(xfer_buf[17]),
    .S(_272_),
    .Y(_000_[5])
  );
  \$_MUX_  _627_ (
    .A(dbg_bw),
    .B(xfer_buf[18]),
    .S(_272_),
    .Y(_001_)
  );
  \$_MUX_  _628_ (
    .A(dbg_bw),
    .B(mem_bw),
    .S(mem_burst),
    .Y(_273_)
  );
  \$_MUX_  _629_ (
    .A(xfer_buf[3]),
    .B(xfer_buf[12]),
    .S(_273_),
    .Y(dbg_din[0])
  );
  \$_INV_  _630_ (
    .A(_273_),
    .Y(_274_)
  );
  \$_AND_  _631_ (
    .A(_274_),
    .B(xfer_buf[14]),
    .Y(dbg_din[10])
  );
  \$_AND_  _632_ (
    .A(_274_),
    .B(xfer_buf[15]),
    .Y(dbg_din[11])
  );
  \$_AND_  _633_ (
    .A(_274_),
    .B(xfer_buf[16]),
    .Y(dbg_din[12])
  );
  \$_AND_  _634_ (
    .A(_274_),
    .B(xfer_buf[17]),
    .Y(dbg_din[13])
  );
  \$_AND_  _635_ (
    .A(_274_),
    .B(xfer_buf[18]),
    .Y(dbg_din[14])
  );
  \$_AND_  _636_ (
    .A(_274_),
    .B(xfer_buf[19]),
    .Y(dbg_din[15])
  );
  \$_MUX_  _637_ (
    .A(xfer_buf[4]),
    .B(xfer_buf[13]),
    .S(_273_),
    .Y(dbg_din[1])
  );
  \$_MUX_  _638_ (
    .A(xfer_buf[5]),
    .B(xfer_buf[14]),
    .S(_273_),
    .Y(dbg_din[2])
  );
  \$_MUX_  _639_ (
    .A(xfer_buf[6]),
    .B(xfer_buf[15]),
    .S(_273_),
    .Y(dbg_din[3])
  );
  \$_MUX_  _640_ (
    .A(xfer_buf[7]),
    .B(xfer_buf[16]),
    .S(_273_),
    .Y(dbg_din[4])
  );
  \$_MUX_  _641_ (
    .A(xfer_buf[8]),
    .B(xfer_buf[17]),
    .S(_273_),
    .Y(dbg_din[5])
  );
  \$_MUX_  _642_ (
    .A(xfer_buf[9]),
    .B(xfer_buf[18]),
    .S(_273_),
    .Y(dbg_din[6])
  );
  \$_MUX_  _643_ (
    .A(xfer_buf[10]),
    .B(xfer_buf[19]),
    .S(_273_),
    .Y(dbg_din[7])
  );
  \$_AND_  _644_ (
    .A(_274_),
    .B(xfer_buf[12]),
    .Y(dbg_din[8])
  );
  \$_AND_  _645_ (
    .A(_274_),
    .B(xfer_buf[13]),
    .Y(dbg_din[9])
  );
  \$_AND_  _646_ (
    .A(uart_state[3]),
    .B(mem_burst),
    .Y(_275_)
  );
  \$_AND_  _647_ (
    .A(_275_),
    .B(_025_),
    .Y(_276_)
  );
  \$_AND_  _648_ (
    .A(_272_),
    .B(_047_),
    .Y(_277_)
  );
  \$_OR_  _649_ (
    .A(_277_),
    .B(mem_burst_rd),
    .Y(_278_)
  );
  \$_AND_  _650_ (
    .A(_278_),
    .B(_041_),
    .Y(_279_)
  );
  \$_OR_  _651_ (
    .A(_279_),
    .B(_276_),
    .Y(dbg_rd)
  );
  \$_DFF_PP0_  \uart_state_reg[0]  /* _652_ */ (
    .C(dbg_clk),
    .D(_280_),
    .Q(uart_state[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \uart_state_reg[1]  /* _653_ */ (
    .C(dbg_clk),
    .D(_281_),
    .Q(uart_state[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \uart_state_reg[2]  /* _654_ */ (
    .C(dbg_clk),
    .D(_282_),
    .Q(uart_state[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \uart_state_reg[3]  /* _655_ */ (
    .C(dbg_clk),
    .D(_283_),
    .Q(uart_state[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \uart_state_reg[4]  /* _656_ */ (
    .C(dbg_clk),
    .D(_284_),
    .Q(uart_state[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \rxd_buf_reg[0]  /* _657_ */ (
    .C(dbg_clk),
    .D(uart_rxd),
    .Q(rxd_buf[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \rxd_buf_reg[1]  /* _658_ */ (
    .C(dbg_clk),
    .D(rxd_buf[0]),
    .Q(rxd_buf[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  rxd_maj_reg /* _659_ */ (
    .C(dbg_clk),
    .D(rxd_maj_nxt),
    .Q(rxd_maj),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  sync_busy_reg /* _660_ */ (
    .C(dbg_clk),
    .D(_003_),
    .Q(sync_busy),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \sync_cnt_reg[0]  /* _661_ */ (
    .C(dbg_clk),
    .D(_004_[0]),
    .Q(sync_cnt[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[7]  /* _662_ */ (
    .C(dbg_clk),
    .D(_004_[10]),
    .Q(bit_cnt_max[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[8]  /* _663_ */ (
    .C(dbg_clk),
    .D(_004_[11]),
    .Q(bit_cnt_max[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[9]  /* _664_ */ (
    .C(dbg_clk),
    .D(_004_[12]),
    .Q(bit_cnt_max[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[10]  /* _665_ */ (
    .C(dbg_clk),
    .D(_004_[13]),
    .Q(bit_cnt_max[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[11]  /* _666_ */ (
    .C(dbg_clk),
    .D(_004_[14]),
    .Q(bit_cnt_max[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[12]  /* _667_ */ (
    .C(dbg_clk),
    .D(_004_[15]),
    .Q(bit_cnt_max[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[13]  /* _668_ */ (
    .C(dbg_clk),
    .D(_004_[16]),
    .Q(bit_cnt_max[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[14]  /* _669_ */ (
    .C(dbg_clk),
    .D(_004_[17]),
    .Q(bit_cnt_max[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[15]  /* _670_ */ (
    .C(dbg_clk),
    .D(_004_[18]),
    .Q(bit_cnt_max[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \sync_cnt_reg[1]  /* _671_ */ (
    .C(dbg_clk),
    .D(_004_[1]),
    .Q(sync_cnt[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \sync_cnt_reg[2]  /* _672_ */ (
    .C(dbg_clk),
    .D(_004_[2]),
    .Q(sync_cnt[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[0]  /* _673_ */ (
    .C(dbg_clk),
    .D(_004_[3]),
    .Q(bit_cnt_max[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[1]  /* _674_ */ (
    .C(dbg_clk),
    .D(_004_[4]),
    .Q(bit_cnt_max[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[2]  /* _675_ */ (
    .C(dbg_clk),
    .D(_004_[5]),
    .Q(bit_cnt_max[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[3]  /* _676_ */ (
    .C(dbg_clk),
    .D(_004_[6]),
    .Q(bit_cnt_max[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[4]  /* _677_ */ (
    .C(dbg_clk),
    .D(_004_[7]),
    .Q(bit_cnt_max[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[5]  /* _678_ */ (
    .C(dbg_clk),
    .D(_004_[8]),
    .Q(bit_cnt_max[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  \bit_cnt_max_reg[6]  /* _679_ */ (
    .C(dbg_clk),
    .D(_004_[9]),
    .Q(bit_cnt_max[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_bit_reg[0]  /* _680_ */ (
    .C(dbg_clk),
    .D(_005_[0]),
    .Q(xfer_bit[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_bit_reg[1]  /* _681_ */ (
    .C(dbg_clk),
    .D(_005_[1]),
    .Q(xfer_bit[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_bit_reg[2]  /* _682_ */ (
    .C(dbg_clk),
    .D(_005_[2]),
    .Q(xfer_bit[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_bit_reg[3]  /* _683_ */ (
    .C(dbg_clk),
    .D(_005_[3]),
    .Q(xfer_bit[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[0]  /* _684_ */ (
    .C(dbg_clk),
    .D(_007_[0]),
    .Q(xfer_cnt[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[10]  /* _685_ */ (
    .C(dbg_clk),
    .D(_007_[10]),
    .Q(xfer_cnt[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[11]  /* _686_ */ (
    .C(dbg_clk),
    .D(_007_[11]),
    .Q(xfer_cnt[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[12]  /* _687_ */ (
    .C(dbg_clk),
    .D(_007_[12]),
    .Q(xfer_cnt[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[13]  /* _688_ */ (
    .C(dbg_clk),
    .D(_007_[13]),
    .Q(xfer_cnt[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[14]  /* _689_ */ (
    .C(dbg_clk),
    .D(_007_[14]),
    .Q(xfer_cnt[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[15]  /* _690_ */ (
    .C(dbg_clk),
    .D(_007_[15]),
    .Q(xfer_cnt[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[1]  /* _691_ */ (
    .C(dbg_clk),
    .D(_007_[1]),
    .Q(xfer_cnt[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[2]  /* _692_ */ (
    .C(dbg_clk),
    .D(_007_[2]),
    .Q(xfer_cnt[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[3]  /* _693_ */ (
    .C(dbg_clk),
    .D(_007_[3]),
    .Q(xfer_cnt[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[4]  /* _694_ */ (
    .C(dbg_clk),
    .D(_007_[4]),
    .Q(xfer_cnt[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[5]  /* _695_ */ (
    .C(dbg_clk),
    .D(_007_[5]),
    .Q(xfer_cnt[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[6]  /* _696_ */ (
    .C(dbg_clk),
    .D(_007_[6]),
    .Q(xfer_cnt[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[7]  /* _697_ */ (
    .C(dbg_clk),
    .D(_007_[7]),
    .Q(xfer_cnt[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[8]  /* _698_ */ (
    .C(dbg_clk),
    .D(_007_[8]),
    .Q(xfer_cnt[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_cnt_reg[9]  /* _699_ */ (
    .C(dbg_clk),
    .D(_007_[9]),
    .Q(xfer_cnt[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[0]  /* _700_ */ (
    .C(dbg_clk),
    .D(_006_[0]),
    .Q(xfer_buf[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[10]  /* _701_ */ (
    .C(dbg_clk),
    .D(_006_[10]),
    .Q(xfer_buf[10]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[11]  /* _702_ */ (
    .C(dbg_clk),
    .D(_006_[11]),
    .Q(xfer_buf[11]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[12]  /* _703_ */ (
    .C(dbg_clk),
    .D(_006_[12]),
    .Q(xfer_buf[12]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[13]  /* _704_ */ (
    .C(dbg_clk),
    .D(_006_[13]),
    .Q(xfer_buf[13]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[14]  /* _705_ */ (
    .C(dbg_clk),
    .D(_006_[14]),
    .Q(xfer_buf[14]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[15]  /* _706_ */ (
    .C(dbg_clk),
    .D(_006_[15]),
    .Q(xfer_buf[15]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[16]  /* _707_ */ (
    .C(dbg_clk),
    .D(_006_[16]),
    .Q(xfer_buf[16]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[17]  /* _708_ */ (
    .C(dbg_clk),
    .D(_006_[17]),
    .Q(xfer_buf[17]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[18]  /* _709_ */ (
    .C(dbg_clk),
    .D(_006_[18]),
    .Q(xfer_buf[18]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[19]  /* _710_ */ (
    .C(dbg_clk),
    .D(_006_[19]),
    .Q(xfer_buf[19]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[1]  /* _711_ */ (
    .C(dbg_clk),
    .D(_006_[1]),
    .Q(xfer_buf[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[2]  /* _712_ */ (
    .C(dbg_clk),
    .D(_006_[2]),
    .Q(xfer_buf[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[3]  /* _713_ */ (
    .C(dbg_clk),
    .D(_006_[3]),
    .Q(xfer_buf[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[4]  /* _714_ */ (
    .C(dbg_clk),
    .D(_006_[4]),
    .Q(xfer_buf[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[5]  /* _715_ */ (
    .C(dbg_clk),
    .D(_006_[5]),
    .Q(xfer_buf[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[6]  /* _716_ */ (
    .C(dbg_clk),
    .D(_006_[6]),
    .Q(xfer_buf[6]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[7]  /* _717_ */ (
    .C(dbg_clk),
    .D(_006_[7]),
    .Q(xfer_buf[7]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[8]  /* _718_ */ (
    .C(dbg_clk),
    .D(_006_[8]),
    .Q(xfer_buf[8]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \xfer_buf_reg[9]  /* _719_ */ (
    .C(dbg_clk),
    .D(_006_[9]),
    .Q(xfer_buf[9]),
    .R(dbg_rst)
  );
  \$_DFF_PP1_  dbg_uart_txd_reg /* _720_ */ (
    .C(dbg_clk),
    .D(_002_),
    .Q(dbg_uart_txd),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[0]  /* _721_ */ (
    .C(dbg_clk),
    .D(_000_[0]),
    .Q(dbg_addr[0]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[1]  /* _722_ */ (
    .C(dbg_clk),
    .D(_000_[1]),
    .Q(dbg_addr[1]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[2]  /* _723_ */ (
    .C(dbg_clk),
    .D(_000_[2]),
    .Q(dbg_addr[2]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[3]  /* _724_ */ (
    .C(dbg_clk),
    .D(_000_[3]),
    .Q(dbg_addr[3]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[4]  /* _725_ */ (
    .C(dbg_clk),
    .D(_000_[4]),
    .Q(dbg_addr[4]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  \dbg_addr_reg[5]  /* _726_ */ (
    .C(dbg_clk),
    .D(_000_[5]),
    .Q(dbg_addr[5]),
    .R(dbg_rst)
  );
  \$_DFF_PP0_  dbg_bw_reg /* _727_ */ (
    .C(dbg_clk),
    .D(_001_),
    .Q(dbg_bw),
    .R(dbg_rst)
  );
  omsp_sync_cell sync_cell_uart_rxd (
    .clk(dbg_clk),
    .data_in(_285_),
    .data_out(uart_rxd_n),
    .rst(dbg_rst)
  );
  assign rxd_s = rxd_maj;
  assign sync_cnt[18:3] = bit_cnt_max;
  assign xfer_buf_nxt = { rxd_maj, xfer_buf[19:1] };
endmodule

module omsp_execution_unit(cpuoff, dbg_reg_din, gie, mab, mb_en, mb_wr, mdb_out, oscoff, pc_sw, pc_sw_wr, scg0, scg1, dbg_halt_st, dbg_mem_dout, dbg_reg_wr, e_state, exec_done, inst_ad, inst_as, inst_alu, inst_bw, inst_dest, inst_dext, inst_irq_rst, inst_jmp, inst_mov, inst_sext, inst_so, inst_src, inst_type, mclk, mdb_in, pc, pc_nxt, puc_rst, scan_enable);
  wire _000_;
  wire [15:0] _001_;
  wire _002_;
  wire _003_;
  wire [15:0] _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire [15:0] alu_out;
  wire [15:0] alu_out_add;
  wire [3:0] alu_stat;
  wire [3:0] alu_stat_wr;
  output cpuoff;
  input dbg_halt_st;
  input [15:0] dbg_mem_dout;
  output [15:0] dbg_reg_din;
  input dbg_reg_wr;
  input [3:0] e_state;
  wire exec_cycle;
  input exec_done;
  output gie;
  input [7:0] inst_ad;
  input [11:0] inst_alu;
  input [7:0] inst_as;
  input inst_bw;
  input [15:0] inst_dest;
  input [15:0] inst_dext;
  input inst_irq_rst;
  input [7:0] inst_jmp;
  input inst_mov;
  input [15:0] inst_sext;
  input [7:0] inst_so;
  input [15:0] inst_src;
  input [2:0] inst_type;
  output [15:0] mab;
  wire mab_lsb;
  output mb_en;
  output [1:0] mb_wr;
  input mclk;
  wire mclk_mdb_in_buf;
  wire mclk_mdb_out_nxt;
  input [15:0] mdb_in;
  wire [15:0] mdb_in_buf;
  wire mdb_in_buf_en;
  wire mdb_in_buf_valid;
  wire [15:0] mdb_in_bw;
  output [15:0] mdb_out;
  wire [15:0] mdb_out_nxt;
  wire [15:0] op_dst;
  wire [15:0] op_src;
  output oscoff;
  input [15:0] pc;
  input [15:0] pc_nxt;
  output [15:0] pc_sw;
  output pc_sw_wr;
  input puc_rst;
  wire [15:0] reg_dest;
  wire reg_dest_wr;
  wire reg_incr;
  wire reg_pc_call;
  wire reg_sp_wr;
  wire reg_sr_clr;
  wire reg_sr_wr;
  wire [15:0] reg_src;
  input scan_enable;
  output scg0;
  output scg1;
  wire [3:0] status;
  \$_INV_  _299_ (
    .A(e_state[2]),
    .Y(_005_)
  );
  \$_AND_  _300_ (
    .A(e_state[1]),
    .B(e_state[0]),
    .Y(_006_)
  );
  \$_AND_  _301_ (
    .A(_006_),
    .B(_005_),
    .Y(_007_)
  );
  \$_AND_  _302_ (
    .A(_007_),
    .B(e_state[3]),
    .Y(exec_cycle)
  );
  \$_INV_  _303_ (
    .A(e_state[0]),
    .Y(_008_)
  );
  \$_AND_  _304_ (
    .A(e_state[1]),
    .B(_008_),
    .Y(_009_)
  );
  \$_INV_  _305_ (
    .A(e_state[3]),
    .Y(_010_)
  );
  \$_AND_  _306_ (
    .A(_010_),
    .B(e_state[2]),
    .Y(_011_)
  );
  \$_AND_  _307_ (
    .A(_011_),
    .B(_009_),
    .Y(_002_)
  );
  \$_INV_  _308_ (
    .A(e_state[1]),
    .Y(_012_)
  );
  \$_AND_  _309_ (
    .A(_012_),
    .B(e_state[0]),
    .Y(_013_)
  );
  \$_AND_  _310_ (
    .A(_013_),
    .B(_005_),
    .Y(_014_)
  );
  \$_AND_  _311_ (
    .A(_014_),
    .B(e_state[3]),
    .Y(_015_)
  );
  \$_AND_  _312_ (
    .A(_015_),
    .B(inst_so[6]),
    .Y(reg_sr_wr)
  );
  \$_AND_  _313_ (
    .A(_014_),
    .B(_010_),
    .Y(_016_)
  );
  \$_AND_  _314_ (
    .A(_007_),
    .B(_010_),
    .Y(_017_)
  );
  \$_OR_  _315_ (
    .A(_017_),
    .B(_016_),
    .Y(_018_)
  );
  \$_AND_  _316_ (
    .A(_009_),
    .B(_005_),
    .Y(_019_)
  );
  \$_AND_  _317_ (
    .A(_019_),
    .B(e_state[3]),
    .Y(_020_)
  );
  \$_AND_  _318_ (
    .A(_011_),
    .B(_006_),
    .Y(_021_)
  );
  \$_OR_  _319_ (
    .A(_021_),
    .B(_020_),
    .Y(_022_)
  );
  \$_OR_  _320_ (
    .A(_022_),
    .B(_018_),
    .Y(_023_)
  );
  \$_INV_  _321_ (
    .A(inst_alu[11]),
    .Y(_024_)
  );
  \$_INV_  _322_ (
    .A(inst_bw),
    .Y(_025_)
  );
  \$_INV_  _323_ (
    .A(alu_out_add[0]),
    .Y(_026_)
  );
  \$_OR_  _324_ (
    .A(_026_),
    .B(_025_),
    .Y(_027_)
  );
  \$_AND_  _325_ (
    .A(_027_),
    .B(_024_),
    .Y(_028_)
  );
  \$_AND_  _326_ (
    .A(_028_),
    .B(_023_),
    .Y(mb_wr[0])
  );
  \$_OR_  _327_ (
    .A(alu_out_add[0]),
    .B(_025_),
    .Y(_029_)
  );
  \$_AND_  _328_ (
    .A(_029_),
    .B(_024_),
    .Y(_030_)
  );
  \$_AND_  _329_ (
    .A(_030_),
    .B(_023_),
    .Y(mb_wr[1])
  );
  \$_INV_  _330_ (
    .A(inst_so[6]),
    .Y(_031_)
  );
  \$_OR_  _331_ (
    .A(inst_so[4]),
    .B(inst_so[5]),
    .Y(_032_)
  );
  \$_INV_  _332_ (
    .A(_032_),
    .Y(_033_)
  );
  \$_AND_  _333_ (
    .A(_033_),
    .B(_031_),
    .Y(_034_)
  );
  \$_AND_  _334_ (
    .A(inst_type[0]),
    .B(inst_as[0]),
    .Y(_035_)
  );
  \$_AND_  _335_ (
    .A(_035_),
    .B(_034_),
    .Y(_036_)
  );
  \$_AND_  _336_ (
    .A(inst_type[2]),
    .B(inst_ad[0]),
    .Y(_037_)
  );
  \$_AND_  _337_ (
    .A(_037_),
    .B(_024_),
    .Y(_038_)
  );
  \$_OR_  _338_ (
    .A(_038_),
    .B(inst_type[1]),
    .Y(_039_)
  );
  \$_OR_  _339_ (
    .A(_039_),
    .B(_036_),
    .Y(_040_)
  );
  \$_AND_  _340_ (
    .A(_040_),
    .B(exec_cycle),
    .Y(_041_)
  );
  \$_OR_  _341_ (
    .A(_041_),
    .B(dbg_reg_wr),
    .Y(reg_dest_wr)
  );
  \$_INV_  _342_ (
    .A(inst_irq_rst),
    .Y(_042_)
  );
  \$_AND_  _343_ (
    .A(_018_),
    .B(_042_),
    .Y(_043_)
  );
  \$_OR_  _344_ (
    .A(inst_as[2]),
    .B(inst_as[3]),
    .Y(_044_)
  );
  \$_AND_  _345_ (
    .A(_044_),
    .B(inst_src[1]),
    .Y(_045_)
  );
  \$_AND_  _346_ (
    .A(_032_),
    .B(_002_),
    .Y(_046_)
  );
  \$_AND_  _347_ (
    .A(_046_),
    .B(_045_),
    .Y(_047_)
  );
  \$_INV_  _348_ (
    .A(_045_),
    .Y(_048_)
  );
  \$_INV_  _349_ (
    .A(inst_as[1]),
    .Y(_049_)
  );
  \$_AND_  _350_ (
    .A(_032_),
    .B(_049_),
    .Y(_050_)
  );
  \$_AND_  _351_ (
    .A(_050_),
    .B(_048_),
    .Y(_051_)
  );
  \$_AND_  _352_ (
    .A(_051_),
    .B(_015_),
    .Y(_052_)
  );
  \$_AND_  _353_ (
    .A(_013_),
    .B(_011_),
    .Y(_053_)
  );
  \$_AND_  _354_ (
    .A(_032_),
    .B(inst_as[1]),
    .Y(_054_)
  );
  \$_AND_  _355_ (
    .A(_054_),
    .B(_053_),
    .Y(_055_)
  );
  \$_OR_  _356_ (
    .A(_055_),
    .B(_052_),
    .Y(_056_)
  );
  \$_OR_  _357_ (
    .A(_056_),
    .B(_047_),
    .Y(_057_)
  );
  \$_OR_  _358_ (
    .A(_057_),
    .B(_043_),
    .Y(reg_sp_wr)
  );
  \$_AND_  _359_ (
    .A(exec_cycle),
    .B(inst_so[5]),
    .Y(_058_)
  );
  \$_OR_  _360_ (
    .A(_012_),
    .B(e_state[0]),
    .Y(_059_)
  );
  \$_OR_  _361_ (
    .A(_059_),
    .B(e_state[2]),
    .Y(_060_)
  );
  \$_OR_  _362_ (
    .A(_060_),
    .B(_010_),
    .Y(_061_)
  );
  \$_OR_  _363_ (
    .A(_061_),
    .B(_031_),
    .Y(_062_)
  );
  \$_INV_  _364_ (
    .A(_062_),
    .Y(_063_)
  );
  \$_OR_  _365_ (
    .A(_063_),
    .B(_058_),
    .Y(reg_pc_call)
  );
  \$_AND_  _366_ (
    .A(exec_cycle),
    .B(inst_so[6]),
    .Y(_064_)
  );
  \$_AND_  _367_ (
    .A(exec_done),
    .B(inst_as[3]),
    .Y(_065_)
  );
  \$_AND_  _368_ (
    .A(_002_),
    .B(inst_so[6]),
    .Y(_066_)
  );
  \$_OR_  _369_ (
    .A(_066_),
    .B(_065_),
    .Y(_067_)
  );
  \$_OR_  _370_ (
    .A(_067_),
    .B(_064_),
    .Y(reg_incr)
  );
  \$_AND_  _371_ (
    .A(_008_),
    .B(_005_),
    .Y(_068_)
  );
  \$_AND_  _372_ (
    .A(_010_),
    .B(_012_),
    .Y(_069_)
  );
  \$_AND_  _373_ (
    .A(_069_),
    .B(_068_),
    .Y(reg_sr_clr)
  );
  \$_INV_  _374_ (
    .A(inst_as[5]),
    .Y(_070_)
  );
  \$_AND_  _375_ (
    .A(_002_),
    .B(_070_),
    .Y(_071_)
  );
  \$_OR_  _376_ (
    .A(_071_),
    .B(_022_),
    .Y(_072_)
  );
  \$_AND_  _377_ (
    .A(_016_),
    .B(_042_),
    .Y(_073_)
  );
  \$_OR_  _378_ (
    .A(_073_),
    .B(_064_),
    .Y(_074_)
  );
  \$_AND_  _379_ (
    .A(_017_),
    .B(_042_),
    .Y(_075_)
  );
  \$_INV_  _380_ (
    .A(inst_type[0]),
    .Y(_076_)
  );
  \$_INV_  _381_ (
    .A(inst_mov),
    .Y(_077_)
  );
  \$_AND_  _382_ (
    .A(_077_),
    .B(_076_),
    .Y(_078_)
  );
  \$_AND_  _383_ (
    .A(_078_),
    .B(_015_),
    .Y(_079_)
  );
  \$_OR_  _384_ (
    .A(_079_),
    .B(_075_),
    .Y(_080_)
  );
  \$_OR_  _385_ (
    .A(_080_),
    .B(_074_),
    .Y(_081_)
  );
  \$_OR_  _386_ (
    .A(_081_),
    .B(_072_),
    .Y(mb_en)
  );
  \$_INV_  _387_ (
    .A(inst_so[5]),
    .Y(_082_)
  );
  \$_AND_  _388_ (
    .A(exec_cycle),
    .B(_082_),
    .Y(_083_)
  );
  \$_AND_  _389_ (
    .A(_019_),
    .B(_010_),
    .Y(_084_)
  );
  \$_OR_  _390_ (
    .A(_084_),
    .B(reg_sr_clr),
    .Y(_085_)
  );
  \$_OR_  _391_ (
    .A(_085_),
    .B(_083_),
    .Y(_086_)
  );
  \$_MUX_  _392_ (
    .A(mdb_out[0]),
    .B(alu_out[0]),
    .S(_086_),
    .Y(_087_)
  );
  \$_MUX_  _393_ (
    .A(_087_),
    .B(pc_nxt[0]),
    .S(_015_),
    .Y(_004_[0])
  );
  \$_MUX_  _394_ (
    .A(mdb_out_nxt[10]),
    .B(alu_out[10]),
    .S(_086_),
    .Y(_088_)
  );
  \$_MUX_  _395_ (
    .A(_088_),
    .B(pc_nxt[10]),
    .S(_015_),
    .Y(_004_[10])
  );
  \$_MUX_  _396_ (
    .A(mdb_out_nxt[11]),
    .B(alu_out[11]),
    .S(_086_),
    .Y(_089_)
  );
  \$_MUX_  _397_ (
    .A(_089_),
    .B(pc_nxt[11]),
    .S(_015_),
    .Y(_004_[11])
  );
  \$_MUX_  _398_ (
    .A(mdb_out_nxt[12]),
    .B(alu_out[12]),
    .S(_086_),
    .Y(_090_)
  );
  \$_MUX_  _399_ (
    .A(_090_),
    .B(pc_nxt[12]),
    .S(_015_),
    .Y(_004_[12])
  );
  \$_MUX_  _400_ (
    .A(mdb_out_nxt[13]),
    .B(alu_out[13]),
    .S(_086_),
    .Y(_091_)
  );
  \$_MUX_  _401_ (
    .A(_091_),
    .B(pc_nxt[13]),
    .S(_015_),
    .Y(_004_[13])
  );
  \$_MUX_  _402_ (
    .A(mdb_out_nxt[14]),
    .B(alu_out[14]),
    .S(_086_),
    .Y(_092_)
  );
  \$_MUX_  _403_ (
    .A(_092_),
    .B(pc_nxt[14]),
    .S(_015_),
    .Y(_004_[14])
  );
  \$_MUX_  _404_ (
    .A(mdb_out_nxt[15]),
    .B(alu_out[15]),
    .S(_086_),
    .Y(_093_)
  );
  \$_MUX_  _405_ (
    .A(_093_),
    .B(pc_nxt[15]),
    .S(_015_),
    .Y(_004_[15])
  );
  \$_MUX_  _406_ (
    .A(mdb_out[1]),
    .B(alu_out[1]),
    .S(_086_),
    .Y(_094_)
  );
  \$_MUX_  _407_ (
    .A(_094_),
    .B(pc_nxt[1]),
    .S(_015_),
    .Y(_004_[1])
  );
  \$_MUX_  _408_ (
    .A(mdb_out[2]),
    .B(alu_out[2]),
    .S(_086_),
    .Y(_095_)
  );
  \$_MUX_  _409_ (
    .A(_095_),
    .B(pc_nxt[2]),
    .S(_015_),
    .Y(_004_[2])
  );
  \$_MUX_  _410_ (
    .A(mdb_out[3]),
    .B(alu_out[3]),
    .S(_086_),
    .Y(_096_)
  );
  \$_MUX_  _411_ (
    .A(_096_),
    .B(pc_nxt[3]),
    .S(_015_),
    .Y(_004_[3])
  );
  \$_MUX_  _412_ (
    .A(mdb_out[4]),
    .B(alu_out[4]),
    .S(_086_),
    .Y(_097_)
  );
  \$_MUX_  _413_ (
    .A(_097_),
    .B(pc_nxt[4]),
    .S(_015_),
    .Y(_004_[4])
  );
  \$_MUX_  _414_ (
    .A(mdb_out[5]),
    .B(alu_out[5]),
    .S(_086_),
    .Y(_098_)
  );
  \$_MUX_  _415_ (
    .A(_098_),
    .B(pc_nxt[5]),
    .S(_015_),
    .Y(_004_[5])
  );
  \$_MUX_  _416_ (
    .A(mdb_out[6]),
    .B(alu_out[6]),
    .S(_086_),
    .Y(_099_)
  );
  \$_MUX_  _417_ (
    .A(_099_),
    .B(pc_nxt[6]),
    .S(_015_),
    .Y(_004_[6])
  );
  \$_MUX_  _418_ (
    .A(mdb_out[7]),
    .B(alu_out[7]),
    .S(_086_),
    .Y(_100_)
  );
  \$_MUX_  _419_ (
    .A(_100_),
    .B(pc_nxt[7]),
    .S(_015_),
    .Y(_004_[7])
  );
  \$_MUX_  _420_ (
    .A(mdb_out_nxt[8]),
    .B(alu_out[8]),
    .S(_086_),
    .Y(_101_)
  );
  \$_MUX_  _421_ (
    .A(_101_),
    .B(pc_nxt[8]),
    .S(_015_),
    .Y(_004_[8])
  );
  \$_MUX_  _422_ (
    .A(mdb_out_nxt[9]),
    .B(alu_out[9]),
    .S(_086_),
    .Y(_102_)
  );
  \$_MUX_  _423_ (
    .A(_102_),
    .B(pc_nxt[9]),
    .S(_015_),
    .Y(_004_[9])
  );
  \$_MUX_  _424_ (
    .A(mab_lsb),
    .B(alu_out_add[0]),
    .S(mb_en),
    .Y(_000_)
  );
  \$_INV_  _425_ (
    .A(exec_cycle),
    .Y(_103_)
  );
  \$_OR_  _426_ (
    .A(mdb_in_buf_valid),
    .B(mdb_in_buf_en),
    .Y(_104_)
  );
  \$_AND_  _427_ (
    .A(_104_),
    .B(_103_),
    .Y(_003_)
  );
  \$_INV_  _428_ (
    .A(mdb_in_buf_en),
    .Y(_105_)
  );
  \$_MUX_  _429_ (
    .A(mdb_in[0]),
    .B(mdb_in[8]),
    .S(mab_lsb),
    .Y(_106_)
  );
  \$_MUX_  _430_ (
    .A(_106_),
    .B(mdb_in[0]),
    .S(_025_),
    .Y(_107_)
  );
  \$_MUX_  _431_ (
    .A(_107_),
    .B(mdb_in_buf[0]),
    .S(_105_),
    .Y(_001_[0])
  );
  \$_MUX_  _432_ (
    .A(mdb_in_buf[10]),
    .B(mdb_in[10]),
    .S(mdb_in_buf_en),
    .Y(_001_[10])
  );
  \$_MUX_  _433_ (
    .A(mdb_in_buf[11]),
    .B(mdb_in[11]),
    .S(mdb_in_buf_en),
    .Y(_001_[11])
  );
  \$_MUX_  _434_ (
    .A(mdb_in_buf[12]),
    .B(mdb_in[12]),
    .S(mdb_in_buf_en),
    .Y(_001_[12])
  );
  \$_MUX_  _435_ (
    .A(mdb_in_buf[13]),
    .B(mdb_in[13]),
    .S(mdb_in_buf_en),
    .Y(_001_[13])
  );
  \$_MUX_  _436_ (
    .A(mdb_in_buf[14]),
    .B(mdb_in[14]),
    .S(mdb_in_buf_en),
    .Y(_001_[14])
  );
  \$_MUX_  _437_ (
    .A(mdb_in_buf[15]),
    .B(mdb_in[15]),
    .S(mdb_in_buf_en),
    .Y(_001_[15])
  );
  \$_MUX_  _438_ (
    .A(mdb_in[1]),
    .B(mdb_in[9]),
    .S(mab_lsb),
    .Y(_108_)
  );
  \$_MUX_  _439_ (
    .A(_108_),
    .B(mdb_in[1]),
    .S(_025_),
    .Y(_109_)
  );
  \$_MUX_  _440_ (
    .A(_109_),
    .B(mdb_in_buf[1]),
    .S(_105_),
    .Y(_001_[1])
  );
  \$_MUX_  _441_ (
    .A(mdb_in[2]),
    .B(mdb_in[10]),
    .S(mab_lsb),
    .Y(_110_)
  );
  \$_MUX_  _442_ (
    .A(_110_),
    .B(mdb_in[2]),
    .S(_025_),
    .Y(_111_)
  );
  \$_MUX_  _443_ (
    .A(_111_),
    .B(mdb_in_buf[2]),
    .S(_105_),
    .Y(_001_[2])
  );
  \$_MUX_  _444_ (
    .A(mdb_in[3]),
    .B(mdb_in[11]),
    .S(mab_lsb),
    .Y(_112_)
  );
  \$_MUX_  _445_ (
    .A(_112_),
    .B(mdb_in[3]),
    .S(_025_),
    .Y(_113_)
  );
  \$_MUX_  _446_ (
    .A(_113_),
    .B(mdb_in_buf[3]),
    .S(_105_),
    .Y(_001_[3])
  );
  \$_MUX_  _447_ (
    .A(mdb_in[4]),
    .B(mdb_in[12]),
    .S(mab_lsb),
    .Y(_114_)
  );
  \$_MUX_  _448_ (
    .A(_114_),
    .B(mdb_in[4]),
    .S(_025_),
    .Y(_115_)
  );
  \$_MUX_  _449_ (
    .A(_115_),
    .B(mdb_in_buf[4]),
    .S(_105_),
    .Y(_001_[4])
  );
  \$_MUX_  _450_ (
    .A(mdb_in[5]),
    .B(mdb_in[13]),
    .S(mab_lsb),
    .Y(_116_)
  );
  \$_MUX_  _451_ (
    .A(_116_),
    .B(mdb_in[5]),
    .S(_025_),
    .Y(_117_)
  );
  \$_MUX_  _452_ (
    .A(_117_),
    .B(mdb_in_buf[5]),
    .S(_105_),
    .Y(_001_[5])
  );
  \$_MUX_  _453_ (
    .A(mdb_in[6]),
    .B(mdb_in[14]),
    .S(mab_lsb),
    .Y(_118_)
  );
  \$_MUX_  _454_ (
    .A(_118_),
    .B(mdb_in[6]),
    .S(_025_),
    .Y(_119_)
  );
  \$_MUX_  _455_ (
    .A(_119_),
    .B(mdb_in_buf[6]),
    .S(_105_),
    .Y(_001_[6])
  );
  \$_MUX_  _456_ (
    .A(mdb_in[7]),
    .B(mdb_in[15]),
    .S(mab_lsb),
    .Y(_120_)
  );
  \$_MUX_  _457_ (
    .A(_120_),
    .B(mdb_in[7]),
    .S(_025_),
    .Y(_121_)
  );
  \$_MUX_  _458_ (
    .A(_121_),
    .B(mdb_in_buf[7]),
    .S(_105_),
    .Y(_001_[7])
  );
  \$_MUX_  _459_ (
    .A(mdb_in_buf[8]),
    .B(mdb_in[8]),
    .S(mdb_in_buf_en),
    .Y(_001_[8])
  );
  \$_MUX_  _460_ (
    .A(mdb_in_buf[9]),
    .B(mdb_in[9]),
    .S(mdb_in_buf_en),
    .Y(_001_[9])
  );
  \$_INV_  _461_ (
    .A(inst_type[1]),
    .Y(_122_)
  );
  \$_AND_  _462_ (
    .A(_122_),
    .B(inst_as[0]),
    .Y(_123_)
  );
  \$_AND_  _463_ (
    .A(_123_),
    .B(exec_cycle),
    .Y(_124_)
  );
  \$_INV_  _464_ (
    .A(inst_as[6]),
    .Y(_125_)
  );
  \$_AND_  _465_ (
    .A(_002_),
    .B(_125_),
    .Y(_126_)
  );
  \$_AND_  _466_ (
    .A(_021_),
    .B(_125_),
    .Y(_127_)
  );
  \$_OR_  _467_ (
    .A(_127_),
    .B(_126_),
    .Y(_128_)
  );
  \$_OR_  _468_ (
    .A(_128_),
    .B(_085_),
    .Y(_129_)
  );
  \$_OR_  _469_ (
    .A(_129_),
    .B(_124_),
    .Y(_130_)
  );
  \$_AND_  _470_ (
    .A(_032_),
    .B(_015_),
    .Y(_131_)
  );
  \$_OR_  _471_ (
    .A(_055_),
    .B(_018_),
    .Y(_132_)
  );
  \$_OR_  _472_ (
    .A(_132_),
    .B(_131_),
    .Y(_133_)
  );
  \$_OR_  _473_ (
    .A(inst_as[6]),
    .B(inst_as[1]),
    .Y(_134_)
  );
  \$_OR_  _474_ (
    .A(_134_),
    .B(inst_as[4]),
    .Y(_135_)
  );
  \$_OR_  _475_ (
    .A(_135_),
    .B(_044_),
    .Y(_136_)
  );
  \$_AND_  _476_ (
    .A(_136_),
    .B(exec_cycle),
    .Y(_137_)
  );
  \$_OR_  _477_ (
    .A(_137_),
    .B(reg_sr_wr),
    .Y(_138_)
  );
  \$_MUX_  _478_ (
    .A(_107_),
    .B(mdb_in_buf[0]),
    .S(mdb_in_buf_valid),
    .Y(_139_)
  );
  \$_AND_  _479_ (
    .A(_033_),
    .B(_015_),
    .Y(_140_)
  );
  \$_AND_  _480_ (
    .A(_034_),
    .B(_020_),
    .Y(_141_)
  );
  \$_OR_  _481_ (
    .A(_141_),
    .B(_140_),
    .Y(_142_)
  );
  \$_OR_  _482_ (
    .A(inst_type[1]),
    .B(inst_so[6]),
    .Y(_143_)
  );
  \$_OR_  _483_ (
    .A(inst_as[7]),
    .B(inst_as[5]),
    .Y(_144_)
  );
  \$_OR_  _484_ (
    .A(_144_),
    .B(_143_),
    .Y(_145_)
  );
  \$_AND_  _485_ (
    .A(_145_),
    .B(exec_cycle),
    .Y(_146_)
  );
  \$_AND_  _486_ (
    .A(_146_),
    .B(inst_sext[0]),
    .Y(_147_)
  );
  \$_MUX_  _487_ (
    .A(_147_),
    .B(inst_dext[0]),
    .S(_142_),
    .Y(_148_)
  );
  \$_MUX_  _488_ (
    .A(_148_),
    .B(_139_),
    .S(_138_),
    .Y(_149_)
  );
  \$_MUX_  _489_ (
    .A(_149_),
    .B(dbg_reg_din[0]),
    .S(_133_),
    .Y(_150_)
  );
  \$_MUX_  _490_ (
    .A(_150_),
    .B(reg_src[0]),
    .S(_130_),
    .Y(op_src[0])
  );
  \$_MUX_  _491_ (
    .A(mdb_in[10]),
    .B(mdb_in_buf[10]),
    .S(mdb_in_buf_valid),
    .Y(_151_)
  );
  \$_AND_  _492_ (
    .A(_146_),
    .B(inst_sext[10]),
    .Y(_152_)
  );
  \$_MUX_  _493_ (
    .A(_152_),
    .B(inst_dext[10]),
    .S(_142_),
    .Y(_153_)
  );
  \$_MUX_  _494_ (
    .A(_153_),
    .B(_151_),
    .S(_138_),
    .Y(_154_)
  );
  \$_MUX_  _495_ (
    .A(_154_),
    .B(dbg_reg_din[10]),
    .S(_133_),
    .Y(_155_)
  );
  \$_MUX_  _496_ (
    .A(_155_),
    .B(reg_src[10]),
    .S(_130_),
    .Y(op_src[10])
  );
  \$_MUX_  _497_ (
    .A(mdb_in[11]),
    .B(mdb_in_buf[11]),
    .S(mdb_in_buf_valid),
    .Y(_156_)
  );
  \$_AND_  _498_ (
    .A(_146_),
    .B(inst_sext[11]),
    .Y(_157_)
  );
  \$_MUX_  _499_ (
    .A(_157_),
    .B(inst_dext[11]),
    .S(_142_),
    .Y(_158_)
  );
  \$_MUX_  _500_ (
    .A(_158_),
    .B(_156_),
    .S(_138_),
    .Y(_159_)
  );
  \$_MUX_  _501_ (
    .A(_159_),
    .B(dbg_reg_din[11]),
    .S(_133_),
    .Y(_160_)
  );
  \$_MUX_  _502_ (
    .A(_160_),
    .B(reg_src[11]),
    .S(_130_),
    .Y(op_src[11])
  );
  \$_MUX_  _503_ (
    .A(mdb_in[12]),
    .B(mdb_in_buf[12]),
    .S(mdb_in_buf_valid),
    .Y(_161_)
  );
  \$_AND_  _504_ (
    .A(_146_),
    .B(inst_sext[12]),
    .Y(_162_)
  );
  \$_MUX_  _505_ (
    .A(_162_),
    .B(inst_dext[12]),
    .S(_142_),
    .Y(_163_)
  );
  \$_MUX_  _506_ (
    .A(_163_),
    .B(_161_),
    .S(_138_),
    .Y(_164_)
  );
  \$_MUX_  _507_ (
    .A(_164_),
    .B(dbg_reg_din[12]),
    .S(_133_),
    .Y(_165_)
  );
  \$_MUX_  _508_ (
    .A(_165_),
    .B(reg_src[12]),
    .S(_130_),
    .Y(op_src[12])
  );
  \$_MUX_  _509_ (
    .A(mdb_in[13]),
    .B(mdb_in_buf[13]),
    .S(mdb_in_buf_valid),
    .Y(_166_)
  );
  \$_AND_  _510_ (
    .A(_146_),
    .B(inst_sext[13]),
    .Y(_167_)
  );
  \$_MUX_  _511_ (
    .A(_167_),
    .B(inst_dext[13]),
    .S(_142_),
    .Y(_168_)
  );
  \$_MUX_  _512_ (
    .A(_168_),
    .B(_166_),
    .S(_138_),
    .Y(_169_)
  );
  \$_MUX_  _513_ (
    .A(_169_),
    .B(dbg_reg_din[13]),
    .S(_133_),
    .Y(_170_)
  );
  \$_MUX_  _514_ (
    .A(_170_),
    .B(reg_src[13]),
    .S(_130_),
    .Y(op_src[13])
  );
  \$_MUX_  _515_ (
    .A(mdb_in[14]),
    .B(mdb_in_buf[14]),
    .S(mdb_in_buf_valid),
    .Y(_171_)
  );
  \$_AND_  _516_ (
    .A(_146_),
    .B(inst_sext[14]),
    .Y(_172_)
  );
  \$_MUX_  _517_ (
    .A(_172_),
    .B(inst_dext[14]),
    .S(_142_),
    .Y(_173_)
  );
  \$_MUX_  _518_ (
    .A(_173_),
    .B(_171_),
    .S(_138_),
    .Y(_174_)
  );
  \$_MUX_  _519_ (
    .A(_174_),
    .B(dbg_reg_din[14]),
    .S(_133_),
    .Y(_175_)
  );
  \$_MUX_  _520_ (
    .A(_175_),
    .B(reg_src[14]),
    .S(_130_),
    .Y(op_src[14])
  );
  \$_MUX_  _521_ (
    .A(mdb_in[15]),
    .B(mdb_in_buf[15]),
    .S(mdb_in_buf_valid),
    .Y(_176_)
  );
  \$_AND_  _522_ (
    .A(_146_),
    .B(inst_sext[15]),
    .Y(_177_)
  );
  \$_MUX_  _523_ (
    .A(_177_),
    .B(inst_dext[15]),
    .S(_142_),
    .Y(_178_)
  );
  \$_MUX_  _524_ (
    .A(_178_),
    .B(_176_),
    .S(_138_),
    .Y(_179_)
  );
  \$_MUX_  _525_ (
    .A(_179_),
    .B(dbg_reg_din[15]),
    .S(_133_),
    .Y(_180_)
  );
  \$_MUX_  _526_ (
    .A(_180_),
    .B(reg_src[15]),
    .S(_130_),
    .Y(op_src[15])
  );
  \$_MUX_  _527_ (
    .A(_109_),
    .B(mdb_in_buf[1]),
    .S(mdb_in_buf_valid),
    .Y(_181_)
  );
  \$_AND_  _528_ (
    .A(_146_),
    .B(inst_sext[1]),
    .Y(_182_)
  );
  \$_MUX_  _529_ (
    .A(_182_),
    .B(inst_dext[1]),
    .S(_142_),
    .Y(_183_)
  );
  \$_MUX_  _530_ (
    .A(_183_),
    .B(_181_),
    .S(_138_),
    .Y(_184_)
  );
  \$_MUX_  _531_ (
    .A(_184_),
    .B(dbg_reg_din[1]),
    .S(_133_),
    .Y(_185_)
  );
  \$_MUX_  _532_ (
    .A(_185_),
    .B(reg_src[1]),
    .S(_130_),
    .Y(op_src[1])
  );
  \$_MUX_  _533_ (
    .A(_111_),
    .B(mdb_in_buf[2]),
    .S(mdb_in_buf_valid),
    .Y(_186_)
  );
  \$_AND_  _534_ (
    .A(_146_),
    .B(inst_sext[2]),
    .Y(_187_)
  );
  \$_MUX_  _535_ (
    .A(_187_),
    .B(inst_dext[2]),
    .S(_142_),
    .Y(_188_)
  );
  \$_MUX_  _536_ (
    .A(_188_),
    .B(_186_),
    .S(_138_),
    .Y(_189_)
  );
  \$_MUX_  _537_ (
    .A(_189_),
    .B(dbg_reg_din[2]),
    .S(_133_),
    .Y(_190_)
  );
  \$_MUX_  _538_ (
    .A(_190_),
    .B(reg_src[2]),
    .S(_130_),
    .Y(op_src[2])
  );
  \$_MUX_  _539_ (
    .A(_113_),
    .B(mdb_in_buf[3]),
    .S(mdb_in_buf_valid),
    .Y(_191_)
  );
  \$_AND_  _540_ (
    .A(_146_),
    .B(inst_sext[3]),
    .Y(_192_)
  );
  \$_MUX_  _541_ (
    .A(_192_),
    .B(inst_dext[3]),
    .S(_142_),
    .Y(_193_)
  );
  \$_MUX_  _542_ (
    .A(_193_),
    .B(_191_),
    .S(_138_),
    .Y(_194_)
  );
  \$_MUX_  _543_ (
    .A(_194_),
    .B(dbg_reg_din[3]),
    .S(_133_),
    .Y(_195_)
  );
  \$_MUX_  _544_ (
    .A(_195_),
    .B(reg_src[3]),
    .S(_130_),
    .Y(op_src[3])
  );
  \$_MUX_  _545_ (
    .A(_115_),
    .B(mdb_in_buf[4]),
    .S(mdb_in_buf_valid),
    .Y(_196_)
  );
  \$_AND_  _546_ (
    .A(_146_),
    .B(inst_sext[4]),
    .Y(_197_)
  );
  \$_MUX_  _547_ (
    .A(_197_),
    .B(inst_dext[4]),
    .S(_142_),
    .Y(_198_)
  );
  \$_MUX_  _548_ (
    .A(_198_),
    .B(_196_),
    .S(_138_),
    .Y(_199_)
  );
  \$_MUX_  _549_ (
    .A(_199_),
    .B(dbg_reg_din[4]),
    .S(_133_),
    .Y(_200_)
  );
  \$_MUX_  _550_ (
    .A(_200_),
    .B(reg_src[4]),
    .S(_130_),
    .Y(op_src[4])
  );
  \$_MUX_  _551_ (
    .A(_117_),
    .B(mdb_in_buf[5]),
    .S(mdb_in_buf_valid),
    .Y(_201_)
  );
  \$_AND_  _552_ (
    .A(_146_),
    .B(inst_sext[5]),
    .Y(_202_)
  );
  \$_MUX_  _553_ (
    .A(_202_),
    .B(inst_dext[5]),
    .S(_142_),
    .Y(_203_)
  );
  \$_MUX_  _554_ (
    .A(_203_),
    .B(_201_),
    .S(_138_),
    .Y(_204_)
  );
  \$_MUX_  _555_ (
    .A(_204_),
    .B(dbg_reg_din[5]),
    .S(_133_),
    .Y(_205_)
  );
  \$_MUX_  _556_ (
    .A(_205_),
    .B(reg_src[5]),
    .S(_130_),
    .Y(op_src[5])
  );
  \$_MUX_  _557_ (
    .A(_119_),
    .B(mdb_in_buf[6]),
    .S(mdb_in_buf_valid),
    .Y(_206_)
  );
  \$_AND_  _558_ (
    .A(_146_),
    .B(inst_sext[6]),
    .Y(_207_)
  );
  \$_MUX_  _559_ (
    .A(_207_),
    .B(inst_dext[6]),
    .S(_142_),
    .Y(_208_)
  );
  \$_MUX_  _560_ (
    .A(_208_),
    .B(_206_),
    .S(_138_),
    .Y(_209_)
  );
  \$_MUX_  _561_ (
    .A(_209_),
    .B(dbg_reg_din[6]),
    .S(_133_),
    .Y(_210_)
  );
  \$_MUX_  _562_ (
    .A(_210_),
    .B(reg_src[6]),
    .S(_130_),
    .Y(op_src[6])
  );
  \$_MUX_  _563_ (
    .A(_121_),
    .B(mdb_in_buf[7]),
    .S(mdb_in_buf_valid),
    .Y(_211_)
  );
  \$_AND_  _564_ (
    .A(_146_),
    .B(inst_sext[7]),
    .Y(_212_)
  );
  \$_MUX_  _565_ (
    .A(_212_),
    .B(inst_dext[7]),
    .S(_142_),
    .Y(_213_)
  );
  \$_MUX_  _566_ (
    .A(_213_),
    .B(_211_),
    .S(_138_),
    .Y(_214_)
  );
  \$_MUX_  _567_ (
    .A(_214_),
    .B(dbg_reg_din[7]),
    .S(_133_),
    .Y(_215_)
  );
  \$_MUX_  _568_ (
    .A(_215_),
    .B(reg_src[7]),
    .S(_130_),
    .Y(op_src[7])
  );
  \$_MUX_  _569_ (
    .A(mdb_in[8]),
    .B(mdb_in_buf[8]),
    .S(mdb_in_buf_valid),
    .Y(_216_)
  );
  \$_AND_  _570_ (
    .A(_146_),
    .B(inst_sext[8]),
    .Y(_217_)
  );
  \$_MUX_  _571_ (
    .A(_217_),
    .B(inst_dext[8]),
    .S(_142_),
    .Y(_218_)
  );
  \$_MUX_  _572_ (
    .A(_218_),
    .B(_216_),
    .S(_138_),
    .Y(_219_)
  );
  \$_MUX_  _573_ (
    .A(_219_),
    .B(dbg_reg_din[8]),
    .S(_133_),
    .Y(_220_)
  );
  \$_MUX_  _574_ (
    .A(_220_),
    .B(reg_src[8]),
    .S(_130_),
    .Y(op_src[8])
  );
  \$_MUX_  _575_ (
    .A(mdb_in[9]),
    .B(mdb_in_buf[9]),
    .S(mdb_in_buf_valid),
    .Y(_221_)
  );
  \$_AND_  _576_ (
    .A(_146_),
    .B(inst_sext[9]),
    .Y(_222_)
  );
  \$_MUX_  _577_ (
    .A(_222_),
    .B(inst_dext[9]),
    .S(_142_),
    .Y(_223_)
  );
  \$_MUX_  _578_ (
    .A(_223_),
    .B(_221_),
    .S(_138_),
    .Y(_224_)
  );
  \$_MUX_  _579_ (
    .A(_224_),
    .B(dbg_reg_din[9]),
    .S(_133_),
    .Y(_225_)
  );
  \$_MUX_  _580_ (
    .A(_225_),
    .B(reg_src[9]),
    .S(_130_),
    .Y(op_src[9])
  );
  \$_AND_  _581_ (
    .A(_135_),
    .B(_002_),
    .Y(_226_)
  );
  \$_AND_  _582_ (
    .A(_135_),
    .B(_021_),
    .Y(_227_)
  );
  \$_OR_  _583_ (
    .A(_227_),
    .B(_226_),
    .Y(_228_)
  );
  \$_OR_  _584_ (
    .A(inst_type[0]),
    .B(inst_ad[0]),
    .Y(_229_)
  );
  \$_OR_  _585_ (
    .A(_229_),
    .B(inst_type[1]),
    .Y(_230_)
  );
  \$_OR_  _586_ (
    .A(_230_),
    .B(inst_so[6]),
    .Y(_231_)
  );
  \$_OR_  _587_ (
    .A(_231_),
    .B(_103_),
    .Y(_232_)
  );
  \$_AND_  _588_ (
    .A(_232_),
    .B(_062_),
    .Y(_233_)
  );
  \$_INV_  _589_ (
    .A(_233_),
    .Y(_234_)
  );
  \$_AND_  _590_ (
    .A(_234_),
    .B(_107_),
    .Y(_235_)
  );
  \$_AND_  _591_ (
    .A(_230_),
    .B(_031_),
    .Y(_236_)
  );
  \$_AND_  _592_ (
    .A(_236_),
    .B(exec_cycle),
    .Y(_237_)
  );
  \$_INV_  _593_ (
    .A(inst_ad[6]),
    .Y(_238_)
  );
  \$_AND_  _594_ (
    .A(_238_),
    .B(_031_),
    .Y(_239_)
  );
  \$_AND_  _595_ (
    .A(_239_),
    .B(_033_),
    .Y(_240_)
  );
  \$_AND_  _596_ (
    .A(_240_),
    .B(_015_),
    .Y(_241_)
  );
  \$_AND_  _597_ (
    .A(_020_),
    .B(_238_),
    .Y(_242_)
  );
  \$_OR_  _598_ (
    .A(_242_),
    .B(_241_),
    .Y(_243_)
  );
  \$_OR_  _599_ (
    .A(_243_),
    .B(_237_),
    .Y(_244_)
  );
  \$_AND_  _600_ (
    .A(_233_),
    .B(dbg_reg_din[0]),
    .Y(_245_)
  );
  \$_AND_  _601_ (
    .A(_245_),
    .B(_244_),
    .Y(_246_)
  );
  \$_OR_  _602_ (
    .A(_246_),
    .B(_235_),
    .Y(_247_)
  );
  \$_MUX_  _603_ (
    .A(_247_),
    .B(inst_sext[0]),
    .S(_228_),
    .Y(_248_)
  );
  \$_MUX_  _604_ (
    .A(_248_),
    .B(dbg_mem_dout[0]),
    .S(dbg_halt_st),
    .Y(op_dst[0])
  );
  \$_AND_  _605_ (
    .A(_131_),
    .B(_031_),
    .Y(_249_)
  );
  \$_OR_  _606_ (
    .A(_084_),
    .B(_055_),
    .Y(_250_)
  );
  \$_OR_  _607_ (
    .A(_250_),
    .B(_018_),
    .Y(_251_)
  );
  \$_OR_  _608_ (
    .A(_251_),
    .B(_047_),
    .Y(_252_)
  );
  \$_OR_  _609_ (
    .A(_252_),
    .B(_249_),
    .Y(_253_)
  );
  \$_MUX_  _610_ (
    .A(_253_),
    .B(dbg_reg_din[10]),
    .S(_244_),
    .Y(_254_)
  );
  \$_MUX_  _611_ (
    .A(_254_),
    .B(mdb_in[10]),
    .S(_234_),
    .Y(_255_)
  );
  \$_MUX_  _612_ (
    .A(_255_),
    .B(inst_sext[10]),
    .S(_228_),
    .Y(_256_)
  );
  \$_MUX_  _613_ (
    .A(_256_),
    .B(dbg_mem_dout[10]),
    .S(dbg_halt_st),
    .Y(op_dst[10])
  );
  \$_MUX_  _614_ (
    .A(_253_),
    .B(dbg_reg_din[11]),
    .S(_244_),
    .Y(_257_)
  );
  \$_MUX_  _615_ (
    .A(_257_),
    .B(mdb_in[11]),
    .S(_234_),
    .Y(_258_)
  );
  \$_MUX_  _616_ (
    .A(_258_),
    .B(inst_sext[11]),
    .S(_228_),
    .Y(_259_)
  );
  \$_MUX_  _617_ (
    .A(_259_),
    .B(dbg_mem_dout[11]),
    .S(dbg_halt_st),
    .Y(op_dst[11])
  );
  \$_MUX_  _618_ (
    .A(_253_),
    .B(dbg_reg_din[12]),
    .S(_244_),
    .Y(_260_)
  );
  \$_MUX_  _619_ (
    .A(_260_),
    .B(mdb_in[12]),
    .S(_234_),
    .Y(_261_)
  );
  \$_MUX_  _620_ (
    .A(_261_),
    .B(inst_sext[12]),
    .S(_228_),
    .Y(_262_)
  );
  \$_MUX_  _621_ (
    .A(_262_),
    .B(dbg_mem_dout[12]),
    .S(dbg_halt_st),
    .Y(op_dst[12])
  );
  \$_MUX_  _622_ (
    .A(_253_),
    .B(dbg_reg_din[13]),
    .S(_244_),
    .Y(_263_)
  );
  \$_MUX_  _623_ (
    .A(_263_),
    .B(mdb_in[13]),
    .S(_234_),
    .Y(_264_)
  );
  \$_MUX_  _624_ (
    .A(_264_),
    .B(inst_sext[13]),
    .S(_228_),
    .Y(_265_)
  );
  \$_MUX_  _625_ (
    .A(_265_),
    .B(dbg_mem_dout[13]),
    .S(dbg_halt_st),
    .Y(op_dst[13])
  );
  \$_MUX_  _626_ (
    .A(_253_),
    .B(dbg_reg_din[14]),
    .S(_244_),
    .Y(_266_)
  );
  \$_MUX_  _627_ (
    .A(_266_),
    .B(mdb_in[14]),
    .S(_234_),
    .Y(_267_)
  );
  \$_MUX_  _628_ (
    .A(_267_),
    .B(inst_sext[14]),
    .S(_228_),
    .Y(_268_)
  );
  \$_MUX_  _629_ (
    .A(_268_),
    .B(dbg_mem_dout[14]),
    .S(dbg_halt_st),
    .Y(op_dst[14])
  );
  \$_MUX_  _630_ (
    .A(_253_),
    .B(dbg_reg_din[15]),
    .S(_244_),
    .Y(_269_)
  );
  \$_MUX_  _631_ (
    .A(_269_),
    .B(mdb_in[15]),
    .S(_234_),
    .Y(_270_)
  );
  \$_MUX_  _632_ (
    .A(_270_),
    .B(inst_sext[15]),
    .S(_228_),
    .Y(_271_)
  );
  \$_MUX_  _633_ (
    .A(_271_),
    .B(dbg_mem_dout[15]),
    .S(dbg_halt_st),
    .Y(op_dst[15])
  );
  \$_MUX_  _634_ (
    .A(_253_),
    .B(dbg_reg_din[1]),
    .S(_244_),
    .Y(_272_)
  );
  \$_MUX_  _635_ (
    .A(_272_),
    .B(_109_),
    .S(_234_),
    .Y(_273_)
  );
  \$_MUX_  _636_ (
    .A(_273_),
    .B(inst_sext[1]),
    .S(_228_),
    .Y(_274_)
  );
  \$_MUX_  _637_ (
    .A(_274_),
    .B(dbg_mem_dout[1]),
    .S(dbg_halt_st),
    .Y(op_dst[1])
  );
  \$_MUX_  _638_ (
    .A(_253_),
    .B(dbg_reg_din[2]),
    .S(_244_),
    .Y(_275_)
  );
  \$_MUX_  _639_ (
    .A(_275_),
    .B(_111_),
    .S(_234_),
    .Y(_276_)
  );
  \$_MUX_  _640_ (
    .A(_276_),
    .B(inst_sext[2]),
    .S(_228_),
    .Y(_277_)
  );
  \$_MUX_  _641_ (
    .A(_277_),
    .B(dbg_mem_dout[2]),
    .S(dbg_halt_st),
    .Y(op_dst[2])
  );
  \$_MUX_  _642_ (
    .A(_253_),
    .B(dbg_reg_din[3]),
    .S(_244_),
    .Y(_278_)
  );
  \$_MUX_  _643_ (
    .A(_278_),
    .B(_113_),
    .S(_234_),
    .Y(_279_)
  );
  \$_MUX_  _644_ (
    .A(_279_),
    .B(inst_sext[3]),
    .S(_228_),
    .Y(_280_)
  );
  \$_MUX_  _645_ (
    .A(_280_),
    .B(dbg_mem_dout[3]),
    .S(dbg_halt_st),
    .Y(op_dst[3])
  );
  \$_MUX_  _646_ (
    .A(_253_),
    .B(dbg_reg_din[4]),
    .S(_244_),
    .Y(_281_)
  );
  \$_MUX_  _647_ (
    .A(_281_),
    .B(_115_),
    .S(_234_),
    .Y(_282_)
  );
  \$_MUX_  _648_ (
    .A(_282_),
    .B(inst_sext[4]),
    .S(_228_),
    .Y(_283_)
  );
  \$_MUX_  _649_ (
    .A(_283_),
    .B(dbg_mem_dout[4]),
    .S(dbg_halt_st),
    .Y(op_dst[4])
  );
  \$_MUX_  _650_ (
    .A(_253_),
    .B(dbg_reg_din[5]),
    .S(_244_),
    .Y(_284_)
  );
  \$_MUX_  _651_ (
    .A(_284_),
    .B(_117_),
    .S(_234_),
    .Y(_285_)
  );
  \$_MUX_  _652_ (
    .A(_285_),
    .B(inst_sext[5]),
    .S(_228_),
    .Y(_286_)
  );
  \$_MUX_  _653_ (
    .A(_286_),
    .B(dbg_mem_dout[5]),
    .S(dbg_halt_st),
    .Y(op_dst[5])
  );
  \$_MUX_  _654_ (
    .A(_253_),
    .B(dbg_reg_din[6]),
    .S(_244_),
    .Y(_287_)
  );
  \$_MUX_  _655_ (
    .A(_287_),
    .B(_119_),
    .S(_234_),
    .Y(_288_)
  );
  \$_MUX_  _656_ (
    .A(_288_),
    .B(inst_sext[6]),
    .S(_228_),
    .Y(_289_)
  );
  \$_MUX_  _657_ (
    .A(_289_),
    .B(dbg_mem_dout[6]),
    .S(dbg_halt_st),
    .Y(op_dst[6])
  );
  \$_MUX_  _658_ (
    .A(_253_),
    .B(dbg_reg_din[7]),
    .S(_244_),
    .Y(_290_)
  );
  \$_MUX_  _659_ (
    .A(_290_),
    .B(_121_),
    .S(_234_),
    .Y(_291_)
  );
  \$_MUX_  _660_ (
    .A(_291_),
    .B(inst_sext[7]),
    .S(_228_),
    .Y(_292_)
  );
  \$_MUX_  _661_ (
    .A(_292_),
    .B(dbg_mem_dout[7]),
    .S(dbg_halt_st),
    .Y(op_dst[7])
  );
  \$_MUX_  _662_ (
    .A(_253_),
    .B(dbg_reg_din[8]),
    .S(_244_),
    .Y(_293_)
  );
  \$_MUX_  _663_ (
    .A(_293_),
    .B(mdb_in[8]),
    .S(_234_),
    .Y(_294_)
  );
  \$_MUX_  _664_ (
    .A(_294_),
    .B(inst_sext[8]),
    .S(_228_),
    .Y(_295_)
  );
  \$_MUX_  _665_ (
    .A(_295_),
    .B(dbg_mem_dout[8]),
    .S(dbg_halt_st),
    .Y(op_dst[8])
  );
  \$_MUX_  _666_ (
    .A(_253_),
    .B(dbg_reg_din[9]),
    .S(_244_),
    .Y(_296_)
  );
  \$_MUX_  _667_ (
    .A(_296_),
    .B(mdb_in[9]),
    .S(_234_),
    .Y(_297_)
  );
  \$_MUX_  _668_ (
    .A(_297_),
    .B(inst_sext[9]),
    .S(_228_),
    .Y(_298_)
  );
  \$_MUX_  _669_ (
    .A(_298_),
    .B(dbg_mem_dout[9]),
    .S(dbg_halt_st),
    .Y(op_dst[9])
  );
  \$_MUX_  _670_ (
    .A(mdb_out_nxt[10]),
    .B(mdb_out[2]),
    .S(inst_bw),
    .Y(mdb_out[10])
  );
  \$_MUX_  _671_ (
    .A(mdb_out_nxt[11]),
    .B(mdb_out[3]),
    .S(inst_bw),
    .Y(mdb_out[11])
  );
  \$_MUX_  _672_ (
    .A(mdb_out_nxt[12]),
    .B(mdb_out[4]),
    .S(inst_bw),
    .Y(mdb_out[12])
  );
  \$_MUX_  _673_ (
    .A(mdb_out_nxt[13]),
    .B(mdb_out[5]),
    .S(inst_bw),
    .Y(mdb_out[13])
  );
  \$_MUX_  _674_ (
    .A(mdb_out_nxt[14]),
    .B(mdb_out[6]),
    .S(inst_bw),
    .Y(mdb_out[14])
  );
  \$_MUX_  _675_ (
    .A(mdb_out_nxt[15]),
    .B(mdb_out[7]),
    .S(inst_bw),
    .Y(mdb_out[15])
  );
  \$_MUX_  _676_ (
    .A(mdb_out_nxt[8]),
    .B(mdb_out[0]),
    .S(inst_bw),
    .Y(mdb_out[8])
  );
  \$_MUX_  _677_ (
    .A(mdb_out_nxt[9]),
    .B(mdb_out[1]),
    .S(inst_bw),
    .Y(mdb_out[9])
  );
  \$_DFF_PP0_  \mdb_out_reg[0]  /* _678_ */ (
    .C(mclk),
    .D(_004_[0]),
    .Q(mdb_out[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[10]  /* _679_ */ (
    .C(mclk),
    .D(_004_[10]),
    .Q(mdb_out_nxt[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[11]  /* _680_ */ (
    .C(mclk),
    .D(_004_[11]),
    .Q(mdb_out_nxt[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[12]  /* _681_ */ (
    .C(mclk),
    .D(_004_[12]),
    .Q(mdb_out_nxt[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[13]  /* _682_ */ (
    .C(mclk),
    .D(_004_[13]),
    .Q(mdb_out_nxt[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[14]  /* _683_ */ (
    .C(mclk),
    .D(_004_[14]),
    .Q(mdb_out_nxt[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[15]  /* _684_ */ (
    .C(mclk),
    .D(_004_[15]),
    .Q(mdb_out_nxt[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[1]  /* _685_ */ (
    .C(mclk),
    .D(_004_[1]),
    .Q(mdb_out[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[2]  /* _686_ */ (
    .C(mclk),
    .D(_004_[2]),
    .Q(mdb_out[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[3]  /* _687_ */ (
    .C(mclk),
    .D(_004_[3]),
    .Q(mdb_out[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[4]  /* _688_ */ (
    .C(mclk),
    .D(_004_[4]),
    .Q(mdb_out[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[5]  /* _689_ */ (
    .C(mclk),
    .D(_004_[5]),
    .Q(mdb_out[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[6]  /* _690_ */ (
    .C(mclk),
    .D(_004_[6]),
    .Q(mdb_out[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_reg[7]  /* _691_ */ (
    .C(mclk),
    .D(_004_[7]),
    .Q(mdb_out[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[8]  /* _692_ */ (
    .C(mclk),
    .D(_004_[8]),
    .Q(mdb_out_nxt[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_out_nxt_reg[9]  /* _693_ */ (
    .C(mclk),
    .D(_004_[9]),
    .Q(mdb_out_nxt[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  mab_lsb_reg /* _694_ */ (
    .C(mclk),
    .D(_000_),
    .Q(mab_lsb),
    .R(puc_rst)
  );
  \$_DFF_PP0_  mdb_in_buf_en_reg /* _695_ */ (
    .C(mclk),
    .D(_002_),
    .Q(mdb_in_buf_en),
    .R(puc_rst)
  );
  \$_DFF_PP0_  mdb_in_buf_valid_reg /* _696_ */ (
    .C(mclk),
    .D(_003_),
    .Q(mdb_in_buf_valid),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[0]  /* _697_ */ (
    .C(mclk),
    .D(_001_[0]),
    .Q(mdb_in_buf[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[10]  /* _698_ */ (
    .C(mclk),
    .D(_001_[10]),
    .Q(mdb_in_buf[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[11]  /* _699_ */ (
    .C(mclk),
    .D(_001_[11]),
    .Q(mdb_in_buf[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[12]  /* _700_ */ (
    .C(mclk),
    .D(_001_[12]),
    .Q(mdb_in_buf[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[13]  /* _701_ */ (
    .C(mclk),
    .D(_001_[13]),
    .Q(mdb_in_buf[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[14]  /* _702_ */ (
    .C(mclk),
    .D(_001_[14]),
    .Q(mdb_in_buf[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[15]  /* _703_ */ (
    .C(mclk),
    .D(_001_[15]),
    .Q(mdb_in_buf[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[1]  /* _704_ */ (
    .C(mclk),
    .D(_001_[1]),
    .Q(mdb_in_buf[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[2]  /* _705_ */ (
    .C(mclk),
    .D(_001_[2]),
    .Q(mdb_in_buf[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[3]  /* _706_ */ (
    .C(mclk),
    .D(_001_[3]),
    .Q(mdb_in_buf[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[4]  /* _707_ */ (
    .C(mclk),
    .D(_001_[4]),
    .Q(mdb_in_buf[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[5]  /* _708_ */ (
    .C(mclk),
    .D(_001_[5]),
    .Q(mdb_in_buf[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[6]  /* _709_ */ (
    .C(mclk),
    .D(_001_[6]),
    .Q(mdb_in_buf[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[7]  /* _710_ */ (
    .C(mclk),
    .D(_001_[7]),
    .Q(mdb_in_buf[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[8]  /* _711_ */ (
    .C(mclk),
    .D(_001_[8]),
    .Q(mdb_in_buf[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \mdb_in_buf_reg[9]  /* _712_ */ (
    .C(mclk),
    .D(_001_[9]),
    .Q(mdb_in_buf[9]),
    .R(puc_rst)
  );
  omsp_alu alu_0 (
    .alu_out(alu_out),
    .alu_out_add(alu_out_add),
    .alu_stat(alu_stat),
    .alu_stat_wr(alu_stat_wr),
    .dbg_halt_st(dbg_halt_st),
    .exec_cycle(exec_cycle),
    .inst_alu(inst_alu),
    .inst_bw(inst_bw),
    .inst_jmp(inst_jmp),
    .inst_so(inst_so),
    .op_dst(op_dst),
    .op_src(op_src),
    .status(status)
  );
  omsp_register_file register_file_0 (
    .alu_stat(alu_stat),
    .alu_stat_wr(alu_stat_wr),
    .cpuoff(cpuoff),
    .gie(gie),
    .inst_bw(inst_bw),
    .inst_dest(inst_dest),
    .inst_src(inst_src),
    .mclk(mclk),
    .oscoff(oscoff),
    .pc(pc),
    .pc_sw(pc_sw),
    .pc_sw_wr(pc_sw_wr),
    .puc_rst(puc_rst),
    .reg_dest(dbg_reg_din),
    .reg_dest_val(alu_out),
    .reg_dest_wr(reg_dest_wr),
    .reg_incr(reg_incr),
    .reg_pc_call(reg_pc_call),
    .reg_sp_val(alu_out_add),
    .reg_sp_wr(reg_sp_wr),
    .reg_sr_clr(reg_sr_clr),
    .reg_sr_wr(reg_sr_wr),
    .reg_src(reg_src),
    .scan_enable(scan_enable),
    .scg0(scg0),
    .scg1(scg1),
    .status(status)
  );
  assign mab = alu_out_add;
  assign mclk_mdb_in_buf = mclk;
  assign mclk_mdb_out_nxt = mclk;
  assign mdb_in_bw[15:8] = mdb_in[15:8];
  assign mdb_out_nxt[7:0] = mdb_out[7:0];
  assign reg_dest = dbg_reg_din;
endmodule

module omsp_frontend(dbg_halt_st, decode_noirq, e_state, exec_done, inst_ad, inst_as, inst_alu, inst_bw, inst_dest, inst_dext, inst_irq_rst, inst_jmp, inst_mov, inst_sext, inst_so, inst_src, inst_type, irq_acc, mab, mb_en, mclk_enable, mclk_wkup, nmi_acc, pc, pc_nxt, cpu_en_s, cpuoff, dbg_halt_cmd, dbg_reg_sel, fe_pmem_wait, gie, irq, mclk, mdb_in, nmi_pnd, nmi_wkup, pc_sw, pc_sw_wr, puc_rst, scan_enable, wdt_irq, wdt_wkup, wkup);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire [7:0] _0005_;
  wire [11:0] _0006_;
  wire [7:0] _0007_;
  wire _0008_;
  wire [3:0] _0009_;
  wire [15:0] _0010_;
  wire _0011_;
  wire [2:0] _0012_;
  wire _0013_;
  wire [15:0] _0014_;
  wire [7:0] _0015_;
  wire [3:0] _0016_;
  wire [1:0] _0017_;
  wire [2:0] _0018_;
  wire [3:0] _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire [15:0] _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  input cpu_en_s;
  input cpuoff;
  input dbg_halt_cmd;
  output dbg_halt_st;
  input [3:0] dbg_reg_sel;
  output decode_noirq;
  wire [3:0] dest_reg;
  output [3:0] e_state;
  wire [3:0] e_state_nxt;
  wire exec_dext_rdy;
  output exec_done;
  wire exec_dst_wr;
  wire exec_jmp;
  wire exec_src_wr;
  wire [15:0] ext_nxt;
  input fe_pmem_wait;
  input gie;
  wire [4:0] i_state;
  output [7:0] inst_ad;
  output [11:0] inst_alu;
  output [7:0] inst_as;
  output inst_bw;
  output [15:0] inst_dest;
  wire [3:0] inst_dest_bin;
  output [15:0] inst_dext;
  output inst_irq_rst;
  output [7:0] inst_jmp;
  wire [2:0] inst_jmp_bin;
  output inst_mov;
  output [15:0] inst_sext;
  output [7:0] inst_so;
  output [15:0] inst_src;
  wire [3:0] inst_src_bin;
  wire [1:0] inst_sz;
  output [2:0] inst_type;
  wire [15:0] ir;
  input [13:0] irq;
  output [13:0] irq_acc;
  wire [15:0] irq_acc_all;
  wire [15:0] irq_addr;
  wire [3:0] irq_num;
  output [15:0] mab;
  output mb_en;
  input mclk;
  wire mclk_decode;
  output mclk_enable;
  wire mclk_inst_dext;
  wire mclk_inst_sext;
  wire mclk_irq_num;
  wire mclk_pc;
  output mclk_wkup;
  input [15:0] mdb_in;
  output nmi_acc;
  input nmi_pnd;
  input nmi_wkup;
  output [15:0] pc;
  wire [15:0] pc_incr;
  output [15:0] pc_nxt;
  input [15:0] pc_sw;
  input pc_sw_wr;
  wire pmem_busy;
  input puc_rst;
  input scan_enable;
  input wdt_irq;
  input wdt_wkup;
  input wkup;
  \$_INV_  _1147_ (
    .A(e_state[1]),
    .Y(_0566_)
  );
  \$_INV_  _1148_ (
    .A(e_state[0]),
    .Y(_0567_)
  );
  \$_AND_  _1149_ (
    .A(_0567_),
    .B(_0566_),
    .Y(_0568_)
  );
  \$_AND_  _1150_ (
    .A(_0568_),
    .B(e_state[2]),
    .Y(_0569_)
  );
  \$_AND_  _1151_ (
    .A(_0569_),
    .B(e_state[3]),
    .Y(_0570_)
  );
  \$_INV_  _1152_ (
    .A(e_state[2]),
    .Y(_0571_)
  );
  \$_AND_  _1153_ (
    .A(_0567_),
    .B(e_state[1]),
    .Y(_0572_)
  );
  \$_AND_  _1154_ (
    .A(_0572_),
    .B(_0571_),
    .Y(_0573_)
  );
  \$_AND_  _1155_ (
    .A(_0573_),
    .B(e_state[3]),
    .Y(_0574_)
  );
  \$_AND_  _1156_ (
    .A(e_state[0]),
    .B(e_state[1]),
    .Y(_0575_)
  );
  \$_INV_  _1157_ (
    .A(e_state[3]),
    .Y(_0576_)
  );
  \$_AND_  _1158_ (
    .A(_0576_),
    .B(e_state[2]),
    .Y(_0577_)
  );
  \$_AND_  _1159_ (
    .A(_0577_),
    .B(_0575_),
    .Y(_0578_)
  );
  \$_AND_  _1160_ (
    .A(_0575_),
    .B(_0571_),
    .Y(_0579_)
  );
  \$_AND_  _1161_ (
    .A(_0579_),
    .B(e_state[3]),
    .Y(_0580_)
  );
  \$_MUX_  _1162_ (
    .A(_0580_),
    .B(_0578_),
    .S(exec_src_wr),
    .Y(_0581_)
  );
  \$_MUX_  _1163_ (
    .A(_0581_),
    .B(_0574_),
    .S(exec_dst_wr),
    .Y(_0582_)
  );
  \$_MUX_  _1164_ (
    .A(_0582_),
    .B(_0570_),
    .S(exec_jmp),
    .Y(exec_done)
  );
  \$_INV_  _1165_ (
    .A(exec_done),
    .Y(_0583_)
  );
  \$_AND_  _1166_ (
    .A(e_state[0]),
    .B(_0566_),
    .Y(_0584_)
  );
  \$_AND_  _1167_ (
    .A(_0584_),
    .B(e_state[2]),
    .Y(_0585_)
  );
  \$_AND_  _1168_ (
    .A(_0585_),
    .B(e_state[3]),
    .Y(_0586_)
  );
  \$_INV_  _1169_ (
    .A(_0586_),
    .Y(_0587_)
  );
  \$_AND_  _1170_ (
    .A(_0587_),
    .B(_0583_),
    .Y(_0588_)
  );
  \$_INV_  _1171_ (
    .A(_0588_),
    .Y(_0589_)
  );
  \$_AND_  _1172_ (
    .A(_0589_),
    .B(i_state[1]),
    .Y(decode_noirq)
  );
  \$_INV_  _1173_ (
    .A(mdb_in[11]),
    .Y(_0590_)
  );
  \$_INV_  _1174_ (
    .A(mdb_in[3]),
    .Y(_0591_)
  );
  \$_OR_  _1175_ (
    .A(exec_done),
    .B(i_state[3]),
    .Y(_0592_)
  );
  \$_OR_  _1176_ (
    .A(irq[1]),
    .B(irq[0]),
    .Y(_0593_)
  );
  \$_OR_  _1177_ (
    .A(_0593_),
    .B(irq[2]),
    .Y(_0594_)
  );
  \$_OR_  _1178_ (
    .A(irq[4]),
    .B(irq[3]),
    .Y(_0595_)
  );
  \$_OR_  _1179_ (
    .A(_0595_),
    .B(_0594_),
    .Y(_0596_)
  );
  \$_OR_  _1180_ (
    .A(irq[6]),
    .B(irq[5]),
    .Y(_0597_)
  );
  \$_OR_  _1181_ (
    .A(irq[8]),
    .B(irq[7]),
    .Y(_0598_)
  );
  \$_OR_  _1182_ (
    .A(_0598_),
    .B(_0597_),
    .Y(_0599_)
  );
  \$_OR_  _1183_ (
    .A(_0599_),
    .B(_0596_),
    .Y(_0600_)
  );
  \$_OR_  _1184_ (
    .A(irq[10]),
    .B(wdt_irq),
    .Y(_0601_)
  );
  \$_OR_  _1185_ (
    .A(irq[12]),
    .B(irq[11]),
    .Y(_0602_)
  );
  \$_OR_  _1186_ (
    .A(irq[9]),
    .B(irq[13]),
    .Y(_0603_)
  );
  \$_OR_  _1187_ (
    .A(_0603_),
    .B(_0602_),
    .Y(_0604_)
  );
  \$_OR_  _1188_ (
    .A(_0604_),
    .B(_0601_),
    .Y(_0605_)
  );
  \$_OR_  _1189_ (
    .A(_0605_),
    .B(_0600_),
    .Y(_0606_)
  );
  \$_AND_  _1190_ (
    .A(_0606_),
    .B(gie),
    .Y(_0607_)
  );
  \$_OR_  _1191_ (
    .A(_0607_),
    .B(nmi_pnd),
    .Y(_0608_)
  );
  \$_INV_  _1192_ (
    .A(dbg_halt_st),
    .Y(_0609_)
  );
  \$_INV_  _1193_ (
    .A(dbg_halt_cmd),
    .Y(_0610_)
  );
  \$_AND_  _1194_ (
    .A(_0610_),
    .B(cpu_en_s),
    .Y(_0611_)
  );
  \$_AND_  _1195_ (
    .A(_0611_),
    .B(_0609_),
    .Y(_0612_)
  );
  \$_AND_  _1196_ (
    .A(_0612_),
    .B(_0608_),
    .Y(_0613_)
  );
  \$_AND_  _1197_ (
    .A(_0613_),
    .B(_0592_),
    .Y(_0614_)
  );
  \$_INV_  _1198_ (
    .A(mdb_in[15]),
    .Y(_0615_)
  );
  \$_INV_  _1199_ (
    .A(mdb_in[13]),
    .Y(_0616_)
  );
  \$_INV_  _1200_ (
    .A(mdb_in[14]),
    .Y(_0617_)
  );
  \$_AND_  _1201_ (
    .A(_0617_),
    .B(_0616_),
    .Y(_0618_)
  );
  \$_AND_  _1202_ (
    .A(_0618_),
    .B(_0615_),
    .Y(_0619_)
  );
  \$_INV_  _1203_ (
    .A(_0619_),
    .Y(_0620_)
  );
  \$_OR_  _1204_ (
    .A(_0620_),
    .B(_0614_),
    .Y(_0621_)
  );
  \$_MUX_  _1205_ (
    .A(_0591_),
    .B(_0590_),
    .S(_0621_),
    .Y(_0622_)
  );
  \$_INV_  _1206_ (
    .A(mdb_in[10]),
    .Y(_0623_)
  );
  \$_INV_  _1207_ (
    .A(mdb_in[2]),
    .Y(_0624_)
  );
  \$_MUX_  _1208_ (
    .A(_0624_),
    .B(_0623_),
    .S(_0621_),
    .Y(_0625_)
  );
  \$_AND_  _1209_ (
    .A(_0625_),
    .B(_0622_),
    .Y(_0626_)
  );
  \$_MUX_  _1210_ (
    .A(mdb_in[1]),
    .B(mdb_in[9]),
    .S(_0621_),
    .Y(_0627_)
  );
  \$_INV_  _1211_ (
    .A(mdb_in[8]),
    .Y(_0628_)
  );
  \$_INV_  _1212_ (
    .A(mdb_in[0]),
    .Y(_0629_)
  );
  \$_MUX_  _1213_ (
    .A(_0629_),
    .B(_0628_),
    .S(_0621_),
    .Y(_0630_)
  );
  \$_AND_  _1214_ (
    .A(_0630_),
    .B(_0627_),
    .Y(_0631_)
  );
  \$_AND_  _1215_ (
    .A(_0631_),
    .B(_0626_),
    .Y(_0632_)
  );
  \$_MUX_  _1216_ (
    .A(mdb_in[3]),
    .B(mdb_in[11]),
    .S(_0621_),
    .Y(_0633_)
  );
  \$_MUX_  _1217_ (
    .A(mdb_in[2]),
    .B(mdb_in[10]),
    .S(_0621_),
    .Y(_0634_)
  );
  \$_OR_  _1218_ (
    .A(_0634_),
    .B(_0633_),
    .Y(_0635_)
  );
  \$_INV_  _1219_ (
    .A(mdb_in[1]),
    .Y(_0636_)
  );
  \$_INV_  _1220_ (
    .A(mdb_in[9]),
    .Y(_0637_)
  );
  \$_MUX_  _1221_ (
    .A(_0636_),
    .B(_0637_),
    .S(_0621_),
    .Y(_0638_)
  );
  \$_OR_  _1222_ (
    .A(_0630_),
    .B(_0638_),
    .Y(_0639_)
  );
  \$_OR_  _1223_ (
    .A(_0639_),
    .B(_0635_),
    .Y(_0640_)
  );
  \$_AND_  _1224_ (
    .A(_0617_),
    .B(mdb_in[13]),
    .Y(_0641_)
  );
  \$_AND_  _1225_ (
    .A(_0641_),
    .B(_0615_),
    .Y(_0642_)
  );
  \$_INV_  _1226_ (
    .A(_0642_),
    .Y(_0643_)
  );
  \$_OR_  _1227_ (
    .A(_0643_),
    .B(_0614_),
    .Y(_0644_)
  );
  \$_INV_  _1228_ (
    .A(mdb_in[5]),
    .Y(_0645_)
  );
  \$_AND_  _1229_ (
    .A(_0645_),
    .B(mdb_in[4]),
    .Y(_0646_)
  );
  \$_AND_  _1230_ (
    .A(_0646_),
    .B(_0644_),
    .Y(_0647_)
  );
  \$_AND_  _1231_ (
    .A(_0647_),
    .B(_0640_),
    .Y(_0648_)
  );
  \$_AND_  _1232_ (
    .A(_0648_),
    .B(_0632_),
    .Y(_0649_)
  );
  \$_MUX_  _1233_ (
    .A(mdb_in[0]),
    .B(mdb_in[8]),
    .S(_0621_),
    .Y(_0650_)
  );
  \$_OR_  _1234_ (
    .A(_0650_),
    .B(_0638_),
    .Y(_0651_)
  );
  \$_OR_  _1235_ (
    .A(_0651_),
    .B(_0635_),
    .Y(_0652_)
  );
  \$_AND_  _1236_ (
    .A(_0630_),
    .B(_0638_),
    .Y(_0653_)
  );
  \$_AND_  _1237_ (
    .A(_0653_),
    .B(_0626_),
    .Y(_0654_)
  );
  \$_AND_  _1238_ (
    .A(mdb_in[5]),
    .B(mdb_in[4]),
    .Y(_0655_)
  );
  \$_AND_  _1239_ (
    .A(_0655_),
    .B(_0644_),
    .Y(_0656_)
  );
  \$_AND_  _1240_ (
    .A(_0656_),
    .B(_0640_),
    .Y(_0657_)
  );
  \$_AND_  _1241_ (
    .A(_0657_),
    .B(_0654_),
    .Y(_0658_)
  );
  \$_OR_  _1242_ (
    .A(_0658_),
    .B(_0648_),
    .Y(_0659_)
  );
  \$_INV_  _1243_ (
    .A(_0621_),
    .Y(_0660_)
  );
  \$_INV_  _1244_ (
    .A(mdb_in[7]),
    .Y(_0661_)
  );
  \$_AND_  _1245_ (
    .A(_0615_),
    .B(_0617_),
    .Y(_0662_)
  );
  \$_OR_  _1246_ (
    .A(_0662_),
    .B(_0614_),
    .Y(_0663_)
  );
  \$_AND_  _1247_ (
    .A(_0624_),
    .B(mdb_in[1]),
    .Y(_0664_)
  );
  \$_AND_  _1248_ (
    .A(_0629_),
    .B(_0591_),
    .Y(_0665_)
  );
  \$_AND_  _1249_ (
    .A(_0665_),
    .B(_0664_),
    .Y(_0666_)
  );
  \$_AND_  _1250_ (
    .A(_0624_),
    .B(_0636_),
    .Y(_0667_)
  );
  \$_AND_  _1251_ (
    .A(_0667_),
    .B(_0665_),
    .Y(_0668_)
  );
  \$_OR_  _1252_ (
    .A(_0663_),
    .B(_0661_),
    .Y(_0669_)
  );
  \$_INV_  _1253_ (
    .A(_0669_),
    .Y(_0670_)
  );
  \$_OR_  _1254_ (
    .A(_0670_),
    .B(_0659_),
    .Y(_0671_)
  );
  \$_INV_  _1255_ (
    .A(_0614_),
    .Y(_0672_)
  );
  \$_INV_  _1256_ (
    .A(cpuoff),
    .Y(_0673_)
  );
  \$_AND_  _1257_ (
    .A(_0611_),
    .B(_0673_),
    .Y(_0674_)
  );
  \$_INV_  _1258_ (
    .A(_0674_),
    .Y(_0675_)
  );
  \$_AND_  _1259_ (
    .A(_0675_),
    .B(exec_done),
    .Y(_0676_)
  );
  \$_INV_  _1260_ (
    .A(_0676_),
    .Y(_0677_)
  );
  \$_INV_  _1261_ (
    .A(pc_sw_wr),
    .Y(_0678_)
  );
  \$_INV_  _1262_ (
    .A(_0611_),
    .Y(_0679_)
  );
  \$_AND_  _1263_ (
    .A(_0679_),
    .B(_0586_),
    .Y(_0680_)
  );
  \$_INV_  _1264_ (
    .A(_0680_),
    .Y(_0681_)
  );
  \$_AND_  _1265_ (
    .A(_0681_),
    .B(_0678_),
    .Y(_0682_)
  );
  \$_AND_  _1266_ (
    .A(_0682_),
    .B(_0677_),
    .Y(_0683_)
  );
  \$_AND_  _1267_ (
    .A(_0683_),
    .B(_0672_),
    .Y(_0684_)
  );
  \$_AND_  _1268_ (
    .A(_0684_),
    .B(_0589_),
    .Y(_0685_)
  );
  \$_AND_  _1269_ (
    .A(_0685_),
    .B(i_state[1]),
    .Y(_0686_)
  );
  \$_INV_  _1270_ (
    .A(_0686_),
    .Y(_0687_)
  );
  \$_OR_  _1271_ (
    .A(_0687_),
    .B(_0671_),
    .Y(_0688_)
  );
  \$_AND_  _1272_ (
    .A(_0588_),
    .B(i_state[1]),
    .Y(_0689_)
  );
  \$_AND_  _1273_ (
    .A(_0689_),
    .B(_0684_),
    .Y(_0690_)
  );
  \$_AND_  _1274_ (
    .A(_0674_),
    .B(i_state[3]),
    .Y(_0691_)
  );
  \$_AND_  _1275_ (
    .A(_0691_),
    .B(_0672_),
    .Y(_0692_)
  );
  \$_AND_  _1276_ (
    .A(pc_sw_wr),
    .B(i_state[1]),
    .Y(_0693_)
  );
  \$_AND_  _1277_ (
    .A(_0693_),
    .B(_0681_),
    .Y(_0694_)
  );
  \$_AND_  _1278_ (
    .A(_0694_),
    .B(_0677_),
    .Y(_0695_)
  );
  \$_AND_  _1279_ (
    .A(_0695_),
    .B(_0672_),
    .Y(_0696_)
  );
  \$_AND_  _1280_ (
    .A(pc_sw_wr),
    .B(i_state[4]),
    .Y(_0697_)
  );
  \$_INV_  _1281_ (
    .A(inst_sz[1]),
    .Y(_0698_)
  );
  \$_AND_  _1282_ (
    .A(_0698_),
    .B(inst_sz[0]),
    .Y(_0699_)
  );
  \$_AND_  _1283_ (
    .A(_0678_),
    .B(i_state[4]),
    .Y(_0700_)
  );
  \$_AND_  _1284_ (
    .A(_0700_),
    .B(_0699_),
    .Y(_0701_)
  );
  \$_OR_  _1285_ (
    .A(_0701_),
    .B(_0697_),
    .Y(_0702_)
  );
  \$_OR_  _1286_ (
    .A(_0702_),
    .B(_0696_),
    .Y(_0703_)
  );
  \$_OR_  _1287_ (
    .A(_0703_),
    .B(_0692_),
    .Y(_0704_)
  );
  \$_OR_  _1288_ (
    .A(_0704_),
    .B(_0690_),
    .Y(_0705_)
  );
  \$_INV_  _1289_ (
    .A(_0705_),
    .Y(_0706_)
  );
  \$_AND_  _1290_ (
    .A(_0706_),
    .B(_0688_),
    .Y(_0707_)
  );
  \$_AND_  _1291_ (
    .A(_0650_),
    .B(_0627_),
    .Y(_0708_)
  );
  \$_AND_  _1292_ (
    .A(_0708_),
    .B(_0626_),
    .Y(_0709_)
  );
  \$_INV_  _1293_ (
    .A(_0647_),
    .Y(_0710_)
  );
  \$_OR_  _1294_ (
    .A(_0710_),
    .B(_0709_),
    .Y(_0711_)
  );
  \$_OR_  _1295_ (
    .A(_0650_),
    .B(_0627_),
    .Y(_0712_)
  );
  \$_OR_  _1296_ (
    .A(_0712_),
    .B(_0635_),
    .Y(_0713_)
  );
  \$_INV_  _1297_ (
    .A(_0656_),
    .Y(_0714_)
  );
  \$_OR_  _1298_ (
    .A(_0714_),
    .B(_0709_),
    .Y(_0715_)
  );
  \$_OR_  _1299_ (
    .A(_0715_),
    .B(_0713_),
    .Y(_0716_)
  );
  \$_AND_  _1300_ (
    .A(_0716_),
    .B(_0711_),
    .Y(_0717_)
  );
  \$_AND_  _1301_ (
    .A(_0669_),
    .B(_0717_),
    .Y(_0718_)
  );
  \$_OR_  _1302_ (
    .A(_0687_),
    .B(_0718_),
    .Y(_0719_)
  );
  \$_OR_  _1303_ (
    .A(i_state[2]),
    .B(i_state[0]),
    .Y(_0720_)
  );
  \$_INV_  _1304_ (
    .A(_0720_),
    .Y(_0721_)
  );
  \$_AND_  _1305_ (
    .A(_0721_),
    .B(_0719_),
    .Y(_0722_)
  );
  \$_AND_  _1306_ (
    .A(_0722_),
    .B(_0707_),
    .Y(_0723_)
  );
  \$_INV_  _1307_ (
    .A(i_state[1]),
    .Y(_0724_)
  );
  \$_INV_  _1308_ (
    .A(i_state[4]),
    .Y(_0725_)
  );
  \$_AND_  _1309_ (
    .A(_0725_),
    .B(_0724_),
    .Y(_0726_)
  );
  \$_INV_  _1310_ (
    .A(i_state[3]),
    .Y(_0727_)
  );
  \$_AND_  _1311_ (
    .A(_0721_),
    .B(_0727_),
    .Y(_0728_)
  );
  \$_AND_  _1312_ (
    .A(_0728_),
    .B(_0726_),
    .Y(_1142_[15])
  );
  \$_INV_  _1313_ (
    .A(_1142_[15]),
    .Y(_0729_)
  );
  \$_AND_  _1314_ (
    .A(_0675_),
    .B(i_state[3]),
    .Y(_0730_)
  );
  \$_AND_  _1315_ (
    .A(_0730_),
    .B(_0672_),
    .Y(_0731_)
  );
  \$_INV_  _1316_ (
    .A(_0731_),
    .Y(_0732_)
  );
  \$_AND_  _1317_ (
    .A(_0676_),
    .B(i_state[1]),
    .Y(_0733_)
  );
  \$_AND_  _1318_ (
    .A(_0733_),
    .B(_0672_),
    .Y(_0734_)
  );
  \$_INV_  _1319_ (
    .A(_0734_),
    .Y(_0735_)
  );
  \$_AND_  _1320_ (
    .A(_0680_),
    .B(i_state[1]),
    .Y(_0736_)
  );
  \$_INV_  _1321_ (
    .A(_0736_),
    .Y(_0737_)
  );
  \$_AND_  _1322_ (
    .A(_0737_),
    .B(_0735_),
    .Y(_0738_)
  );
  \$_AND_  _1323_ (
    .A(_0738_),
    .B(_0732_),
    .Y(_0739_)
  );
  \$_AND_  _1324_ (
    .A(_0739_),
    .B(_0729_),
    .Y(_0740_)
  );
  \$_AND_  _1325_ (
    .A(_0740_),
    .B(_0719_),
    .Y(_0741_)
  );
  \$_INV_  _1326_ (
    .A(_0741_),
    .Y(_0742_)
  );
  \$_INV_  _1327_ (
    .A(_0699_),
    .Y(_0743_)
  );
  \$_AND_  _1328_ (
    .A(_0700_),
    .B(_0743_),
    .Y(_1143_)
  );
  \$_OR_  _1329_ (
    .A(_1143_),
    .B(_0734_),
    .Y(_0744_)
  );
  \$_OR_  _1330_ (
    .A(_0744_),
    .B(_0736_),
    .Y(_0745_)
  );
  \$_OR_  _1331_ (
    .A(_0745_),
    .B(_0731_),
    .Y(_0746_)
  );
  \$_AND_  _1332_ (
    .A(_0746_),
    .B(_0679_),
    .Y(_0747_)
  );
  \$_AND_  _1333_ (
    .A(_0747_),
    .B(_0742_),
    .Y(_0748_)
  );
  \$_AND_  _1334_ (
    .A(_0748_),
    .B(_0723_),
    .Y(_0000_)
  );
  \$_INV_  _1335_ (
    .A(irq_addr[4]),
    .Y(_0749_)
  );
  \$_INV_  _1336_ (
    .A(irq_addr[3]),
    .Y(_0750_)
  );
  \$_INV_  _1337_ (
    .A(irq_addr[1]),
    .Y(_0751_)
  );
  \$_INV_  _1338_ (
    .A(irq_addr[2]),
    .Y(_0752_)
  );
  \$_AND_  _1339_ (
    .A(_0752_),
    .B(_0751_),
    .Y(_0753_)
  );
  \$_AND_  _1340_ (
    .A(_0753_),
    .B(_0750_),
    .Y(_0754_)
  );
  \$_AND_  _1341_ (
    .A(_0754_),
    .B(_0749_),
    .Y(_0755_)
  );
  \$_AND_  _1342_ (
    .A(_0755_),
    .B(_1142_[15]),
    .Y(irq_acc[0])
  );
  \$_AND_  _1343_ (
    .A(irq_addr[2]),
    .B(_0751_),
    .Y(_0756_)
  );
  \$_AND_  _1344_ (
    .A(_0756_),
    .B(_0750_),
    .Y(_0757_)
  );
  \$_AND_  _1345_ (
    .A(_0757_),
    .B(irq_addr[4]),
    .Y(_0758_)
  );
  \$_AND_  _1346_ (
    .A(_0758_),
    .B(_1142_[15]),
    .Y(irq_acc[10])
  );
  \$_AND_  _1347_ (
    .A(irq_addr[2]),
    .B(irq_addr[1]),
    .Y(_0759_)
  );
  \$_AND_  _1348_ (
    .A(_0759_),
    .B(_0750_),
    .Y(_0760_)
  );
  \$_AND_  _1349_ (
    .A(_0760_),
    .B(irq_addr[4]),
    .Y(_0761_)
  );
  \$_AND_  _1350_ (
    .A(_0761_),
    .B(_1142_[15]),
    .Y(irq_acc[11])
  );
  \$_AND_  _1351_ (
    .A(_0753_),
    .B(irq_addr[3]),
    .Y(_0762_)
  );
  \$_AND_  _1352_ (
    .A(_0762_),
    .B(irq_addr[4]),
    .Y(_0763_)
  );
  \$_AND_  _1353_ (
    .A(_0763_),
    .B(_1142_[15]),
    .Y(irq_acc[12])
  );
  \$_AND_  _1354_ (
    .A(_0752_),
    .B(irq_addr[1]),
    .Y(_0764_)
  );
  \$_AND_  _1355_ (
    .A(_0764_),
    .B(irq_addr[3]),
    .Y(_0765_)
  );
  \$_AND_  _1356_ (
    .A(_0765_),
    .B(irq_addr[4]),
    .Y(_0766_)
  );
  \$_AND_  _1357_ (
    .A(_0766_),
    .B(_1142_[15]),
    .Y(irq_acc[13])
  );
  \$_AND_  _1358_ (
    .A(_0756_),
    .B(irq_addr[3]),
    .Y(_0767_)
  );
  \$_AND_  _1359_ (
    .A(_0767_),
    .B(irq_addr[4]),
    .Y(_0768_)
  );
  \$_AND_  _1360_ (
    .A(_0768_),
    .B(_1142_[15]),
    .Y(irq_acc_all[14])
  );
  \$_AND_  _1361_ (
    .A(_0764_),
    .B(_0750_),
    .Y(_0769_)
  );
  \$_AND_  _1362_ (
    .A(_0769_),
    .B(_0749_),
    .Y(_0770_)
  );
  \$_AND_  _1363_ (
    .A(_0770_),
    .B(_1142_[15]),
    .Y(irq_acc[1])
  );
  \$_AND_  _1364_ (
    .A(_0757_),
    .B(_0749_),
    .Y(_0771_)
  );
  \$_AND_  _1365_ (
    .A(_0771_),
    .B(_1142_[15]),
    .Y(irq_acc[2])
  );
  \$_AND_  _1366_ (
    .A(_0760_),
    .B(_0749_),
    .Y(_0772_)
  );
  \$_AND_  _1367_ (
    .A(_0772_),
    .B(_1142_[15]),
    .Y(irq_acc[3])
  );
  \$_AND_  _1368_ (
    .A(_0762_),
    .B(_0749_),
    .Y(_0773_)
  );
  \$_AND_  _1369_ (
    .A(_0773_),
    .B(_1142_[15]),
    .Y(irq_acc[4])
  );
  \$_AND_  _1370_ (
    .A(_0765_),
    .B(_0749_),
    .Y(_0774_)
  );
  \$_AND_  _1371_ (
    .A(_0774_),
    .B(_1142_[15]),
    .Y(irq_acc[5])
  );
  \$_AND_  _1372_ (
    .A(_0767_),
    .B(_0749_),
    .Y(_0775_)
  );
  \$_AND_  _1373_ (
    .A(_0775_),
    .B(_1142_[15]),
    .Y(irq_acc[6])
  );
  \$_AND_  _1374_ (
    .A(_0749_),
    .B(irq_addr[3]),
    .Y(_0776_)
  );
  \$_AND_  _1375_ (
    .A(_0776_),
    .B(_0759_),
    .Y(_0777_)
  );
  \$_AND_  _1376_ (
    .A(_0777_),
    .B(_1142_[15]),
    .Y(irq_acc[7])
  );
  \$_AND_  _1377_ (
    .A(_0754_),
    .B(irq_addr[4]),
    .Y(_0778_)
  );
  \$_AND_  _1378_ (
    .A(_0778_),
    .B(_1142_[15]),
    .Y(irq_acc[8])
  );
  \$_AND_  _1379_ (
    .A(_0769_),
    .B(irq_addr[4]),
    .Y(_0779_)
  );
  \$_AND_  _1380_ (
    .A(_0779_),
    .B(_1142_[15]),
    .Y(irq_acc[9])
  );
  \$_INV_  _1381_ (
    .A(inst_jmp_bin[2]),
    .Y(_0780_)
  );
  \$_INV_  _1382_ (
    .A(inst_jmp_bin[0]),
    .Y(_0781_)
  );
  \$_INV_  _1383_ (
    .A(inst_jmp_bin[1]),
    .Y(_0782_)
  );
  \$_AND_  _1384_ (
    .A(_0782_),
    .B(_0781_),
    .Y(_0783_)
  );
  \$_AND_  _1385_ (
    .A(_0783_),
    .B(_0780_),
    .Y(_0784_)
  );
  \$_AND_  _1386_ (
    .A(_0784_),
    .B(inst_type[1]),
    .Y(inst_jmp[0])
  );
  \$_AND_  _1387_ (
    .A(_0782_),
    .B(inst_jmp_bin[0]),
    .Y(_0785_)
  );
  \$_AND_  _1388_ (
    .A(_0785_),
    .B(_0780_),
    .Y(_0786_)
  );
  \$_AND_  _1389_ (
    .A(_0786_),
    .B(inst_type[1]),
    .Y(inst_jmp[1])
  );
  \$_AND_  _1390_ (
    .A(inst_jmp_bin[1]),
    .B(_0781_),
    .Y(_0787_)
  );
  \$_AND_  _1391_ (
    .A(_0787_),
    .B(_0780_),
    .Y(_0788_)
  );
  \$_AND_  _1392_ (
    .A(_0788_),
    .B(inst_type[1]),
    .Y(inst_jmp[2])
  );
  \$_AND_  _1393_ (
    .A(inst_jmp_bin[1]),
    .B(inst_jmp_bin[0]),
    .Y(_0789_)
  );
  \$_AND_  _1394_ (
    .A(_0789_),
    .B(_0780_),
    .Y(_0790_)
  );
  \$_AND_  _1395_ (
    .A(_0790_),
    .B(inst_type[1]),
    .Y(inst_jmp[3])
  );
  \$_AND_  _1396_ (
    .A(_0783_),
    .B(inst_jmp_bin[2]),
    .Y(_0791_)
  );
  \$_AND_  _1397_ (
    .A(_0791_),
    .B(inst_type[1]),
    .Y(inst_jmp[4])
  );
  \$_AND_  _1398_ (
    .A(_0785_),
    .B(inst_jmp_bin[2]),
    .Y(_0792_)
  );
  \$_AND_  _1399_ (
    .A(_0792_),
    .B(inst_type[1]),
    .Y(inst_jmp[5])
  );
  \$_AND_  _1400_ (
    .A(_0787_),
    .B(inst_jmp_bin[2]),
    .Y(_0793_)
  );
  \$_AND_  _1401_ (
    .A(_0793_),
    .B(inst_type[1]),
    .Y(inst_jmp[6])
  );
  \$_INV_  _1402_ (
    .A(_0783_),
    .Y(_0794_)
  );
  \$_INV_  _1403_ (
    .A(_0789_),
    .Y(_0795_)
  );
  \$_MUX_  _1404_ (
    .A(_0795_),
    .B(_0794_),
    .S(inst_jmp_bin[2]),
    .Y(_0796_)
  );
  \$_INV_  _1405_ (
    .A(_0792_),
    .Y(_0797_)
  );
  \$_INV_  _1406_ (
    .A(_0793_),
    .Y(_0798_)
  );
  \$_AND_  _1407_ (
    .A(_0798_),
    .B(_0797_),
    .Y(_0799_)
  );
  \$_AND_  _1408_ (
    .A(_0799_),
    .B(_0796_),
    .Y(_0800_)
  );
  \$_INV_  _1409_ (
    .A(_0784_),
    .Y(_0801_)
  );
  \$_AND_  _1410_ (
    .A(_0801_),
    .B(inst_type[1]),
    .Y(_0802_)
  );
  \$_INV_  _1411_ (
    .A(_0786_),
    .Y(_0803_)
  );
  \$_INV_  _1412_ (
    .A(_0788_),
    .Y(_0804_)
  );
  \$_AND_  _1413_ (
    .A(_0804_),
    .B(_0803_),
    .Y(_0805_)
  );
  \$_AND_  _1414_ (
    .A(_0805_),
    .B(_0802_),
    .Y(_0806_)
  );
  \$_AND_  _1415_ (
    .A(_0806_),
    .B(_0800_),
    .Y(inst_jmp[7])
  );
  \$_INV_  _1416_ (
    .A(_0719_),
    .Y(_1144_)
  );
  \$_INV_  _1417_ (
    .A(_0707_),
    .Y(_0807_)
  );
  \$_OR_  _1418_ (
    .A(_0720_),
    .B(_0807_),
    .Y(_1145_)
  );
  \$_INV_  _1419_ (
    .A(_0739_),
    .Y(_1146_)
  );
  \$_INV_  _1420_ (
    .A(_0689_),
    .Y(_0808_)
  );
  \$_INV_  _1421_ (
    .A(_0573_),
    .Y(_0809_)
  );
  \$_INV_  _1422_ (
    .A(_0579_),
    .Y(_0810_)
  );
  \$_MUX_  _1423_ (
    .A(_0810_),
    .B(_0809_),
    .S(_0576_),
    .Y(_0811_)
  );
  \$_AND_  _1424_ (
    .A(_0584_),
    .B(_0571_),
    .Y(_0812_)
  );
  \$_AND_  _1425_ (
    .A(_0812_),
    .B(_0576_),
    .Y(_0813_)
  );
  \$_AND_  _1426_ (
    .A(_0568_),
    .B(_0571_),
    .Y(_0814_)
  );
  \$_AND_  _1427_ (
    .A(_0814_),
    .B(_0576_),
    .Y(_0815_)
  );
  \$_OR_  _1428_ (
    .A(_0815_),
    .B(_0813_),
    .Y(_0816_)
  );
  \$_INV_  _1429_ (
    .A(_0816_),
    .Y(_0817_)
  );
  \$_AND_  _1430_ (
    .A(_0817_),
    .B(_0811_),
    .Y(_0818_)
  );
  \$_MUX_  _1431_ (
    .A(_0812_),
    .B(_0569_),
    .S(_0576_),
    .Y(_0819_)
  );
  \$_INV_  _1432_ (
    .A(_0819_),
    .Y(_0820_)
  );
  \$_INV_  _1433_ (
    .A(_0574_),
    .Y(_0821_)
  );
  \$_AND_  _1434_ (
    .A(_0577_),
    .B(_0572_),
    .Y(_0822_)
  );
  \$_INV_  _1435_ (
    .A(_0822_),
    .Y(_0823_)
  );
  \$_AND_  _1436_ (
    .A(_0823_),
    .B(_0821_),
    .Y(_0824_)
  );
  \$_AND_  _1437_ (
    .A(_0824_),
    .B(_0820_),
    .Y(_0825_)
  );
  \$_AND_  _1438_ (
    .A(_0825_),
    .B(_0818_),
    .Y(_0826_)
  );
  \$_INV_  _1439_ (
    .A(_0570_),
    .Y(_0827_)
  );
  \$_INV_  _1440_ (
    .A(_0578_),
    .Y(_0828_)
  );
  \$_AND_  _1441_ (
    .A(_0828_),
    .B(_0827_),
    .Y(_0829_)
  );
  \$_AND_  _1442_ (
    .A(_0829_),
    .B(_0587_),
    .Y(_0830_)
  );
  \$_AND_  _1443_ (
    .A(_0814_),
    .B(e_state[3]),
    .Y(_0831_)
  );
  \$_INV_  _1444_ (
    .A(_0831_),
    .Y(_0832_)
  );
  \$_AND_  _1445_ (
    .A(_0579_),
    .B(_0576_),
    .Y(_0833_)
  );
  \$_AND_  _1446_ (
    .A(_0585_),
    .B(_0576_),
    .Y(_0834_)
  );
  \$_OR_  _1447_ (
    .A(_0834_),
    .B(_0833_),
    .Y(_0835_)
  );
  \$_INV_  _1448_ (
    .A(_0835_),
    .Y(_0836_)
  );
  \$_AND_  _1449_ (
    .A(_0836_),
    .B(_0832_),
    .Y(_0837_)
  );
  \$_AND_  _1450_ (
    .A(_0837_),
    .B(_0830_),
    .Y(_0838_)
  );
  \$_AND_  _1451_ (
    .A(_0838_),
    .B(_0826_),
    .Y(_0839_)
  );
  \$_INV_  _1452_ (
    .A(exec_jmp),
    .Y(_0840_)
  );
  \$_INV_  _1453_ (
    .A(exec_src_wr),
    .Y(_0841_)
  );
  \$_AND_  _1454_ (
    .A(mdb_in[8]),
    .B(_0661_),
    .Y(_0842_)
  );
  \$_AND_  _1455_ (
    .A(_0842_),
    .B(mdb_in[9]),
    .Y(_0843_)
  );
  \$_INV_  _1456_ (
    .A(_0843_),
    .Y(_0844_)
  );
  \$_AND_  _1457_ (
    .A(_0628_),
    .B(_0661_),
    .Y(_0845_)
  );
  \$_AND_  _1458_ (
    .A(_0845_),
    .B(mdb_in[9]),
    .Y(_0846_)
  );
  \$_INV_  _1459_ (
    .A(_0846_),
    .Y(_0847_)
  );
  \$_AND_  _1460_ (
    .A(_0628_),
    .B(mdb_in[7]),
    .Y(_0848_)
  );
  \$_AND_  _1461_ (
    .A(_0848_),
    .B(mdb_in[9]),
    .Y(_0849_)
  );
  \$_INV_  _1462_ (
    .A(_0849_),
    .Y(_0850_)
  );
  \$_AND_  _1463_ (
    .A(_0850_),
    .B(_0847_),
    .Y(_0851_)
  );
  \$_AND_  _1464_ (
    .A(_0851_),
    .B(_0844_),
    .Y(_0852_)
  );
  \$_AND_  _1465_ (
    .A(_0845_),
    .B(_0637_),
    .Y(_0853_)
  );
  \$_AND_  _1466_ (
    .A(_0848_),
    .B(_0637_),
    .Y(_0854_)
  );
  \$_AND_  _1467_ (
    .A(_0842_),
    .B(_0637_),
    .Y(_0855_)
  );
  \$_AND_  _1468_ (
    .A(mdb_in[8]),
    .B(mdb_in[7]),
    .Y(_0856_)
  );
  \$_AND_  _1469_ (
    .A(_0856_),
    .B(_0637_),
    .Y(_0857_)
  );
  \$_INV_  _1470_ (
    .A(_0637_),
    .Y(_0858_)
  );
  \$_AND_  _1471_ (
    .A(_0858_),
    .B(_0852_),
    .Y(_0859_)
  );
  \$_AND_  _1472_ (
    .A(_0859_),
    .B(_0672_),
    .Y(_0860_)
  );
  \$_AND_  _1473_ (
    .A(_0860_),
    .B(_0660_),
    .Y(_0861_)
  );
  \$_OR_  _1474_ (
    .A(_0861_),
    .B(_0614_),
    .Y(_0862_)
  );
  \$_AND_  _1475_ (
    .A(_0862_),
    .B(_0609_),
    .Y(_0863_)
  );
  \$_AND_  _1476_ (
    .A(_0611_),
    .B(_0727_),
    .Y(_0864_)
  );
  \$_AND_  _1477_ (
    .A(_0843_),
    .B(_0672_),
    .Y(_0865_)
  );
  \$_AND_  _1478_ (
    .A(_0865_),
    .B(_0660_),
    .Y(_0866_)
  );
  \$_INV_  _1479_ (
    .A(_0866_),
    .Y(_0867_)
  );
  \$_AND_  _1480_ (
    .A(_0867_),
    .B(_0716_),
    .Y(_0868_)
  );
  \$_INV_  _1481_ (
    .A(mdb_in[4]),
    .Y(_0869_)
  );
  \$_AND_  _1482_ (
    .A(mdb_in[5]),
    .B(_0869_),
    .Y(_0870_)
  );
  \$_AND_  _1483_ (
    .A(_0870_),
    .B(_0644_),
    .Y(_0871_)
  );
  \$_AND_  _1484_ (
    .A(_0871_),
    .B(_0640_),
    .Y(_0872_)
  );
  \$_AND_  _1485_ (
    .A(_0872_),
    .B(_0652_),
    .Y(_0873_)
  );
  \$_AND_  _1486_ (
    .A(_0713_),
    .B(_0652_),
    .Y(_0874_)
  );
  \$_AND_  _1487_ (
    .A(_0657_),
    .B(_0874_),
    .Y(_0875_)
  );
  \$_OR_  _1488_ (
    .A(_0875_),
    .B(_0873_),
    .Y(_0876_)
  );
  \$_INV_  _1489_ (
    .A(_0876_),
    .Y(_0877_)
  );
  \$_AND_  _1490_ (
    .A(_0877_),
    .B(_0868_),
    .Y(_0878_)
  );
  \$_AND_  _1491_ (
    .A(_0944_),
    .B(_0864_),
    .Y(_0879_)
  );
  \$_OR_  _1492_ (
    .A(_0879_),
    .B(_0863_),
    .Y(_0880_)
  );
  \$_AND_  _1493_ (
    .A(_0880_),
    .B(_0841_),
    .Y(_0881_)
  );
  \$_AND_  _1494_ (
    .A(_0881_),
    .B(_0840_),
    .Y(_0882_)
  );
  \$_INV_  _1495_ (
    .A(_0882_),
    .Y(_0883_)
  );
  \$_INV_  _1496_ (
    .A(exec_dst_wr),
    .Y(_0884_)
  );
  \$_AND_  _1497_ (
    .A(_0580_),
    .B(_0884_),
    .Y(_0885_)
  );
  \$_AND_  _1498_ (
    .A(_0885_),
    .B(_0883_),
    .Y(_0886_)
  );
  \$_INV_  _1499_ (
    .A(_0886_),
    .Y(_0887_)
  );
  \$_AND_  _1500_ (
    .A(_0880_),
    .B(_0840_),
    .Y(_0888_)
  );
  \$_OR_  _1501_ (
    .A(_0888_),
    .B(_0821_),
    .Y(_0889_)
  );
  \$_OR_  _1502_ (
    .A(_0880_),
    .B(_0830_),
    .Y(_0890_)
  );
  \$_AND_  _1503_ (
    .A(_0890_),
    .B(_0836_),
    .Y(_0891_)
  );
  \$_AND_  _1504_ (
    .A(_0891_),
    .B(_0889_),
    .Y(_0892_)
  );
  \$_AND_  _1505_ (
    .A(_0892_),
    .B(_0887_),
    .Y(_0893_)
  );
  \$_INV_  _1506_ (
    .A(_0839_),
    .Y(_0894_)
  );
  \$_INV_  _1507_ (
    .A(_0863_),
    .Y(_0895_)
  );
  \$_INV_  _1508_ (
    .A(_0864_),
    .Y(_0896_)
  );
  \$_AND_  _1509_ (
    .A(_0669_),
    .B(_0711_),
    .Y(_0897_)
  );
  \$_AND_  _1510_ (
    .A(_0897_),
    .B(_0878_),
    .Y(_0898_)
  );
  \$_OR_  _1511_ (
    .A(_0898_),
    .B(_0648_),
    .Y(_0899_)
  );
  \$_OR_  _1512_ (
    .A(_0899_),
    .B(cpuoff),
    .Y(_0900_)
  );
  \$_OR_  _1513_ (
    .A(_0900_),
    .B(_0896_),
    .Y(_0901_)
  );
  \$_AND_  _1514_ (
    .A(_0901_),
    .B(_0895_),
    .Y(_0902_)
  );
  \$_INV_  _1515_ (
    .A(_0902_),
    .Y(_0903_)
  );
  \$_AND_  _1516_ (
    .A(_0903_),
    .B(_0841_),
    .Y(_0904_)
  );
  \$_INV_  _1517_ (
    .A(_0904_),
    .Y(_0905_)
  );
  \$_AND_  _1518_ (
    .A(_0884_),
    .B(_0840_),
    .Y(_0906_)
  );
  \$_AND_  _1519_ (
    .A(_0906_),
    .B(_0580_),
    .Y(_0907_)
  );
  \$_AND_  _1520_ (
    .A(_0907_),
    .B(_0905_),
    .Y(_0908_)
  );
  \$_INV_  _1521_ (
    .A(_0830_),
    .Y(_0909_)
  );
  \$_AND_  _1522_ (
    .A(_0902_),
    .B(_0909_),
    .Y(_0910_)
  );
  \$_AND_  _1523_ (
    .A(_0574_),
    .B(_0840_),
    .Y(_0911_)
  );
  \$_AND_  _1524_ (
    .A(_0911_),
    .B(_0902_),
    .Y(_0912_)
  );
  \$_INV_  _1525_ (
    .A(i_state[0]),
    .Y(_0913_)
  );
  \$_OR_  _1526_ (
    .A(inst_as[1]),
    .B(inst_as[4]),
    .Y(_0914_)
  );
  \$_OR_  _1527_ (
    .A(inst_as[5]),
    .B(inst_as[6]),
    .Y(_0915_)
  );
  \$_OR_  _1528_ (
    .A(_0915_),
    .B(_0914_),
    .Y(_0916_)
  );
  \$_INV_  _1529_ (
    .A(_0916_),
    .Y(_0917_)
  );
  \$_AND_  _1530_ (
    .A(_0917_),
    .B(i_state[4]),
    .Y(_0918_)
  );
  \$_INV_  _1531_ (
    .A(_0918_),
    .Y(_0919_)
  );
  \$_AND_  _1532_ (
    .A(_0919_),
    .B(_0913_),
    .Y(_0920_)
  );
  \$_INV_  _1533_ (
    .A(_0920_),
    .Y(_0921_)
  );
  \$_OR_  _1534_ (
    .A(_0921_),
    .B(exec_dext_rdy),
    .Y(_0922_)
  );
  \$_AND_  _1535_ (
    .A(_0922_),
    .B(_0831_),
    .Y(_0923_)
  );
  \$_INV_  _1536_ (
    .A(inst_ad[6]),
    .Y(_0924_)
  );
  \$_INV_  _1537_ (
    .A(inst_ad[4]),
    .Y(_0925_)
  );
  \$_INV_  _1538_ (
    .A(inst_ad[1]),
    .Y(_0926_)
  );
  \$_AND_  _1539_ (
    .A(_0926_),
    .B(_0925_),
    .Y(_0927_)
  );
  \$_AND_  _1540_ (
    .A(_0927_),
    .B(_0924_),
    .Y(_0928_)
  );
  \$_AND_  _1541_ (
    .A(_0928_),
    .B(_0822_),
    .Y(_0929_)
  );
  \$_AND_  _1542_ (
    .A(_0573_),
    .B(_0576_),
    .Y(_0930_)
  );
  \$_OR_  _1543_ (
    .A(_0815_),
    .B(_0930_),
    .Y(_0931_)
  );
  \$_OR_  _1544_ (
    .A(_0931_),
    .B(_0929_),
    .Y(_0932_)
  );
  \$_AND_  _1545_ (
    .A(_0916_),
    .B(i_state[4]),
    .Y(_0933_)
  );
  \$_INV_  _1546_ (
    .A(_0933_),
    .Y(_0934_)
  );
  \$_AND_  _1547_ (
    .A(_0934_),
    .B(_0834_),
    .Y(_0935_)
  );
  \$_OR_  _1548_ (
    .A(_0935_),
    .B(_0819_),
    .Y(_0936_)
  );
  \$_OR_  _1549_ (
    .A(_0936_),
    .B(_0932_),
    .Y(_0937_)
  );
  \$_OR_  _1550_ (
    .A(_0937_),
    .B(_0923_),
    .Y(_0938_)
  );
  \$_OR_  _1551_ (
    .A(_0938_),
    .B(_0912_),
    .Y(_0939_)
  );
  \$_OR_  _1552_ (
    .A(_0939_),
    .B(_0910_),
    .Y(_0940_)
  );
  \$_OR_  _1553_ (
    .A(_0940_),
    .B(_0908_),
    .Y(_0941_)
  );
  \$_AND_  _1554_ (
    .A(_0941_),
    .B(_0894_),
    .Y(e_state_nxt[0])
  );
  \$_INV_  _1555_ (
    .A(e_state_nxt[0]),
    .Y(_0942_)
  );
  \$_AND_  _1556_ (
    .A(_0711_),
    .B(_0673_),
    .Y(_0943_)
  );
  \$_AND_  _1557_ (
    .A(_0943_),
    .B(_0878_),
    .Y(_0944_)
  );
  \$_OR_  _1558_ (
    .A(_0944_),
    .B(cpuoff),
    .Y(_0945_)
  );
  \$_OR_  _1559_ (
    .A(_0945_),
    .B(_0896_),
    .Y(_0946_)
  );
  \$_AND_  _1560_ (
    .A(_0946_),
    .B(_0895_),
    .Y(_0947_)
  );
  \$_AND_  _1561_ (
    .A(_0841_),
    .B(_0840_),
    .Y(_0948_)
  );
  \$_AND_  _1562_ (
    .A(_0948_),
    .B(_0947_),
    .Y(_0949_)
  );
  \$_OR_  _1563_ (
    .A(_0949_),
    .B(exec_jmp),
    .Y(_0950_)
  );
  \$_OR_  _1564_ (
    .A(_0950_),
    .B(exec_dst_wr),
    .Y(_0951_)
  );
  \$_AND_  _1565_ (
    .A(_0951_),
    .B(_0580_),
    .Y(_0952_)
  );
  \$_INV_  _1566_ (
    .A(_0952_),
    .Y(_0953_)
  );
  \$_INV_  _1567_ (
    .A(_0947_),
    .Y(_0954_)
  );
  \$_AND_  _1568_ (
    .A(_0954_),
    .B(_0840_),
    .Y(_0955_)
  );
  \$_OR_  _1569_ (
    .A(_0955_),
    .B(_0821_),
    .Y(_0956_)
  );
  \$_AND_  _1570_ (
    .A(_0947_),
    .B(_0909_),
    .Y(_0957_)
  );
  \$_INV_  _1571_ (
    .A(_0957_),
    .Y(_0958_)
  );
  \$_AND_  _1572_ (
    .A(_0832_),
    .B(_0823_),
    .Y(_0959_)
  );
  \$_AND_  _1573_ (
    .A(_0959_),
    .B(_0820_),
    .Y(_0960_)
  );
  \$_AND_  _1574_ (
    .A(_0960_),
    .B(_0958_),
    .Y(_0961_)
  );
  \$_AND_  _1575_ (
    .A(_0961_),
    .B(_0956_),
    .Y(_0962_)
  );
  \$_AND_  _1576_ (
    .A(_0962_),
    .B(_0953_),
    .Y(_0963_)
  );
  \$_INV_  _1577_ (
    .A(_0878_),
    .Y(_0964_)
  );
  \$_OR_  _1578_ (
    .A(_0666_),
    .B(_0661_),
    .Y(_0965_)
  );
  \$_OR_  _1579_ (
    .A(_0965_),
    .B(_0668_),
    .Y(_0966_)
  );
  \$_OR_  _1580_ (
    .A(_0966_),
    .B(_0663_),
    .Y(_0967_)
  );
  \$_AND_  _1581_ (
    .A(_0867_),
    .B(_0967_),
    .Y(_0968_)
  );
  \$_AND_  _1582_ (
    .A(_0846_),
    .B(_0672_),
    .Y(_0969_)
  );
  \$_AND_  _1583_ (
    .A(_0969_),
    .B(_0660_),
    .Y(_0970_)
  );
  \$_INV_  _1584_ (
    .A(_0970_),
    .Y(_0971_)
  );
  \$_AND_  _1585_ (
    .A(_0849_),
    .B(_0672_),
    .Y(_0972_)
  );
  \$_AND_  _1586_ (
    .A(_0972_),
    .B(_0660_),
    .Y(_0973_)
  );
  \$_INV_  _1587_ (
    .A(_0973_),
    .Y(_0974_)
  );
  \$_AND_  _1588_ (
    .A(_0974_),
    .B(_0971_),
    .Y(_0975_)
  );
  \$_AND_  _1589_ (
    .A(_0975_),
    .B(_0968_),
    .Y(_0976_)
  );
  \$_AND_  _1590_ (
    .A(_0976_),
    .B(_0669_),
    .Y(_0977_)
  );
  \$_OR_  _1591_ (
    .A(_0977_),
    .B(_0964_),
    .Y(_0978_)
  );
  \$_AND_  _1592_ (
    .A(_0864_),
    .B(_0673_),
    .Y(_0979_)
  );
  \$_AND_  _1593_ (
    .A(_0979_),
    .B(_0895_),
    .Y(_0980_)
  );
  \$_AND_  _1594_ (
    .A(_0980_),
    .B(_0711_),
    .Y(_0981_)
  );
  \$_AND_  _1595_ (
    .A(_0981_),
    .B(_0978_),
    .Y(_0982_)
  );
  \$_OR_  _1596_ (
    .A(_0982_),
    .B(_0863_),
    .Y(_0983_)
  );
  \$_OR_  _1597_ (
    .A(_0983_),
    .B(exec_src_wr),
    .Y(_0984_)
  );
  \$_AND_  _1598_ (
    .A(_0984_),
    .B(_0906_),
    .Y(_0985_)
  );
  \$_OR_  _1599_ (
    .A(_0985_),
    .B(exec_dst_wr),
    .Y(_0986_)
  );
  \$_AND_  _1600_ (
    .A(_0986_),
    .B(_0580_),
    .Y(_0987_)
  );
  \$_AND_  _1601_ (
    .A(_0983_),
    .B(_0909_),
    .Y(_0988_)
  );
  \$_AND_  _1602_ (
    .A(_0983_),
    .B(_0911_),
    .Y(_0989_)
  );
  \$_OR_  _1603_ (
    .A(_0819_),
    .B(_0815_),
    .Y(_0990_)
  );
  \$_AND_  _1604_ (
    .A(_0933_),
    .B(_0834_),
    .Y(_0991_)
  );
  \$_OR_  _1605_ (
    .A(inst_so[5]),
    .B(inst_so[4]),
    .Y(_0992_)
  );
  \$_INV_  _1606_ (
    .A(_0992_),
    .Y(_0993_)
  );
  \$_INV_  _1607_ (
    .A(inst_so[6]),
    .Y(_0994_)
  );
  \$_AND_  _1608_ (
    .A(_0994_),
    .B(_0926_),
    .Y(_0995_)
  );
  \$_AND_  _1609_ (
    .A(_0995_),
    .B(_0993_),
    .Y(_0996_)
  );
  \$_AND_  _1610_ (
    .A(_0996_),
    .B(_0822_),
    .Y(_0997_)
  );
  \$_AND_  _1611_ (
    .A(_0997_),
    .B(_0928_),
    .Y(_0998_)
  );
  \$_OR_  _1612_ (
    .A(_0998_),
    .B(_0991_),
    .Y(_0999_)
  );
  \$_OR_  _1613_ (
    .A(_0999_),
    .B(_0990_),
    .Y(_1000_)
  );
  \$_OR_  _1614_ (
    .A(_1000_),
    .B(_0989_),
    .Y(_1001_)
  );
  \$_OR_  _1615_ (
    .A(_1001_),
    .B(_0988_),
    .Y(_1002_)
  );
  \$_OR_  _1616_ (
    .A(_1002_),
    .B(_0987_),
    .Y(_1003_)
  );
  \$_OR_  _1617_ (
    .A(_1003_),
    .B(_0839_),
    .Y(e_state_nxt[1])
  );
  \$_OR_  _1618_ (
    .A(e_state_nxt[1]),
    .B(_0963_),
    .Y(_1004_)
  );
  \$_OR_  _1619_ (
    .A(_1004_),
    .B(_0942_),
    .Y(_1005_)
  );
  \$_OR_  _1620_ (
    .A(_1005_),
    .B(_0893_),
    .Y(_1006_)
  );
  \$_AND_  _1621_ (
    .A(_1006_),
    .B(_0808_),
    .Y(_1007_)
  );
  \$_AND_  _1622_ (
    .A(_0611_),
    .B(dbg_halt_st),
    .Y(_1008_)
  );
  \$_OR_  _1623_ (
    .A(pmem_busy),
    .B(pc_sw_wr),
    .Y(_1009_)
  );
  \$_OR_  _1624_ (
    .A(_1009_),
    .B(_1008_),
    .Y(_1010_)
  );
  \$_OR_  _1625_ (
    .A(_1010_),
    .B(_1142_[15]),
    .Y(_1011_)
  );
  \$_OR_  _1626_ (
    .A(_1011_),
    .B(_1007_),
    .Y(mb_en)
  );
  \$_AND_  _1627_ (
    .A(_0583_),
    .B(inst_irq_rst),
    .Y(_0011_)
  );
  \$_INV_  _1628_ (
    .A(_0593_),
    .Y(_1012_)
  );
  \$_OR_  _1629_ (
    .A(_1012_),
    .B(irq[1]),
    .Y(_1013_)
  );
  \$_INV_  _1630_ (
    .A(irq[2]),
    .Y(_1014_)
  );
  \$_INV_  _1631_ (
    .A(irq[3]),
    .Y(_1015_)
  );
  \$_AND_  _1632_ (
    .A(_1015_),
    .B(_1014_),
    .Y(_1016_)
  );
  \$_AND_  _1633_ (
    .A(_1016_),
    .B(_1013_),
    .Y(_1017_)
  );
  \$_OR_  _1634_ (
    .A(_1017_),
    .B(irq[3]),
    .Y(_1018_)
  );
  \$_INV_  _1635_ (
    .A(irq[4]),
    .Y(_1019_)
  );
  \$_INV_  _1636_ (
    .A(irq[5]),
    .Y(_1020_)
  );
  \$_AND_  _1637_ (
    .A(_1020_),
    .B(_1019_),
    .Y(_1021_)
  );
  \$_AND_  _1638_ (
    .A(_1021_),
    .B(_1018_),
    .Y(_1022_)
  );
  \$_OR_  _1639_ (
    .A(_1022_),
    .B(irq[5]),
    .Y(_1023_)
  );
  \$_INV_  _1640_ (
    .A(irq[6]),
    .Y(_1024_)
  );
  \$_INV_  _1641_ (
    .A(irq[7]),
    .Y(_1025_)
  );
  \$_AND_  _1642_ (
    .A(_1025_),
    .B(_1024_),
    .Y(_1026_)
  );
  \$_AND_  _1643_ (
    .A(_1026_),
    .B(_1023_),
    .Y(_1027_)
  );
  \$_OR_  _1644_ (
    .A(_1027_),
    .B(irq[7]),
    .Y(_1028_)
  );
  \$_INV_  _1645_ (
    .A(irq[8]),
    .Y(_1029_)
  );
  \$_INV_  _1646_ (
    .A(irq[9]),
    .Y(_1030_)
  );
  \$_AND_  _1647_ (
    .A(_1030_),
    .B(_1029_),
    .Y(_1031_)
  );
  \$_AND_  _1648_ (
    .A(_1031_),
    .B(_1028_),
    .Y(_1032_)
  );
  \$_OR_  _1649_ (
    .A(_1032_),
    .B(irq[9]),
    .Y(_1033_)
  );
  \$_INV_  _1650_ (
    .A(irq[11]),
    .Y(_1034_)
  );
  \$_INV_  _1651_ (
    .A(_0601_),
    .Y(_1035_)
  );
  \$_AND_  _1652_ (
    .A(_1035_),
    .B(_1034_),
    .Y(_1036_)
  );
  \$_AND_  _1653_ (
    .A(_1036_),
    .B(_1033_),
    .Y(_1037_)
  );
  \$_OR_  _1654_ (
    .A(_1037_),
    .B(irq[11]),
    .Y(_1038_)
  );
  \$_INV_  _1655_ (
    .A(irq[12]),
    .Y(_1039_)
  );
  \$_INV_  _1656_ (
    .A(irq[13]),
    .Y(_1040_)
  );
  \$_AND_  _1657_ (
    .A(_1040_),
    .B(_1039_),
    .Y(_1041_)
  );
  \$_AND_  _1658_ (
    .A(_1041_),
    .B(_1038_),
    .Y(_1042_)
  );
  \$_OR_  _1659_ (
    .A(_1042_),
    .B(irq[13]),
    .Y(_1043_)
  );
  \$_INV_  _1660_ (
    .A(nmi_pnd),
    .Y(_1044_)
  );
  \$_AND_  _1661_ (
    .A(_0614_),
    .B(_1044_),
    .Y(_1045_)
  );
  \$_AND_  _1662_ (
    .A(_1045_),
    .B(_1043_),
    .Y(_1046_)
  );
  \$_AND_  _1663_ (
    .A(_0672_),
    .B(irq_addr[1]),
    .Y(_1047_)
  );
  \$_OR_  _1664_ (
    .A(_1047_),
    .B(_1046_),
    .Y(_0019_[0])
  );
  \$_OR_  _1665_ (
    .A(_1012_),
    .B(irq[2]),
    .Y(_1048_)
  );
  \$_OR_  _1666_ (
    .A(_1048_),
    .B(irq[3]),
    .Y(_1049_)
  );
  \$_AND_  _1667_ (
    .A(_1021_),
    .B(_1024_),
    .Y(_1050_)
  );
  \$_AND_  _1668_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_1051_)
  );
  \$_OR_  _1669_ (
    .A(_1051_),
    .B(irq[6]),
    .Y(_1052_)
  );
  \$_OR_  _1670_ (
    .A(_1052_),
    .B(irq[7]),
    .Y(_1053_)
  );
  \$_AND_  _1671_ (
    .A(_1031_),
    .B(_1035_),
    .Y(_1054_)
  );
  \$_AND_  _1672_ (
    .A(_1054_),
    .B(_1053_),
    .Y(_1055_)
  );
  \$_OR_  _1673_ (
    .A(_1055_),
    .B(_0601_),
    .Y(_1056_)
  );
  \$_OR_  _1674_ (
    .A(_1056_),
    .B(irq[11]),
    .Y(_1057_)
  );
  \$_AND_  _1675_ (
    .A(_1039_),
    .B(_1044_),
    .Y(_1058_)
  );
  \$_AND_  _1676_ (
    .A(_1058_),
    .B(_1040_),
    .Y(_1059_)
  );
  \$_AND_  _1677_ (
    .A(_1059_),
    .B(_1057_),
    .Y(_1060_)
  );
  \$_OR_  _1678_ (
    .A(_1060_),
    .B(nmi_pnd),
    .Y(_1061_)
  );
  \$_MUX_  _1679_ (
    .A(_1061_),
    .B(irq_addr[2]),
    .S(_0672_),
    .Y(_0019_[1])
  );
  \$_INV_  _1680_ (
    .A(_0596_),
    .Y(_1062_)
  );
  \$_OR_  _1681_ (
    .A(_1062_),
    .B(irq[4]),
    .Y(_1063_)
  );
  \$_OR_  _1682_ (
    .A(_1063_),
    .B(irq[5]),
    .Y(_1064_)
  );
  \$_OR_  _1683_ (
    .A(_1064_),
    .B(irq[6]),
    .Y(_1065_)
  );
  \$_OR_  _1684_ (
    .A(_1065_),
    .B(irq[7]),
    .Y(_1066_)
  );
  \$_INV_  _1685_ (
    .A(_0602_),
    .Y(_1067_)
  );
  \$_AND_  _1686_ (
    .A(_1054_),
    .B(_1067_),
    .Y(_1068_)
  );
  \$_AND_  _1687_ (
    .A(_1068_),
    .B(_1066_),
    .Y(_1069_)
  );
  \$_OR_  _1688_ (
    .A(_1069_),
    .B(irq[12]),
    .Y(_1070_)
  );
  \$_OR_  _1689_ (
    .A(_1070_),
    .B(irq[13]),
    .Y(_1071_)
  );
  \$_OR_  _1690_ (
    .A(_1071_),
    .B(nmi_pnd),
    .Y(_1072_)
  );
  \$_MUX_  _1691_ (
    .A(_1072_),
    .B(irq_addr[3]),
    .S(_0672_),
    .Y(_0019_[2])
  );
  \$_INV_  _1692_ (
    .A(_0600_),
    .Y(_1073_)
  );
  \$_OR_  _1693_ (
    .A(_1073_),
    .B(irq[8]),
    .Y(_1074_)
  );
  \$_OR_  _1694_ (
    .A(_1074_),
    .B(irq[9]),
    .Y(_1075_)
  );
  \$_OR_  _1695_ (
    .A(_1075_),
    .B(_0601_),
    .Y(_1076_)
  );
  \$_OR_  _1696_ (
    .A(_1076_),
    .B(irq[11]),
    .Y(_1077_)
  );
  \$_OR_  _1697_ (
    .A(_1077_),
    .B(irq[12]),
    .Y(_1078_)
  );
  \$_OR_  _1698_ (
    .A(_1078_),
    .B(irq[13]),
    .Y(_1079_)
  );
  \$_OR_  _1699_ (
    .A(_1079_),
    .B(nmi_pnd),
    .Y(_1080_)
  );
  \$_MUX_  _1700_ (
    .A(_1080_),
    .B(irq_addr[4]),
    .S(_0672_),
    .Y(_0019_[3])
  );
  \$_OR_  _1701_ (
    .A(_0614_),
    .B(decode_noirq),
    .Y(_1081_)
  );
  \$_INV_  _1702_ (
    .A(_1081_),
    .Y(_1082_)
  );
  \$_OR_  _1703_ (
    .A(_0714_),
    .B(_0640_),
    .Y(_1083_)
  );
  \$_AND_  _1704_ (
    .A(_0871_),
    .B(_0709_),
    .Y(_1084_)
  );
  \$_INV_  _1705_ (
    .A(_1084_),
    .Y(_1085_)
  );
  \$_AND_  _1706_ (
    .A(_1085_),
    .B(_1083_),
    .Y(_1086_)
  );
  \$_AND_  _1707_ (
    .A(_0647_),
    .B(_0709_),
    .Y(_1087_)
  );
  \$_INV_  _1708_ (
    .A(_1087_),
    .Y(_1088_)
  );
  \$_AND_  _1709_ (
    .A(_0645_),
    .B(_0869_),
    .Y(_1089_)
  );
  \$_AND_  _1710_ (
    .A(_1089_),
    .B(_0644_),
    .Y(_1090_)
  );
  \$_INV_  _1711_ (
    .A(_1090_),
    .Y(_1091_)
  );
  \$_OR_  _1712_ (
    .A(_1091_),
    .B(_0640_),
    .Y(_1092_)
  );
  \$_AND_  _1713_ (
    .A(_1092_),
    .B(_1088_),
    .Y(_1093_)
  );
  \$_AND_  _1714_ (
    .A(_1093_),
    .B(_1086_),
    .Y(_1094_)
  );
  \$_AND_  _1715_ (
    .A(_0657_),
    .B(_0632_),
    .Y(_1095_)
  );
  \$_INV_  _1716_ (
    .A(_1095_),
    .Y(_1096_)
  );
  \$_AND_  _1717_ (
    .A(_0872_),
    .B(_0632_),
    .Y(_1097_)
  );
  \$_INV_  _1718_ (
    .A(_1097_),
    .Y(_1098_)
  );
  \$_AND_  _1719_ (
    .A(_1098_),
    .B(_1096_),
    .Y(_1099_)
  );
  \$_AND_  _1720_ (
    .A(_1099_),
    .B(_1094_),
    .Y(_1100_)
  );
  \$_OR_  _1721_ (
    .A(_1100_),
    .B(_1082_),
    .Y(_1101_)
  );
  \$_AND_  _1722_ (
    .A(_0656_),
    .B(_0709_),
    .Y(_1102_)
  );
  \$_OR_  _1723_ (
    .A(_1102_),
    .B(_1087_),
    .Y(_1103_)
  );
  \$_INV_  _1724_ (
    .A(_0644_),
    .Y(_1104_)
  );
  \$_AND_  _1725_ (
    .A(_1081_),
    .B(_1104_),
    .Y(_1105_)
  );
  \$_INV_  _1726_ (
    .A(_1105_),
    .Y(_1106_)
  );
  \$_MUX_  _1727_ (
    .A(inst_sext[0]),
    .B(mdb_in[0]),
    .S(_0933_),
    .Y(_1107_)
  );
  \$_AND_  _1728_ (
    .A(_1107_),
    .B(_1106_),
    .Y(_1108_)
  );
  \$_MUX_  _1729_ (
    .A(_1103_),
    .B(_1108_),
    .S(_1101_),
    .Y(_0014_[0])
  );
  \$_INV_  _1730_ (
    .A(_1101_),
    .Y(_1109_)
  );
  \$_AND_  _1731_ (
    .A(_0746_),
    .B(_0741_),
    .Y(_1110_)
  );
  \$_AND_  _1732_ (
    .A(_1110_),
    .B(_0723_),
    .Y(_1111_)
  );
  \$_INV_  _1733_ (
    .A(inst_as[4]),
    .Y(_1112_)
  );
  \$_AND_  _1734_ (
    .A(i_state[4]),
    .B(_1112_),
    .Y(_1113_)
  );
  \$_AND_  _1735_ (
    .A(_1113_),
    .B(inst_ad[4]),
    .Y(_1114_)
  );
  \$_INV_  _1736_ (
    .A(_1114_),
    .Y(_1115_)
  );
  \$_OR_  _1737_ (
    .A(_1115_),
    .B(_1111_),
    .Y(_1116_)
  );
  \$_AND_  _1738_ (
    .A(i_state[4]),
    .B(inst_as[4]),
    .Y(_1117_)
  );
  \$_AND_  _1739_ (
    .A(i_state[0]),
    .B(inst_ad[4]),
    .Y(_1118_)
  );
  \$_OR_  _1740_ (
    .A(_1118_),
    .B(_1117_),
    .Y(_1119_)
  );
  \$_INV_  _1741_ (
    .A(_1119_),
    .Y(_1120_)
  );
  \$_AND_  _1742_ (
    .A(_1120_),
    .B(_1116_),
    .Y(_1121_)
  );
  \$_XOR_  _1743_ (
    .A(_1121_),
    .B(mdb_in[10]),
    .Y(_1122_)
  );
  \$_OR_  _1744_ (
    .A(_1121_),
    .B(_0637_),
    .Y(_1123_)
  );
  \$_XOR_  _1745_ (
    .A(_1121_),
    .B(mdb_in[9]),
    .Y(_1124_)
  );
  \$_OR_  _1746_ (
    .A(_1121_),
    .B(_0628_),
    .Y(_1125_)
  );
  \$_XOR_  _1747_ (
    .A(_1121_),
    .B(mdb_in[8]),
    .Y(_1126_)
  );
  \$_OR_  _1748_ (
    .A(_1121_),
    .B(_0661_),
    .Y(_1127_)
  );
  \$_XOR_  _1749_ (
    .A(_1121_),
    .B(mdb_in[7]),
    .Y(_1128_)
  );
  \$_INV_  _1750_ (
    .A(mdb_in[6]),
    .Y(_1129_)
  );
  \$_OR_  _1751_ (
    .A(_1121_),
    .B(_1129_),
    .Y(_1130_)
  );
  \$_XOR_  _1752_ (
    .A(_1121_),
    .B(mdb_in[6]),
    .Y(_1131_)
  );
  \$_OR_  _1753_ (
    .A(_1121_),
    .B(_0645_),
    .Y(_1132_)
  );
  \$_XOR_  _1754_ (
    .A(_1121_),
    .B(mdb_in[5]),
    .Y(_1133_)
  );
  \$_OR_  _1755_ (
    .A(_1121_),
    .B(_0869_),
    .Y(_1134_)
  );
  \$_XOR_  _1756_ (
    .A(_1121_),
    .B(mdb_in[4]),
    .Y(_1135_)
  );
  \$_OR_  _1757_ (
    .A(_1121_),
    .B(_0591_),
    .Y(_1136_)
  );
  \$_XOR_  _1758_ (
    .A(_1121_),
    .B(mdb_in[3]),
    .Y(_1137_)
  );
  \$_OR_  _1759_ (
    .A(_1121_),
    .B(_0624_),
    .Y(_1138_)
  );
  \$_XOR_  _1760_ (
    .A(_1121_),
    .B(mdb_in[2]),
    .Y(_1139_)
  );
  \$_OR_  _1761_ (
    .A(_1121_),
    .B(_0636_),
    .Y(_1140_)
  );
  \$_OR_  _1762_ (
    .A(_1140_),
    .B(_1139_),
    .Y(_1141_)
  );
  \$_AND_  _1763_ (
    .A(_1141_),
    .B(_1138_),
    .Y(_0020_)
  );
  \$_OR_  _1764_ (
    .A(_0020_),
    .B(_1137_),
    .Y(_0021_)
  );
  \$_AND_  _1765_ (
    .A(_0021_),
    .B(_1136_),
    .Y(_0022_)
  );
  \$_OR_  _1766_ (
    .A(_0022_),
    .B(_1135_),
    .Y(_0023_)
  );
  \$_AND_  _1767_ (
    .A(_0023_),
    .B(_1134_),
    .Y(_0024_)
  );
  \$_OR_  _1768_ (
    .A(_0024_),
    .B(_1133_),
    .Y(_0025_)
  );
  \$_AND_  _1769_ (
    .A(_0025_),
    .B(_1132_),
    .Y(_0026_)
  );
  \$_OR_  _1770_ (
    .A(_0026_),
    .B(_1131_),
    .Y(_0027_)
  );
  \$_AND_  _1771_ (
    .A(_0027_),
    .B(_1130_),
    .Y(_0028_)
  );
  \$_OR_  _1772_ (
    .A(_0028_),
    .B(_1128_),
    .Y(_0029_)
  );
  \$_AND_  _1773_ (
    .A(_0029_),
    .B(_1127_),
    .Y(_0030_)
  );
  \$_OR_  _1774_ (
    .A(_0030_),
    .B(_1126_),
    .Y(_0031_)
  );
  \$_AND_  _1775_ (
    .A(_0031_),
    .B(_1125_),
    .Y(_0032_)
  );
  \$_OR_  _1776_ (
    .A(_0032_),
    .B(_1124_),
    .Y(_0033_)
  );
  \$_AND_  _1777_ (
    .A(_0033_),
    .B(_1123_),
    .Y(_0034_)
  );
  \$_XOR_  _1778_ (
    .A(_0034_),
    .B(_1122_),
    .Y(_0035_)
  );
  \$_MUX_  _1779_ (
    .A(_0035_),
    .B(inst_sext[10]),
    .S(_0934_),
    .Y(_0036_)
  );
  \$_MUX_  _1780_ (
    .A(_0036_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0037_)
  );
  \$_MUX_  _1781_ (
    .A(_0037_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[10])
  );
  \$_XOR_  _1782_ (
    .A(_1121_),
    .B(mdb_in[11]),
    .Y(_0038_)
  );
  \$_OR_  _1783_ (
    .A(_1121_),
    .B(_0623_),
    .Y(_0039_)
  );
  \$_OR_  _1784_ (
    .A(_0034_),
    .B(_1122_),
    .Y(_0040_)
  );
  \$_AND_  _1785_ (
    .A(_0040_),
    .B(_0039_),
    .Y(_0041_)
  );
  \$_XOR_  _1786_ (
    .A(_0041_),
    .B(_0038_),
    .Y(_0042_)
  );
  \$_MUX_  _1787_ (
    .A(_0042_),
    .B(inst_sext[11]),
    .S(_0934_),
    .Y(_0043_)
  );
  \$_MUX_  _1788_ (
    .A(_0043_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0044_)
  );
  \$_MUX_  _1789_ (
    .A(_0044_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[11])
  );
  \$_XOR_  _1790_ (
    .A(_1121_),
    .B(mdb_in[12]),
    .Y(_0045_)
  );
  \$_OR_  _1791_ (
    .A(_1121_),
    .B(_0590_),
    .Y(_0046_)
  );
  \$_OR_  _1792_ (
    .A(_0041_),
    .B(_0038_),
    .Y(_0047_)
  );
  \$_AND_  _1793_ (
    .A(_0047_),
    .B(_0046_),
    .Y(_0048_)
  );
  \$_XOR_  _1794_ (
    .A(_0048_),
    .B(_0045_),
    .Y(_0049_)
  );
  \$_MUX_  _1795_ (
    .A(_0049_),
    .B(inst_sext[12]),
    .S(_0934_),
    .Y(_0050_)
  );
  \$_MUX_  _1796_ (
    .A(_0050_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0051_)
  );
  \$_MUX_  _1797_ (
    .A(_0051_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[12])
  );
  \$_XOR_  _1798_ (
    .A(_1121_),
    .B(mdb_in[13]),
    .Y(_0052_)
  );
  \$_INV_  _1799_ (
    .A(mdb_in[12]),
    .Y(_0053_)
  );
  \$_OR_  _1800_ (
    .A(_1121_),
    .B(_0053_),
    .Y(_0054_)
  );
  \$_OR_  _1801_ (
    .A(_0048_),
    .B(_0045_),
    .Y(_0055_)
  );
  \$_AND_  _1802_ (
    .A(_0055_),
    .B(_0054_),
    .Y(_0056_)
  );
  \$_XOR_  _1803_ (
    .A(_0056_),
    .B(_0052_),
    .Y(_0057_)
  );
  \$_MUX_  _1804_ (
    .A(_0057_),
    .B(inst_sext[13]),
    .S(_0934_),
    .Y(_0058_)
  );
  \$_MUX_  _1805_ (
    .A(_0058_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0059_)
  );
  \$_MUX_  _1806_ (
    .A(_0059_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[13])
  );
  \$_XOR_  _1807_ (
    .A(_1121_),
    .B(mdb_in[14]),
    .Y(_0060_)
  );
  \$_OR_  _1808_ (
    .A(_1121_),
    .B(_0616_),
    .Y(_0061_)
  );
  \$_OR_  _1809_ (
    .A(_0056_),
    .B(_0052_),
    .Y(_0062_)
  );
  \$_AND_  _1810_ (
    .A(_0062_),
    .B(_0061_),
    .Y(_0063_)
  );
  \$_XOR_  _1811_ (
    .A(_0063_),
    .B(_0060_),
    .Y(_0064_)
  );
  \$_MUX_  _1812_ (
    .A(_0064_),
    .B(inst_sext[14]),
    .S(_0934_),
    .Y(_0065_)
  );
  \$_MUX_  _1813_ (
    .A(_0065_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0066_)
  );
  \$_MUX_  _1814_ (
    .A(_0066_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[14])
  );
  \$_XOR_  _1815_ (
    .A(_1121_),
    .B(mdb_in[15]),
    .Y(_0067_)
  );
  \$_OR_  _1816_ (
    .A(_1121_),
    .B(_0617_),
    .Y(_0068_)
  );
  \$_OR_  _1817_ (
    .A(_0063_),
    .B(_0060_),
    .Y(_0069_)
  );
  \$_AND_  _1818_ (
    .A(_0069_),
    .B(_0068_),
    .Y(_0070_)
  );
  \$_XOR_  _1819_ (
    .A(_0070_),
    .B(_0067_),
    .Y(_0071_)
  );
  \$_MUX_  _1820_ (
    .A(_0071_),
    .B(inst_sext[15]),
    .S(_0934_),
    .Y(_0072_)
  );
  \$_MUX_  _1821_ (
    .A(_0072_),
    .B(mdb_in[9]),
    .S(_1105_),
    .Y(_0073_)
  );
  \$_MUX_  _1822_ (
    .A(_0073_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[15])
  );
  \$_OR_  _1823_ (
    .A(_1084_),
    .B(_1102_),
    .Y(_0074_)
  );
  \$_XOR_  _1824_ (
    .A(_1121_),
    .B(_0636_),
    .Y(_0075_)
  );
  \$_MUX_  _1825_ (
    .A(_0075_),
    .B(inst_sext[1]),
    .S(_0934_),
    .Y(_0076_)
  );
  \$_MUX_  _1826_ (
    .A(_0076_),
    .B(mdb_in[0]),
    .S(_1105_),
    .Y(_0077_)
  );
  \$_MUX_  _1827_ (
    .A(_0077_),
    .B(_0074_),
    .S(_1109_),
    .Y(_0014_[1])
  );
  \$_OR_  _1828_ (
    .A(_1102_),
    .B(_1097_),
    .Y(_0078_)
  );
  \$_XOR_  _1829_ (
    .A(_1140_),
    .B(_1139_),
    .Y(_0079_)
  );
  \$_MUX_  _1830_ (
    .A(_0079_),
    .B(inst_sext[2]),
    .S(_0934_),
    .Y(_0080_)
  );
  \$_MUX_  _1831_ (
    .A(_0080_),
    .B(mdb_in[1]),
    .S(_1105_),
    .Y(_0081_)
  );
  \$_MUX_  _1832_ (
    .A(_0081_),
    .B(_0078_),
    .S(_1109_),
    .Y(_0014_[2])
  );
  \$_OR_  _1833_ (
    .A(_1102_),
    .B(_1095_),
    .Y(_0082_)
  );
  \$_AND_  _1834_ (
    .A(_1109_),
    .B(_1098_),
    .Y(_0083_)
  );
  \$_AND_  _1835_ (
    .A(_0083_),
    .B(_0082_),
    .Y(_0084_)
  );
  \$_XOR_  _1836_ (
    .A(_0020_),
    .B(_1137_),
    .Y(_0085_)
  );
  \$_MUX_  _1837_ (
    .A(_0085_),
    .B(inst_sext[3]),
    .S(_0934_),
    .Y(_0086_)
  );
  \$_MUX_  _1838_ (
    .A(_0086_),
    .B(mdb_in[2]),
    .S(_1105_),
    .Y(_0087_)
  );
  \$_AND_  _1839_ (
    .A(_0087_),
    .B(_1101_),
    .Y(_0088_)
  );
  \$_OR_  _1840_ (
    .A(_0088_),
    .B(_0084_),
    .Y(_0014_[3])
  );
  \$_XOR_  _1841_ (
    .A(_0022_),
    .B(_1135_),
    .Y(_0089_)
  );
  \$_MUX_  _1842_ (
    .A(_0089_),
    .B(inst_sext[4]),
    .S(_0934_),
    .Y(_0090_)
  );
  \$_MUX_  _1843_ (
    .A(_0090_),
    .B(mdb_in[3]),
    .S(_1105_),
    .Y(_0091_)
  );
  \$_MUX_  _1844_ (
    .A(_0091_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[4])
  );
  \$_XOR_  _1845_ (
    .A(_0024_),
    .B(_1133_),
    .Y(_0092_)
  );
  \$_MUX_  _1846_ (
    .A(_0092_),
    .B(inst_sext[5]),
    .S(_0934_),
    .Y(_0093_)
  );
  \$_MUX_  _1847_ (
    .A(_0093_),
    .B(mdb_in[4]),
    .S(_1105_),
    .Y(_0094_)
  );
  \$_MUX_  _1848_ (
    .A(_0094_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[5])
  );
  \$_XOR_  _1849_ (
    .A(_0026_),
    .B(_1131_),
    .Y(_0095_)
  );
  \$_MUX_  _1850_ (
    .A(_0095_),
    .B(inst_sext[6]),
    .S(_0934_),
    .Y(_0096_)
  );
  \$_MUX_  _1851_ (
    .A(_0096_),
    .B(mdb_in[5]),
    .S(_1105_),
    .Y(_0097_)
  );
  \$_MUX_  _1852_ (
    .A(_0097_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[6])
  );
  \$_XOR_  _1853_ (
    .A(_0028_),
    .B(_1128_),
    .Y(_0098_)
  );
  \$_MUX_  _1854_ (
    .A(_0098_),
    .B(inst_sext[7]),
    .S(_0934_),
    .Y(_0099_)
  );
  \$_MUX_  _1855_ (
    .A(_0099_),
    .B(mdb_in[6]),
    .S(_1105_),
    .Y(_0100_)
  );
  \$_MUX_  _1856_ (
    .A(_0100_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[7])
  );
  \$_XOR_  _1857_ (
    .A(_0030_),
    .B(_1126_),
    .Y(_0101_)
  );
  \$_MUX_  _1858_ (
    .A(_0101_),
    .B(inst_sext[8]),
    .S(_0934_),
    .Y(_0102_)
  );
  \$_MUX_  _1859_ (
    .A(_0102_),
    .B(mdb_in[7]),
    .S(_1105_),
    .Y(_0103_)
  );
  \$_MUX_  _1860_ (
    .A(_0103_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[8])
  );
  \$_XOR_  _1861_ (
    .A(_0032_),
    .B(_1124_),
    .Y(_0104_)
  );
  \$_MUX_  _1862_ (
    .A(_0104_),
    .B(inst_sext[9]),
    .S(_0934_),
    .Y(_0105_)
  );
  \$_MUX_  _1863_ (
    .A(_0105_),
    .B(mdb_in[8]),
    .S(_1105_),
    .Y(_0106_)
  );
  \$_MUX_  _1864_ (
    .A(_0106_),
    .B(_1102_),
    .S(_1109_),
    .Y(_0014_[9])
  );
  \$_MUX_  _1865_ (
    .A(inst_dext[0]),
    .B(mdb_in[0]),
    .S(i_state[0]),
    .Y(_0107_)
  );
  \$_MUX_  _1866_ (
    .A(_0107_),
    .B(mdb_in[0]),
    .S(_0918_),
    .Y(_0010_[0])
  );
  \$_MUX_  _1867_ (
    .A(_0035_),
    .B(inst_dext[10]),
    .S(_0913_),
    .Y(_0108_)
  );
  \$_MUX_  _1868_ (
    .A(_0108_),
    .B(_0035_),
    .S(_0918_),
    .Y(_0010_[10])
  );
  \$_MUX_  _1869_ (
    .A(_0042_),
    .B(inst_dext[11]),
    .S(_0913_),
    .Y(_0109_)
  );
  \$_MUX_  _1870_ (
    .A(_0109_),
    .B(_0042_),
    .S(_0918_),
    .Y(_0010_[11])
  );
  \$_MUX_  _1871_ (
    .A(_0049_),
    .B(inst_dext[12]),
    .S(_0913_),
    .Y(_0110_)
  );
  \$_MUX_  _1872_ (
    .A(_0110_),
    .B(_0049_),
    .S(_0918_),
    .Y(_0010_[12])
  );
  \$_MUX_  _1873_ (
    .A(_0057_),
    .B(inst_dext[13]),
    .S(_0913_),
    .Y(_0111_)
  );
  \$_MUX_  _1874_ (
    .A(_0111_),
    .B(_0057_),
    .S(_0918_),
    .Y(_0010_[13])
  );
  \$_MUX_  _1875_ (
    .A(_0064_),
    .B(inst_dext[14]),
    .S(_0913_),
    .Y(_0112_)
  );
  \$_MUX_  _1876_ (
    .A(_0112_),
    .B(_0064_),
    .S(_0918_),
    .Y(_0010_[14])
  );
  \$_MUX_  _1877_ (
    .A(_0071_),
    .B(inst_dext[15]),
    .S(_0913_),
    .Y(_0113_)
  );
  \$_MUX_  _1878_ (
    .A(_0113_),
    .B(_0071_),
    .S(_0918_),
    .Y(_0010_[15])
  );
  \$_MUX_  _1879_ (
    .A(_0075_),
    .B(inst_dext[1]),
    .S(_0913_),
    .Y(_0114_)
  );
  \$_MUX_  _1880_ (
    .A(_0114_),
    .B(_0075_),
    .S(_0918_),
    .Y(_0010_[1])
  );
  \$_MUX_  _1881_ (
    .A(_0079_),
    .B(inst_dext[2]),
    .S(_0913_),
    .Y(_0115_)
  );
  \$_MUX_  _1882_ (
    .A(_0115_),
    .B(_0079_),
    .S(_0918_),
    .Y(_0010_[2])
  );
  \$_MUX_  _1883_ (
    .A(_0085_),
    .B(inst_dext[3]),
    .S(_0913_),
    .Y(_0116_)
  );
  \$_MUX_  _1884_ (
    .A(_0116_),
    .B(_0085_),
    .S(_0918_),
    .Y(_0010_[3])
  );
  \$_MUX_  _1885_ (
    .A(_0089_),
    .B(inst_dext[4]),
    .S(_0913_),
    .Y(_0117_)
  );
  \$_MUX_  _1886_ (
    .A(_0117_),
    .B(_0089_),
    .S(_0918_),
    .Y(_0010_[4])
  );
  \$_MUX_  _1887_ (
    .A(_0092_),
    .B(inst_dext[5]),
    .S(_0913_),
    .Y(_0118_)
  );
  \$_MUX_  _1888_ (
    .A(_0118_),
    .B(_0092_),
    .S(_0918_),
    .Y(_0010_[5])
  );
  \$_MUX_  _1889_ (
    .A(_0095_),
    .B(inst_dext[6]),
    .S(_0913_),
    .Y(_0119_)
  );
  \$_MUX_  _1890_ (
    .A(_0119_),
    .B(_0095_),
    .S(_0918_),
    .Y(_0010_[6])
  );
  \$_MUX_  _1891_ (
    .A(_0098_),
    .B(inst_dext[7]),
    .S(_0913_),
    .Y(_0120_)
  );
  \$_MUX_  _1892_ (
    .A(_0120_),
    .B(_0098_),
    .S(_0918_),
    .Y(_0010_[7])
  );
  \$_MUX_  _1893_ (
    .A(_0101_),
    .B(inst_dext[8]),
    .S(_0913_),
    .Y(_0121_)
  );
  \$_MUX_  _1894_ (
    .A(_0121_),
    .B(_0101_),
    .S(_0918_),
    .Y(_0010_[8])
  );
  \$_MUX_  _1895_ (
    .A(_0104_),
    .B(inst_dext[9]),
    .S(_0913_),
    .Y(_0122_)
  );
  \$_MUX_  _1896_ (
    .A(_0122_),
    .B(_0104_),
    .S(_0918_),
    .Y(_0010_[9])
  );
  \$_MUX_  _1897_ (
    .A(inst_type[0]),
    .B(_0660_),
    .S(_1081_),
    .Y(_0018_[0])
  );
  \$_MUX_  _1898_ (
    .A(inst_type[1]),
    .B(_1104_),
    .S(_1081_),
    .Y(_0018_[1])
  );
  \$_INV_  _1899_ (
    .A(_0663_),
    .Y(_0123_)
  );
  \$_MUX_  _1900_ (
    .A(inst_type[2]),
    .B(_0123_),
    .S(_1081_),
    .Y(_0018_[2])
  );
  \$_AND_  _1901_ (
    .A(_0853_),
    .B(_0672_),
    .Y(_0124_)
  );
  \$_AND_  _1902_ (
    .A(_0124_),
    .B(_0660_),
    .Y(_0125_)
  );
  \$_MUX_  _1903_ (
    .A(_0125_),
    .B(inst_so[0]),
    .S(_1082_),
    .Y(_0015_[0])
  );
  \$_AND_  _1904_ (
    .A(_0854_),
    .B(_0672_),
    .Y(_0126_)
  );
  \$_AND_  _1905_ (
    .A(_0126_),
    .B(_0660_),
    .Y(_0127_)
  );
  \$_MUX_  _1906_ (
    .A(_0127_),
    .B(inst_so[1]),
    .S(_1082_),
    .Y(_0015_[1])
  );
  \$_AND_  _1907_ (
    .A(_0855_),
    .B(_0672_),
    .Y(_0128_)
  );
  \$_AND_  _1908_ (
    .A(_0128_),
    .B(_0660_),
    .Y(_0129_)
  );
  \$_MUX_  _1909_ (
    .A(_0129_),
    .B(inst_so[2]),
    .S(_1082_),
    .Y(_0015_[2])
  );
  \$_AND_  _1910_ (
    .A(_0857_),
    .B(_0672_),
    .Y(_0130_)
  );
  \$_AND_  _1911_ (
    .A(_0130_),
    .B(_0660_),
    .Y(_0131_)
  );
  \$_MUX_  _1912_ (
    .A(_0131_),
    .B(inst_so[3]),
    .S(_1082_),
    .Y(_0015_[3])
  );
  \$_MUX_  _1913_ (
    .A(_0970_),
    .B(inst_so[4]),
    .S(_1082_),
    .Y(_0015_[4])
  );
  \$_MUX_  _1914_ (
    .A(_0973_),
    .B(inst_so[5]),
    .S(_1082_),
    .Y(_0015_[5])
  );
  \$_MUX_  _1915_ (
    .A(_0866_),
    .B(inst_so[6]),
    .S(_1082_),
    .Y(_0015_[6])
  );
  \$_MUX_  _1916_ (
    .A(_0862_),
    .B(inst_so[7]),
    .S(_1082_),
    .Y(_0015_[7])
  );
  \$_MUX_  _1917_ (
    .A(inst_jmp_bin[0]),
    .B(mdb_in[10]),
    .S(_1081_),
    .Y(_0012_[0])
  );
  \$_MUX_  _1918_ (
    .A(inst_jmp_bin[1]),
    .B(mdb_in[11]),
    .S(_1081_),
    .Y(_0012_[1])
  );
  \$_MUX_  _1919_ (
    .A(inst_jmp_bin[2]),
    .B(mdb_in[12]),
    .S(_1081_),
    .Y(_0012_[2])
  );
  \$_AND_  _1920_ (
    .A(_0616_),
    .B(_0053_),
    .Y(_0132_)
  );
  \$_AND_  _1921_ (
    .A(_0132_),
    .B(mdb_in[14]),
    .Y(_0133_)
  );
  \$_AND_  _1922_ (
    .A(_0133_),
    .B(_0615_),
    .Y(_0134_)
  );
  \$_AND_  _1923_ (
    .A(_0134_),
    .B(_0123_),
    .Y(_0135_)
  );
  \$_MUX_  _1924_ (
    .A(_0135_),
    .B(inst_mov),
    .S(_1082_),
    .Y(_0013_)
  );
  \$_MUX_  _1925_ (
    .A(inst_dest_bin[0]),
    .B(mdb_in[0]),
    .S(_1081_),
    .Y(_0009_[0])
  );
  \$_MUX_  _1926_ (
    .A(inst_dest_bin[1]),
    .B(mdb_in[1]),
    .S(_1081_),
    .Y(_0009_[1])
  );
  \$_MUX_  _1927_ (
    .A(inst_dest_bin[2]),
    .B(mdb_in[2]),
    .S(_1081_),
    .Y(_0009_[2])
  );
  \$_MUX_  _1928_ (
    .A(inst_dest_bin[3]),
    .B(mdb_in[3]),
    .S(_1081_),
    .Y(_0009_[3])
  );
  \$_MUX_  _1929_ (
    .A(inst_src_bin[0]),
    .B(mdb_in[8]),
    .S(_1081_),
    .Y(_0016_[0])
  );
  \$_MUX_  _1930_ (
    .A(inst_src_bin[1]),
    .B(mdb_in[9]),
    .S(_1081_),
    .Y(_0016_[1])
  );
  \$_MUX_  _1931_ (
    .A(inst_src_bin[2]),
    .B(mdb_in[10]),
    .S(_1081_),
    .Y(_0016_[2])
  );
  \$_MUX_  _1932_ (
    .A(inst_src_bin[3]),
    .B(mdb_in[11]),
    .S(_1081_),
    .Y(_0016_[3])
  );
  \$_AND_  _1933_ (
    .A(_1090_),
    .B(_0640_),
    .Y(_0136_)
  );
  \$_OR_  _1934_ (
    .A(_0136_),
    .B(_1104_),
    .Y(_0137_)
  );
  \$_MUX_  _1935_ (
    .A(_0137_),
    .B(inst_as[0]),
    .S(_1082_),
    .Y(_0007_[0])
  );
  \$_AND_  _1936_ (
    .A(_0874_),
    .B(_0648_),
    .Y(_0138_)
  );
  \$_MUX_  _1937_ (
    .A(_0138_),
    .B(inst_as[1]),
    .S(_1082_),
    .Y(_0007_[1])
  );
  \$_MUX_  _1938_ (
    .A(_0873_),
    .B(inst_as[2]),
    .S(_1082_),
    .Y(_0007_[2])
  );
  \$_MUX_  _1939_ (
    .A(_0875_),
    .B(inst_as[3]),
    .S(_1082_),
    .Y(_0007_[3])
  );
  \$_AND_  _1940_ (
    .A(_0654_),
    .B(_0648_),
    .Y(_0139_)
  );
  \$_MUX_  _1941_ (
    .A(_0139_),
    .B(inst_as[4]),
    .S(_1082_),
    .Y(_0007_[4])
  );
  \$_MUX_  _1942_ (
    .A(_0658_),
    .B(inst_as[5]),
    .S(_1082_),
    .Y(_0007_[5])
  );
  \$_MUX_  _1943_ (
    .A(_0649_),
    .B(inst_as[6]),
    .S(_1082_),
    .Y(_0007_[6])
  );
  \$_INV_  _1944_ (
    .A(_1100_),
    .Y(_0140_)
  );
  \$_MUX_  _1945_ (
    .A(_0140_),
    .B(inst_as[7]),
    .S(_1082_),
    .Y(_0007_[7])
  );
  \$_AND_  _1946_ (
    .A(_0123_),
    .B(_0661_),
    .Y(_0141_)
  );
  \$_MUX_  _1947_ (
    .A(_0141_),
    .B(inst_ad[0]),
    .S(_1082_),
    .Y(_0005_[0])
  );
  \$_INV_  _1948_ (
    .A(_0967_),
    .Y(_0142_)
  );
  \$_MUX_  _1949_ (
    .A(_0142_),
    .B(inst_ad[1]),
    .S(_1082_),
    .Y(_0005_[1])
  );
  \$_AND_  _1950_ (
    .A(_1082_),
    .B(inst_ad[2]),
    .Y(_0005_[2])
  );
  \$_AND_  _1951_ (
    .A(_1082_),
    .B(inst_ad[3]),
    .Y(_0005_[3])
  );
  \$_INV_  _1952_ (
    .A(_0965_),
    .Y(_0143_)
  );
  \$_AND_  _1953_ (
    .A(_0143_),
    .B(_0668_),
    .Y(_0144_)
  );
  \$_AND_  _1954_ (
    .A(_0144_),
    .B(_0123_),
    .Y(_0145_)
  );
  \$_MUX_  _1955_ (
    .A(_0145_),
    .B(inst_ad[4]),
    .S(_1082_),
    .Y(_0005_[4])
  );
  \$_AND_  _1956_ (
    .A(_1082_),
    .B(inst_ad[5]),
    .Y(_0005_[5])
  );
  \$_AND_  _1957_ (
    .A(_0666_),
    .B(mdb_in[7]),
    .Y(_0146_)
  );
  \$_AND_  _1958_ (
    .A(_0146_),
    .B(_0123_),
    .Y(_0147_)
  );
  \$_MUX_  _1959_ (
    .A(_0147_),
    .B(inst_ad[6]),
    .S(_1082_),
    .Y(_0005_[6])
  );
  \$_AND_  _1960_ (
    .A(_1082_),
    .B(inst_ad[7]),
    .Y(_0005_[7])
  );
  \$_AND_  _1961_ (
    .A(_0611_),
    .B(mdb_in[6]),
    .Y(_0148_)
  );
  \$_AND_  _1962_ (
    .A(_0148_),
    .B(_0672_),
    .Y(_0149_)
  );
  \$_AND_  _1963_ (
    .A(_0149_),
    .B(_0644_),
    .Y(_0150_)
  );
  \$_MUX_  _1964_ (
    .A(_0150_),
    .B(inst_bw),
    .S(_1082_),
    .Y(_0008_)
  );
  \$_XOR_  _1965_ (
    .A(_0670_),
    .B(_0659_),
    .Y(_0151_)
  );
  \$_MUX_  _1966_ (
    .A(_0151_),
    .B(inst_sz[0]),
    .S(_1082_),
    .Y(_0017_[0])
  );
  \$_AND_  _1967_ (
    .A(_0670_),
    .B(_0659_),
    .Y(_0152_)
  );
  \$_MUX_  _1968_ (
    .A(_0152_),
    .B(inst_sz[1]),
    .S(_1082_),
    .Y(_0017_[1])
  );
  \$_AND_  _1969_ (
    .A(_0141_),
    .B(_0668_),
    .Y(_0153_)
  );
  \$_OR_  _1970_ (
    .A(_0866_),
    .B(_1104_),
    .Y(_0154_)
  );
  \$_OR_  _1971_ (
    .A(_0154_),
    .B(_0153_),
    .Y(_0155_)
  );
  \$_AND_  _1972_ (
    .A(_0155_),
    .B(_1081_),
    .Y(_0156_)
  );
  \$_AND_  _1973_ (
    .A(_0827_),
    .B(exec_jmp),
    .Y(_0157_)
  );
  \$_OR_  _1974_ (
    .A(_0157_),
    .B(_0156_),
    .Y(_0003_)
  );
  \$_AND_  _1975_ (
    .A(_0812_),
    .B(e_state[3]),
    .Y(_0158_)
  );
  \$_AND_  _1976_ (
    .A(_0821_),
    .B(exec_dst_wr),
    .Y(_0159_)
  );
  \$_OR_  _1977_ (
    .A(_0159_),
    .B(_0158_),
    .Y(_0002_)
  );
  \$_AND_  _1978_ (
    .A(_0822_),
    .B(inst_type[0]),
    .Y(_0160_)
  );
  \$_AND_  _1979_ (
    .A(_0828_),
    .B(exec_src_wr),
    .Y(_0161_)
  );
  \$_AND_  _1980_ (
    .A(_0161_),
    .B(_0821_),
    .Y(_0162_)
  );
  \$_OR_  _1981_ (
    .A(_0162_),
    .B(_0160_),
    .Y(_0004_)
  );
  \$_INV_  _1982_ (
    .A(_0158_),
    .Y(_0163_)
  );
  \$_AND_  _1983_ (
    .A(_0922_),
    .B(_0163_),
    .Y(_0001_)
  );
  \$_AND_  _1984_ (
    .A(_0132_),
    .B(_0617_),
    .Y(_0164_)
  );
  \$_AND_  _1985_ (
    .A(_0164_),
    .B(mdb_in[15]),
    .Y(_0165_)
  );
  \$_AND_  _1986_ (
    .A(_0165_),
    .B(_0123_),
    .Y(_0166_)
  );
  \$_AND_  _1987_ (
    .A(mdb_in[13]),
    .B(mdb_in[12]),
    .Y(_0167_)
  );
  \$_AND_  _1988_ (
    .A(_0615_),
    .B(mdb_in[14]),
    .Y(_0168_)
  );
  \$_AND_  _1989_ (
    .A(_0168_),
    .B(_0167_),
    .Y(_0169_)
  );
  \$_AND_  _1990_ (
    .A(_0169_),
    .B(_0123_),
    .Y(_0170_)
  );
  \$_OR_  _1991_ (
    .A(_0170_),
    .B(_0166_),
    .Y(_0171_)
  );
  \$_AND_  _1992_ (
    .A(_0616_),
    .B(mdb_in[12]),
    .Y(_0172_)
  );
  \$_AND_  _1993_ (
    .A(_0172_),
    .B(_0617_),
    .Y(_0173_)
  );
  \$_AND_  _1994_ (
    .A(_0173_),
    .B(mdb_in[15]),
    .Y(_0174_)
  );
  \$_AND_  _1995_ (
    .A(_0174_),
    .B(_0123_),
    .Y(_0175_)
  );
  \$_AND_  _1996_ (
    .A(_0133_),
    .B(mdb_in[15]),
    .Y(_0176_)
  );
  \$_AND_  _1997_ (
    .A(_0176_),
    .B(_0123_),
    .Y(_0177_)
  );
  \$_OR_  _1998_ (
    .A(_0177_),
    .B(_0175_),
    .Y(_0178_)
  );
  \$_OR_  _1999_ (
    .A(_0178_),
    .B(_0171_),
    .Y(_0179_)
  );
  \$_MUX_  _2000_ (
    .A(_0179_),
    .B(inst_alu[0]),
    .S(_1082_),
    .Y(_0006_[0])
  );
  \$_OR_  _2001_ (
    .A(_0129_),
    .B(_0125_),
    .Y(_0180_)
  );
  \$_MUX_  _2002_ (
    .A(_0180_),
    .B(inst_alu[10]),
    .S(_1082_),
    .Y(_0006_[10])
  );
  \$_AND_  _2003_ (
    .A(_0167_),
    .B(_0617_),
    .Y(_0181_)
  );
  \$_AND_  _2004_ (
    .A(_0181_),
    .B(mdb_in[15]),
    .Y(_0182_)
  );
  \$_AND_  _2005_ (
    .A(_0182_),
    .B(_0123_),
    .Y(_0183_)
  );
  \$_OR_  _2006_ (
    .A(_0183_),
    .B(_0175_),
    .Y(_0184_)
  );
  \$_MUX_  _2007_ (
    .A(_0184_),
    .B(inst_alu[11]),
    .S(_1082_),
    .Y(_0006_[11])
  );
  \$_OR_  _2008_ (
    .A(_0175_),
    .B(_0166_),
    .Y(_0185_)
  );
  \$_MUX_  _2009_ (
    .A(_0185_),
    .B(inst_alu[1]),
    .S(_1082_),
    .Y(_0006_[1])
  );
  \$_AND_  _2010_ (
    .A(mdb_in[13]),
    .B(_0053_),
    .Y(_0186_)
  );
  \$_AND_  _2011_ (
    .A(_0186_),
    .B(_0617_),
    .Y(_0187_)
  );
  \$_AND_  _2012_ (
    .A(_0187_),
    .B(mdb_in[15]),
    .Y(_0188_)
  );
  \$_AND_  _2013_ (
    .A(_0188_),
    .B(_0123_),
    .Y(_0189_)
  );
  \$_AND_  _2014_ (
    .A(_0186_),
    .B(mdb_in[14]),
    .Y(_0190_)
  );
  \$_AND_  _2015_ (
    .A(_0190_),
    .B(_0615_),
    .Y(_0191_)
  );
  \$_AND_  _2016_ (
    .A(_0191_),
    .B(_0123_),
    .Y(_0192_)
  );
  \$_OR_  _2017_ (
    .A(_0192_),
    .B(_0170_),
    .Y(_0193_)
  );
  \$_OR_  _2018_ (
    .A(_0193_),
    .B(_0189_),
    .Y(_0194_)
  );
  \$_MUX_  _2019_ (
    .A(_0194_),
    .B(inst_alu[2]),
    .S(_1082_),
    .Y(_0006_[2])
  );
  \$_AND_  _2020_ (
    .A(_0172_),
    .B(mdb_in[14]),
    .Y(_0195_)
  );
  \$_AND_  _2021_ (
    .A(_0195_),
    .B(_0615_),
    .Y(_0196_)
  );
  \$_AND_  _2022_ (
    .A(_0196_),
    .B(_0123_),
    .Y(_0197_)
  );
  \$_OR_  _2023_ (
    .A(_0192_),
    .B(_0175_),
    .Y(_0198_)
  );
  \$_OR_  _2024_ (
    .A(_0198_),
    .B(_0197_),
    .Y(_0199_)
  );
  \$_OR_  _2025_ (
    .A(_0199_),
    .B(_0171_),
    .Y(_0200_)
  );
  \$_OR_  _2026_ (
    .A(_0200_),
    .B(_0154_),
    .Y(_0201_)
  );
  \$_MUX_  _2027_ (
    .A(_0201_),
    .B(inst_alu[3]),
    .S(_1082_),
    .Y(_0006_[3])
  );
  \$_INV_  _2028_ (
    .A(_0176_),
    .Y(_0202_)
  );
  \$_INV_  _2029_ (
    .A(_0182_),
    .Y(_0203_)
  );
  \$_AND_  _2030_ (
    .A(_0203_),
    .B(_0202_),
    .Y(_0204_)
  );
  \$_INV_  _2031_ (
    .A(_0187_),
    .Y(_0205_)
  );
  \$_INV_  _2032_ (
    .A(_0190_),
    .Y(_0206_)
  );
  \$_MUX_  _2033_ (
    .A(_0206_),
    .B(_0205_),
    .S(mdb_in[15]),
    .Y(_0207_)
  );
  \$_AND_  _2034_ (
    .A(_0207_),
    .B(_0204_),
    .Y(_0208_)
  );
  \$_INV_  _2035_ (
    .A(_0134_),
    .Y(_0209_)
  );
  \$_INV_  _2036_ (
    .A(_0169_),
    .Y(_0210_)
  );
  \$_AND_  _2037_ (
    .A(_0210_),
    .B(_0209_),
    .Y(_0211_)
  );
  \$_INV_  _2038_ (
    .A(_0165_),
    .Y(_0212_)
  );
  \$_INV_  _2039_ (
    .A(_0174_),
    .Y(_0213_)
  );
  \$_AND_  _2040_ (
    .A(_0213_),
    .B(_0212_),
    .Y(_0214_)
  );
  \$_AND_  _2041_ (
    .A(_0214_),
    .B(_0211_),
    .Y(_0215_)
  );
  \$_AND_  _2042_ (
    .A(_0215_),
    .B(_0208_),
    .Y(_0216_)
  );
  \$_AND_  _2043_ (
    .A(_0190_),
    .B(mdb_in[15]),
    .Y(_0217_)
  );
  \$_INV_  _2044_ (
    .A(_0217_),
    .Y(_0218_)
  );
  \$_INV_  _2045_ (
    .A(_0181_),
    .Y(_0219_)
  );
  \$_INV_  _2046_ (
    .A(_0195_),
    .Y(_0220_)
  );
  \$_MUX_  _2047_ (
    .A(_0220_),
    .B(_0219_),
    .S(_0615_),
    .Y(_0221_)
  );
  \$_AND_  _2048_ (
    .A(_0221_),
    .B(_0218_),
    .Y(_0222_)
  );
  \$_INV_  _2049_ (
    .A(_0196_),
    .Y(_0223_)
  );
  \$_INV_  _2050_ (
    .A(_0164_),
    .Y(_0224_)
  );
  \$_OR_  _2051_ (
    .A(_0224_),
    .B(mdb_in[15]),
    .Y(_0225_)
  );
  \$_AND_  _2052_ (
    .A(_0225_),
    .B(_0223_),
    .Y(_0226_)
  );
  \$_INV_  _2053_ (
    .A(_0173_),
    .Y(_0227_)
  );
  \$_OR_  _2054_ (
    .A(_0227_),
    .B(mdb_in[15]),
    .Y(_0228_)
  );
  \$_OR_  _2055_ (
    .A(_0205_),
    .B(mdb_in[15]),
    .Y(_0229_)
  );
  \$_AND_  _2056_ (
    .A(_0229_),
    .B(_0228_),
    .Y(_0230_)
  );
  \$_AND_  _2057_ (
    .A(_0230_),
    .B(_0226_),
    .Y(_0231_)
  );
  \$_AND_  _2058_ (
    .A(_0231_),
    .B(_0222_),
    .Y(_0232_)
  );
  \$_AND_  _2059_ (
    .A(_0232_),
    .B(_0216_),
    .Y(_0233_)
  );
  \$_AND_  _2060_ (
    .A(_0233_),
    .B(_0123_),
    .Y(_0234_)
  );
  \$_OR_  _2061_ (
    .A(_0183_),
    .B(_0177_),
    .Y(_0235_)
  );
  \$_OR_  _2062_ (
    .A(_0235_),
    .B(_0234_),
    .Y(_0236_)
  );
  \$_MUX_  _2063_ (
    .A(_0236_),
    .B(inst_alu[4]),
    .S(_1082_),
    .Y(_0006_[4])
  );
  \$_AND_  _2064_ (
    .A(_0195_),
    .B(mdb_in[15]),
    .Y(_0237_)
  );
  \$_AND_  _2065_ (
    .A(_0237_),
    .B(_0123_),
    .Y(_0238_)
  );
  \$_MUX_  _2066_ (
    .A(_0238_),
    .B(inst_alu[5]),
    .S(_1082_),
    .Y(_0006_[5])
  );
  \$_AND_  _2067_ (
    .A(_0217_),
    .B(_0123_),
    .Y(_0239_)
  );
  \$_MUX_  _2068_ (
    .A(_0239_),
    .B(inst_alu[6]),
    .S(_1082_),
    .Y(_0006_[6])
  );
  \$_MUX_  _2069_ (
    .A(_0189_),
    .B(inst_alu[7]),
    .S(_1082_),
    .Y(_0006_[7])
  );
  \$_OR_  _2070_ (
    .A(_0183_),
    .B(_0131_),
    .Y(_0240_)
  );
  \$_OR_  _2071_ (
    .A(_0240_),
    .B(_0234_),
    .Y(_0241_)
  );
  \$_MUX_  _2072_ (
    .A(_0241_),
    .B(inst_alu[8]),
    .S(_1082_),
    .Y(_0006_[8])
  );
  \$_OR_  _2073_ (
    .A(_0234_),
    .B(_0189_),
    .Y(_0242_)
  );
  \$_OR_  _2074_ (
    .A(_0242_),
    .B(_0239_),
    .Y(_0243_)
  );
  \$_OR_  _2075_ (
    .A(_0240_),
    .B(_0180_),
    .Y(_0244_)
  );
  \$_OR_  _2076_ (
    .A(_0244_),
    .B(_0243_),
    .Y(_0245_)
  );
  \$_OR_  _2077_ (
    .A(_0245_),
    .B(_0200_),
    .Y(_0246_)
  );
  \$_MUX_  _2078_ (
    .A(_0246_),
    .B(inst_alu[9]),
    .S(_1082_),
    .Y(_0006_[9])
  );
  \$_INV_  _2079_ (
    .A(_0893_),
    .Y(e_state_nxt[2])
  );
  \$_INV_  _2080_ (
    .A(_0963_),
    .Y(e_state_nxt[3])
  );
  \$_AND_  _2081_ (
    .A(pc_sw[0]),
    .B(pc_sw_wr),
    .Y(_0247_)
  );
  \$_MUX_  _2082_ (
    .A(pc[0]),
    .B(mdb_in[0]),
    .S(i_state[2]),
    .Y(_0248_)
  );
  \$_AND_  _2083_ (
    .A(_0248_),
    .B(_0678_),
    .Y(_0249_)
  );
  \$_AND_  _2084_ (
    .A(_0249_),
    .B(_0729_),
    .Y(_0250_)
  );
  \$_OR_  _2085_ (
    .A(_0250_),
    .B(_0247_),
    .Y(mab[0])
  );
  \$_AND_  _2086_ (
    .A(_1007_),
    .B(pc[1]),
    .Y(_0251_)
  );
  \$_AND_  _2087_ (
    .A(_0251_),
    .B(pc[2]),
    .Y(_0252_)
  );
  \$_AND_  _2088_ (
    .A(_0252_),
    .B(pc[3]),
    .Y(_0253_)
  );
  \$_AND_  _2089_ (
    .A(_0253_),
    .B(pc[4]),
    .Y(_0254_)
  );
  \$_AND_  _2090_ (
    .A(_0254_),
    .B(pc[5]),
    .Y(_0255_)
  );
  \$_AND_  _2091_ (
    .A(_0255_),
    .B(pc[6]),
    .Y(_0256_)
  );
  \$_AND_  _2092_ (
    .A(_0256_),
    .B(pc[7]),
    .Y(_0257_)
  );
  \$_AND_  _2093_ (
    .A(_0257_),
    .B(pc[8]),
    .Y(_0258_)
  );
  \$_AND_  _2094_ (
    .A(_0258_),
    .B(pc[9]),
    .Y(_0259_)
  );
  \$_XOR_  _2095_ (
    .A(_0259_),
    .B(pc[10]),
    .Y(_0260_)
  );
  \$_MUX_  _2096_ (
    .A(_0260_),
    .B(mdb_in[10]),
    .S(i_state[2]),
    .Y(_0261_)
  );
  \$_OR_  _2097_ (
    .A(_0261_),
    .B(_1142_[15]),
    .Y(_0262_)
  );
  \$_MUX_  _2098_ (
    .A(_0262_),
    .B(pc_sw[10]),
    .S(pc_sw_wr),
    .Y(mab[10])
  );
  \$_AND_  _2099_ (
    .A(_0259_),
    .B(pc[10]),
    .Y(_0263_)
  );
  \$_XOR_  _2100_ (
    .A(_0263_),
    .B(pc[11]),
    .Y(_0264_)
  );
  \$_MUX_  _2101_ (
    .A(_0264_),
    .B(mdb_in[11]),
    .S(i_state[2]),
    .Y(_0265_)
  );
  \$_OR_  _2102_ (
    .A(_0265_),
    .B(_1142_[15]),
    .Y(_0266_)
  );
  \$_MUX_  _2103_ (
    .A(_0266_),
    .B(pc_sw[11]),
    .S(pc_sw_wr),
    .Y(mab[11])
  );
  \$_AND_  _2104_ (
    .A(_0263_),
    .B(pc[11]),
    .Y(_0267_)
  );
  \$_XOR_  _2105_ (
    .A(_0267_),
    .B(pc[12]),
    .Y(_0268_)
  );
  \$_MUX_  _2106_ (
    .A(_0268_),
    .B(mdb_in[12]),
    .S(i_state[2]),
    .Y(_0269_)
  );
  \$_OR_  _2107_ (
    .A(_0269_),
    .B(_1142_[15]),
    .Y(_0270_)
  );
  \$_MUX_  _2108_ (
    .A(_0270_),
    .B(pc_sw[12]),
    .S(pc_sw_wr),
    .Y(mab[12])
  );
  \$_AND_  _2109_ (
    .A(_0267_),
    .B(pc[12]),
    .Y(_0271_)
  );
  \$_XOR_  _2110_ (
    .A(_0271_),
    .B(pc[13]),
    .Y(_0272_)
  );
  \$_MUX_  _2111_ (
    .A(_0272_),
    .B(mdb_in[13]),
    .S(i_state[2]),
    .Y(_0273_)
  );
  \$_OR_  _2112_ (
    .A(_0273_),
    .B(_1142_[15]),
    .Y(_0274_)
  );
  \$_MUX_  _2113_ (
    .A(_0274_),
    .B(pc_sw[13]),
    .S(pc_sw_wr),
    .Y(mab[13])
  );
  \$_AND_  _2114_ (
    .A(_0271_),
    .B(pc[13]),
    .Y(_0275_)
  );
  \$_XOR_  _2115_ (
    .A(_0275_),
    .B(pc[14]),
    .Y(_0276_)
  );
  \$_MUX_  _2116_ (
    .A(_0276_),
    .B(mdb_in[14]),
    .S(i_state[2]),
    .Y(_0277_)
  );
  \$_OR_  _2117_ (
    .A(_0277_),
    .B(_1142_[15]),
    .Y(_0278_)
  );
  \$_MUX_  _2118_ (
    .A(_0278_),
    .B(pc_sw[14]),
    .S(pc_sw_wr),
    .Y(mab[14])
  );
  \$_AND_  _2119_ (
    .A(_0275_),
    .B(pc[14]),
    .Y(_0279_)
  );
  \$_XOR_  _2120_ (
    .A(_0279_),
    .B(pc[15]),
    .Y(_0280_)
  );
  \$_MUX_  _2121_ (
    .A(_0280_),
    .B(mdb_in[15]),
    .S(i_state[2]),
    .Y(_0281_)
  );
  \$_OR_  _2122_ (
    .A(_0281_),
    .B(_1142_[15]),
    .Y(_0282_)
  );
  \$_MUX_  _2123_ (
    .A(_0282_),
    .B(pc_sw[15]),
    .S(pc_sw_wr),
    .Y(mab[15])
  );
  \$_XOR_  _2124_ (
    .A(_1007_),
    .B(pc[1]),
    .Y(_0283_)
  );
  \$_MUX_  _2125_ (
    .A(_0283_),
    .B(mdb_in[1]),
    .S(i_state[2]),
    .Y(_0284_)
  );
  \$_MUX_  _2126_ (
    .A(_0284_),
    .B(irq_addr[1]),
    .S(_1142_[15]),
    .Y(_0285_)
  );
  \$_MUX_  _2127_ (
    .A(_0285_),
    .B(pc_sw[1]),
    .S(pc_sw_wr),
    .Y(mab[1])
  );
  \$_XOR_  _2128_ (
    .A(_0251_),
    .B(pc[2]),
    .Y(_0286_)
  );
  \$_MUX_  _2129_ (
    .A(_0286_),
    .B(mdb_in[2]),
    .S(i_state[2]),
    .Y(_0287_)
  );
  \$_MUX_  _2130_ (
    .A(_0287_),
    .B(irq_addr[2]),
    .S(_1142_[15]),
    .Y(_0288_)
  );
  \$_MUX_  _2131_ (
    .A(_0288_),
    .B(pc_sw[2]),
    .S(pc_sw_wr),
    .Y(mab[2])
  );
  \$_XOR_  _2132_ (
    .A(_0252_),
    .B(pc[3]),
    .Y(_0289_)
  );
  \$_MUX_  _2133_ (
    .A(_0289_),
    .B(mdb_in[3]),
    .S(i_state[2]),
    .Y(_0290_)
  );
  \$_MUX_  _2134_ (
    .A(_0290_),
    .B(irq_addr[3]),
    .S(_1142_[15]),
    .Y(_0291_)
  );
  \$_MUX_  _2135_ (
    .A(_0291_),
    .B(pc_sw[3]),
    .S(pc_sw_wr),
    .Y(mab[3])
  );
  \$_XOR_  _2136_ (
    .A(_0253_),
    .B(pc[4]),
    .Y(_0292_)
  );
  \$_MUX_  _2137_ (
    .A(_0292_),
    .B(mdb_in[4]),
    .S(i_state[2]),
    .Y(_0293_)
  );
  \$_MUX_  _2138_ (
    .A(_0293_),
    .B(irq_addr[4]),
    .S(_1142_[15]),
    .Y(_0294_)
  );
  \$_MUX_  _2139_ (
    .A(_0294_),
    .B(pc_sw[4]),
    .S(pc_sw_wr),
    .Y(mab[4])
  );
  \$_XOR_  _2140_ (
    .A(_0254_),
    .B(pc[5]),
    .Y(_0295_)
  );
  \$_MUX_  _2141_ (
    .A(_0295_),
    .B(mdb_in[5]),
    .S(i_state[2]),
    .Y(_0296_)
  );
  \$_OR_  _2142_ (
    .A(_0296_),
    .B(_1142_[15]),
    .Y(_0297_)
  );
  \$_MUX_  _2143_ (
    .A(_0297_),
    .B(pc_sw[5]),
    .S(pc_sw_wr),
    .Y(mab[5])
  );
  \$_XOR_  _2144_ (
    .A(_0255_),
    .B(pc[6]),
    .Y(_0298_)
  );
  \$_MUX_  _2145_ (
    .A(_0298_),
    .B(mdb_in[6]),
    .S(i_state[2]),
    .Y(_0299_)
  );
  \$_OR_  _2146_ (
    .A(_0299_),
    .B(_1142_[15]),
    .Y(_0300_)
  );
  \$_MUX_  _2147_ (
    .A(_0300_),
    .B(pc_sw[6]),
    .S(pc_sw_wr),
    .Y(mab[6])
  );
  \$_XOR_  _2148_ (
    .A(_0256_),
    .B(pc[7]),
    .Y(_0301_)
  );
  \$_MUX_  _2149_ (
    .A(_0301_),
    .B(mdb_in[7]),
    .S(i_state[2]),
    .Y(_0302_)
  );
  \$_OR_  _2150_ (
    .A(_0302_),
    .B(_1142_[15]),
    .Y(_0303_)
  );
  \$_MUX_  _2151_ (
    .A(_0303_),
    .B(pc_sw[7]),
    .S(pc_sw_wr),
    .Y(mab[7])
  );
  \$_XOR_  _2152_ (
    .A(_0257_),
    .B(pc[8]),
    .Y(_0304_)
  );
  \$_MUX_  _2153_ (
    .A(_0304_),
    .B(mdb_in[8]),
    .S(i_state[2]),
    .Y(_0305_)
  );
  \$_OR_  _2154_ (
    .A(_0305_),
    .B(_1142_[15]),
    .Y(_0306_)
  );
  \$_MUX_  _2155_ (
    .A(_0306_),
    .B(pc_sw[8]),
    .S(pc_sw_wr),
    .Y(mab[8])
  );
  \$_XOR_  _2156_ (
    .A(_0258_),
    .B(pc[9]),
    .Y(_0307_)
  );
  \$_MUX_  _2157_ (
    .A(_0307_),
    .B(mdb_in[9]),
    .S(i_state[2]),
    .Y(_0308_)
  );
  \$_OR_  _2158_ (
    .A(_0308_),
    .B(_1142_[15]),
    .Y(_0309_)
  );
  \$_MUX_  _2159_ (
    .A(_0309_),
    .B(pc_sw[9]),
    .S(pc_sw_wr),
    .Y(mab[9])
  );
  \$_INV_  _2160_ (
    .A(dbg_reg_sel[3]),
    .Y(_0310_)
  );
  \$_INV_  _2161_ (
    .A(dbg_reg_sel[2]),
    .Y(_0311_)
  );
  \$_INV_  _2162_ (
    .A(dbg_reg_sel[0]),
    .Y(_0312_)
  );
  \$_INV_  _2163_ (
    .A(dbg_reg_sel[1]),
    .Y(_0313_)
  );
  \$_AND_  _2164_ (
    .A(_0313_),
    .B(_0312_),
    .Y(_0314_)
  );
  \$_AND_  _2165_ (
    .A(_0314_),
    .B(_0311_),
    .Y(_0315_)
  );
  \$_AND_  _2166_ (
    .A(_0315_),
    .B(_0310_),
    .Y(_0316_)
  );
  \$_INV_  _2167_ (
    .A(inst_dest_bin[3]),
    .Y(_0317_)
  );
  \$_INV_  _2168_ (
    .A(inst_dest_bin[2]),
    .Y(_0318_)
  );
  \$_INV_  _2169_ (
    .A(inst_dest_bin[0]),
    .Y(_0319_)
  );
  \$_INV_  _2170_ (
    .A(inst_dest_bin[1]),
    .Y(_0320_)
  );
  \$_AND_  _2171_ (
    .A(_0320_),
    .B(_0319_),
    .Y(_0321_)
  );
  \$_AND_  _2172_ (
    .A(_0321_),
    .B(_0318_),
    .Y(_0322_)
  );
  \$_AND_  _2173_ (
    .A(_0322_),
    .B(_0317_),
    .Y(_0323_)
  );
  \$_INV_  _2174_ (
    .A(inst_type[1]),
    .Y(_0324_)
  );
  \$_INV_  _2175_ (
    .A(inst_so[7]),
    .Y(_0325_)
  );
  \$_AND_  _2176_ (
    .A(_0993_),
    .B(_0325_),
    .Y(_0326_)
  );
  \$_AND_  _2177_ (
    .A(_0326_),
    .B(_0324_),
    .Y(_0327_)
  );
  \$_AND_  _2178_ (
    .A(_0327_),
    .B(_0323_),
    .Y(_0328_)
  );
  \$_OR_  _2179_ (
    .A(_0328_),
    .B(inst_type[1]),
    .Y(_0329_)
  );
  \$_MUX_  _2180_ (
    .A(_0329_),
    .B(_0316_),
    .S(dbg_halt_st),
    .Y(inst_dest[0])
  );
  \$_AND_  _2181_ (
    .A(dbg_reg_sel[1]),
    .B(_0312_),
    .Y(_0330_)
  );
  \$_AND_  _2182_ (
    .A(_0330_),
    .B(_0311_),
    .Y(_0331_)
  );
  \$_AND_  _2183_ (
    .A(_0331_),
    .B(dbg_reg_sel[3]),
    .Y(_0332_)
  );
  \$_AND_  _2184_ (
    .A(_0332_),
    .B(dbg_halt_st),
    .Y(_0333_)
  );
  \$_AND_  _2185_ (
    .A(inst_dest_bin[1]),
    .B(_0319_),
    .Y(_0334_)
  );
  \$_AND_  _2186_ (
    .A(_0334_),
    .B(_0318_),
    .Y(_0335_)
  );
  \$_AND_  _2187_ (
    .A(_0335_),
    .B(inst_dest_bin[3]),
    .Y(_0336_)
  );
  \$_AND_  _2188_ (
    .A(_0324_),
    .B(_0609_),
    .Y(_0337_)
  );
  \$_AND_  _2189_ (
    .A(_0337_),
    .B(_0326_),
    .Y(_0338_)
  );
  \$_AND_  _2190_ (
    .A(_0338_),
    .B(_0336_),
    .Y(_0339_)
  );
  \$_OR_  _2191_ (
    .A(_0339_),
    .B(_0333_),
    .Y(inst_dest[10])
  );
  \$_AND_  _2192_ (
    .A(dbg_reg_sel[1]),
    .B(dbg_reg_sel[0]),
    .Y(_0340_)
  );
  \$_AND_  _2193_ (
    .A(_0340_),
    .B(_0311_),
    .Y(_0341_)
  );
  \$_AND_  _2194_ (
    .A(_0341_),
    .B(dbg_reg_sel[3]),
    .Y(_0342_)
  );
  \$_AND_  _2195_ (
    .A(_0342_),
    .B(dbg_halt_st),
    .Y(_0343_)
  );
  \$_AND_  _2196_ (
    .A(inst_dest_bin[1]),
    .B(inst_dest_bin[0]),
    .Y(_0344_)
  );
  \$_AND_  _2197_ (
    .A(_0344_),
    .B(_0318_),
    .Y(_0345_)
  );
  \$_AND_  _2198_ (
    .A(_0345_),
    .B(inst_dest_bin[3]),
    .Y(_0346_)
  );
  \$_AND_  _2199_ (
    .A(_0346_),
    .B(_0338_),
    .Y(_0347_)
  );
  \$_OR_  _2200_ (
    .A(_0347_),
    .B(_0343_),
    .Y(inst_dest[11])
  );
  \$_AND_  _2201_ (
    .A(_0314_),
    .B(dbg_reg_sel[2]),
    .Y(_0348_)
  );
  \$_AND_  _2202_ (
    .A(_0348_),
    .B(dbg_reg_sel[3]),
    .Y(_0349_)
  );
  \$_AND_  _2203_ (
    .A(_0349_),
    .B(dbg_halt_st),
    .Y(_0350_)
  );
  \$_AND_  _2204_ (
    .A(_0321_),
    .B(inst_dest_bin[2]),
    .Y(_0351_)
  );
  \$_AND_  _2205_ (
    .A(_0351_),
    .B(inst_dest_bin[3]),
    .Y(_0352_)
  );
  \$_AND_  _2206_ (
    .A(_0352_),
    .B(_0338_),
    .Y(_0353_)
  );
  \$_OR_  _2207_ (
    .A(_0353_),
    .B(_0350_),
    .Y(inst_dest[12])
  );
  \$_AND_  _2208_ (
    .A(_0313_),
    .B(dbg_reg_sel[0]),
    .Y(_0354_)
  );
  \$_AND_  _2209_ (
    .A(_0354_),
    .B(dbg_reg_sel[2]),
    .Y(_0355_)
  );
  \$_AND_  _2210_ (
    .A(_0355_),
    .B(dbg_reg_sel[3]),
    .Y(_0356_)
  );
  \$_AND_  _2211_ (
    .A(_0356_),
    .B(dbg_halt_st),
    .Y(_0357_)
  );
  \$_AND_  _2212_ (
    .A(_0320_),
    .B(inst_dest_bin[0]),
    .Y(_0358_)
  );
  \$_AND_  _2213_ (
    .A(_0358_),
    .B(inst_dest_bin[2]),
    .Y(_0359_)
  );
  \$_AND_  _2214_ (
    .A(_0359_),
    .B(inst_dest_bin[3]),
    .Y(_0360_)
  );
  \$_AND_  _2215_ (
    .A(_0360_),
    .B(_0338_),
    .Y(_0361_)
  );
  \$_OR_  _2216_ (
    .A(_0361_),
    .B(_0357_),
    .Y(inst_dest[13])
  );
  \$_AND_  _2217_ (
    .A(_0330_),
    .B(dbg_reg_sel[2]),
    .Y(_0362_)
  );
  \$_AND_  _2218_ (
    .A(_0362_),
    .B(dbg_reg_sel[3]),
    .Y(_0363_)
  );
  \$_AND_  _2219_ (
    .A(_0363_),
    .B(dbg_halt_st),
    .Y(_0364_)
  );
  \$_AND_  _2220_ (
    .A(_0334_),
    .B(inst_dest_bin[2]),
    .Y(_0365_)
  );
  \$_AND_  _2221_ (
    .A(_0365_),
    .B(inst_dest_bin[3]),
    .Y(_0366_)
  );
  \$_AND_  _2222_ (
    .A(_0366_),
    .B(_0338_),
    .Y(_0367_)
  );
  \$_OR_  _2223_ (
    .A(_0367_),
    .B(_0364_),
    .Y(inst_dest[14])
  );
  \$_INV_  _2224_ (
    .A(_0349_),
    .Y(_0368_)
  );
  \$_INV_  _2225_ (
    .A(_0356_),
    .Y(_0369_)
  );
  \$_AND_  _2226_ (
    .A(_0369_),
    .B(_0368_),
    .Y(_0370_)
  );
  \$_INV_  _2227_ (
    .A(_0362_),
    .Y(_0371_)
  );
  \$_AND_  _2228_ (
    .A(_0354_),
    .B(_0311_),
    .Y(_0372_)
  );
  \$_INV_  _2229_ (
    .A(_0372_),
    .Y(_0373_)
  );
  \$_MUX_  _2230_ (
    .A(_0373_),
    .B(_0371_),
    .S(dbg_reg_sel[3]),
    .Y(_0374_)
  );
  \$_AND_  _2231_ (
    .A(_0374_),
    .B(_0370_),
    .Y(_0375_)
  );
  \$_INV_  _2232_ (
    .A(_0316_),
    .Y(_0376_)
  );
  \$_AND_  _2233_ (
    .A(_0310_),
    .B(dbg_reg_sel[2]),
    .Y(_0377_)
  );
  \$_AND_  _2234_ (
    .A(_0377_),
    .B(_0340_),
    .Y(_0378_)
  );
  \$_INV_  _2235_ (
    .A(_0378_),
    .Y(_0379_)
  );
  \$_AND_  _2236_ (
    .A(_0379_),
    .B(dbg_halt_st),
    .Y(_0380_)
  );
  \$_AND_  _2237_ (
    .A(_0380_),
    .B(_0376_),
    .Y(_0381_)
  );
  \$_INV_  _2238_ (
    .A(_0332_),
    .Y(_0382_)
  );
  \$_INV_  _2239_ (
    .A(_0342_),
    .Y(_0383_)
  );
  \$_AND_  _2240_ (
    .A(_0383_),
    .B(_0382_),
    .Y(_0384_)
  );
  \$_AND_  _2241_ (
    .A(_0384_),
    .B(_0381_),
    .Y(_0385_)
  );
  \$_AND_  _2242_ (
    .A(_0385_),
    .B(_0375_),
    .Y(_0386_)
  );
  \$_AND_  _2243_ (
    .A(_0372_),
    .B(dbg_reg_sel[3]),
    .Y(_0387_)
  );
  \$_INV_  _2244_ (
    .A(_0387_),
    .Y(_0388_)
  );
  \$_INV_  _2245_ (
    .A(_0315_),
    .Y(_0389_)
  );
  \$_MUX_  _2246_ (
    .A(_0371_),
    .B(_0389_),
    .S(dbg_reg_sel[3]),
    .Y(_0390_)
  );
  \$_AND_  _2247_ (
    .A(_0390_),
    .B(_0388_),
    .Y(_0391_)
  );
  \$_AND_  _2248_ (
    .A(_0331_),
    .B(_0310_),
    .Y(_0392_)
  );
  \$_INV_  _2249_ (
    .A(_0392_),
    .Y(_0393_)
  );
  \$_AND_  _2250_ (
    .A(_0341_),
    .B(_0310_),
    .Y(_0394_)
  );
  \$_INV_  _2251_ (
    .A(_0394_),
    .Y(_0395_)
  );
  \$_AND_  _2252_ (
    .A(_0395_),
    .B(_0393_),
    .Y(_0396_)
  );
  \$_AND_  _2253_ (
    .A(_0348_),
    .B(_0310_),
    .Y(_0397_)
  );
  \$_INV_  _2254_ (
    .A(_0397_),
    .Y(_0398_)
  );
  \$_AND_  _2255_ (
    .A(_0355_),
    .B(_0310_),
    .Y(_0399_)
  );
  \$_INV_  _2256_ (
    .A(_0399_),
    .Y(_0400_)
  );
  \$_AND_  _2257_ (
    .A(_0400_),
    .B(_0398_),
    .Y(_0401_)
  );
  \$_AND_  _2258_ (
    .A(_0401_),
    .B(_0396_),
    .Y(_0402_)
  );
  \$_AND_  _2259_ (
    .A(_0402_),
    .B(_0391_),
    .Y(_0403_)
  );
  \$_AND_  _2260_ (
    .A(_0403_),
    .B(_0386_),
    .Y(_0404_)
  );
  \$_INV_  _2261_ (
    .A(_0352_),
    .Y(_0405_)
  );
  \$_INV_  _2262_ (
    .A(_0360_),
    .Y(_0406_)
  );
  \$_AND_  _2263_ (
    .A(_0406_),
    .B(_0405_),
    .Y(_0407_)
  );
  \$_INV_  _2264_ (
    .A(_0365_),
    .Y(_0408_)
  );
  \$_AND_  _2265_ (
    .A(_0358_),
    .B(_0318_),
    .Y(_0409_)
  );
  \$_INV_  _2266_ (
    .A(_0409_),
    .Y(_0410_)
  );
  \$_MUX_  _2267_ (
    .A(_0410_),
    .B(_0408_),
    .S(inst_dest_bin[3]),
    .Y(_0411_)
  );
  \$_AND_  _2268_ (
    .A(_0411_),
    .B(_0407_),
    .Y(_0412_)
  );
  \$_INV_  _2269_ (
    .A(_0323_),
    .Y(_0413_)
  );
  \$_AND_  _2270_ (
    .A(_0317_),
    .B(inst_dest_bin[2]),
    .Y(_0414_)
  );
  \$_AND_  _2271_ (
    .A(_0414_),
    .B(_0344_),
    .Y(_0415_)
  );
  \$_INV_  _2272_ (
    .A(_0415_),
    .Y(_0416_)
  );
  \$_AND_  _2273_ (
    .A(_0416_),
    .B(_0413_),
    .Y(_0417_)
  );
  \$_INV_  _2274_ (
    .A(_0336_),
    .Y(_0418_)
  );
  \$_INV_  _2275_ (
    .A(_0346_),
    .Y(_0419_)
  );
  \$_AND_  _2276_ (
    .A(_0419_),
    .B(_0418_),
    .Y(_0420_)
  );
  \$_AND_  _2277_ (
    .A(_0420_),
    .B(_0417_),
    .Y(_0421_)
  );
  \$_AND_  _2278_ (
    .A(_0421_),
    .B(_0412_),
    .Y(_0422_)
  );
  \$_AND_  _2279_ (
    .A(_0409_),
    .B(inst_dest_bin[3]),
    .Y(_0423_)
  );
  \$_INV_  _2280_ (
    .A(_0423_),
    .Y(_0424_)
  );
  \$_INV_  _2281_ (
    .A(_0322_),
    .Y(_0425_)
  );
  \$_MUX_  _2282_ (
    .A(_0408_),
    .B(_0425_),
    .S(inst_dest_bin[3]),
    .Y(_0426_)
  );
  \$_AND_  _2283_ (
    .A(_0426_),
    .B(_0424_),
    .Y(_0427_)
  );
  \$_AND_  _2284_ (
    .A(_0335_),
    .B(_0317_),
    .Y(_0428_)
  );
  \$_INV_  _2285_ (
    .A(_0428_),
    .Y(_0429_)
  );
  \$_AND_  _2286_ (
    .A(_0345_),
    .B(_0317_),
    .Y(_0430_)
  );
  \$_INV_  _2287_ (
    .A(_0430_),
    .Y(_0431_)
  );
  \$_AND_  _2288_ (
    .A(_0431_),
    .B(_0429_),
    .Y(_0432_)
  );
  \$_AND_  _2289_ (
    .A(_0351_),
    .B(_0317_),
    .Y(_0433_)
  );
  \$_INV_  _2290_ (
    .A(_0433_),
    .Y(_0434_)
  );
  \$_AND_  _2291_ (
    .A(_0359_),
    .B(_0317_),
    .Y(_0435_)
  );
  \$_INV_  _2292_ (
    .A(_0435_),
    .Y(_0436_)
  );
  \$_AND_  _2293_ (
    .A(_0436_),
    .B(_0434_),
    .Y(_0437_)
  );
  \$_AND_  _2294_ (
    .A(_0437_),
    .B(_0432_),
    .Y(_0438_)
  );
  \$_AND_  _2295_ (
    .A(_0438_),
    .B(_0427_),
    .Y(_0439_)
  );
  \$_AND_  _2296_ (
    .A(_0439_),
    .B(_0422_),
    .Y(_0440_)
  );
  \$_AND_  _2297_ (
    .A(_0440_),
    .B(_0338_),
    .Y(_0441_)
  );
  \$_OR_  _2298_ (
    .A(_0441_),
    .B(_0404_),
    .Y(inst_dest[15])
  );
  \$_AND_  _2299_ (
    .A(_0372_),
    .B(_0310_),
    .Y(_0442_)
  );
  \$_AND_  _2300_ (
    .A(_0442_),
    .B(dbg_halt_st),
    .Y(_0443_)
  );
  \$_INV_  _2301_ (
    .A(_0326_),
    .Y(_0444_)
  );
  \$_AND_  _2302_ (
    .A(_0409_),
    .B(_0317_),
    .Y(_0445_)
  );
  \$_OR_  _2303_ (
    .A(_0445_),
    .B(_0444_),
    .Y(_0446_)
  );
  \$_AND_  _2304_ (
    .A(_0446_),
    .B(_0337_),
    .Y(_0447_)
  );
  \$_OR_  _2305_ (
    .A(_0447_),
    .B(_0443_),
    .Y(inst_dest[1])
  );
  \$_AND_  _2306_ (
    .A(_0392_),
    .B(dbg_halt_st),
    .Y(_0448_)
  );
  \$_AND_  _2307_ (
    .A(_0428_),
    .B(_0338_),
    .Y(_0449_)
  );
  \$_OR_  _2308_ (
    .A(_0449_),
    .B(_0448_),
    .Y(inst_dest[2])
  );
  \$_AND_  _2309_ (
    .A(_0394_),
    .B(dbg_halt_st),
    .Y(_0450_)
  );
  \$_AND_  _2310_ (
    .A(_0430_),
    .B(_0338_),
    .Y(_0451_)
  );
  \$_OR_  _2311_ (
    .A(_0451_),
    .B(_0450_),
    .Y(inst_dest[3])
  );
  \$_AND_  _2312_ (
    .A(_0397_),
    .B(dbg_halt_st),
    .Y(_0452_)
  );
  \$_AND_  _2313_ (
    .A(_0433_),
    .B(_0338_),
    .Y(_0453_)
  );
  \$_OR_  _2314_ (
    .A(_0453_),
    .B(_0452_),
    .Y(inst_dest[4])
  );
  \$_AND_  _2315_ (
    .A(_0399_),
    .B(dbg_halt_st),
    .Y(_0454_)
  );
  \$_AND_  _2316_ (
    .A(_0435_),
    .B(_0338_),
    .Y(_0455_)
  );
  \$_OR_  _2317_ (
    .A(_0455_),
    .B(_0454_),
    .Y(inst_dest[5])
  );
  \$_AND_  _2318_ (
    .A(_0362_),
    .B(_0310_),
    .Y(_0456_)
  );
  \$_AND_  _2319_ (
    .A(_0456_),
    .B(dbg_halt_st),
    .Y(_0457_)
  );
  \$_AND_  _2320_ (
    .A(_0365_),
    .B(_0317_),
    .Y(_0458_)
  );
  \$_AND_  _2321_ (
    .A(_0458_),
    .B(_0338_),
    .Y(_0459_)
  );
  \$_OR_  _2322_ (
    .A(_0459_),
    .B(_0457_),
    .Y(inst_dest[6])
  );
  \$_AND_  _2323_ (
    .A(_0378_),
    .B(dbg_halt_st),
    .Y(_0460_)
  );
  \$_AND_  _2324_ (
    .A(_0415_),
    .B(_0338_),
    .Y(_0461_)
  );
  \$_OR_  _2325_ (
    .A(_0461_),
    .B(_0460_),
    .Y(inst_dest[7])
  );
  \$_AND_  _2326_ (
    .A(_0315_),
    .B(dbg_reg_sel[3]),
    .Y(_0462_)
  );
  \$_AND_  _2327_ (
    .A(_0462_),
    .B(dbg_halt_st),
    .Y(_0463_)
  );
  \$_AND_  _2328_ (
    .A(_0322_),
    .B(inst_dest_bin[3]),
    .Y(_0464_)
  );
  \$_AND_  _2329_ (
    .A(_0464_),
    .B(_0338_),
    .Y(_0465_)
  );
  \$_OR_  _2330_ (
    .A(_0465_),
    .B(_0463_),
    .Y(inst_dest[8])
  );
  \$_AND_  _2331_ (
    .A(_0387_),
    .B(dbg_halt_st),
    .Y(_0466_)
  );
  \$_AND_  _2332_ (
    .A(_0423_),
    .B(_0338_),
    .Y(_0467_)
  );
  \$_OR_  _2333_ (
    .A(_0467_),
    .B(_0466_),
    .Y(inst_dest[9])
  );
  \$_INV_  _2334_ (
    .A(inst_src_bin[3]),
    .Y(_0468_)
  );
  \$_INV_  _2335_ (
    .A(inst_src_bin[2]),
    .Y(_0469_)
  );
  \$_INV_  _2336_ (
    .A(inst_src_bin[0]),
    .Y(_0470_)
  );
  \$_INV_  _2337_ (
    .A(inst_src_bin[1]),
    .Y(_0471_)
  );
  \$_AND_  _2338_ (
    .A(_0471_),
    .B(_0470_),
    .Y(_0472_)
  );
  \$_AND_  _2339_ (
    .A(_0472_),
    .B(_0469_),
    .Y(_0473_)
  );
  \$_AND_  _2340_ (
    .A(_0473_),
    .B(_0468_),
    .Y(_0474_)
  );
  \$_AND_  _2341_ (
    .A(_0474_),
    .B(inst_type[2]),
    .Y(_0475_)
  );
  \$_AND_  _2342_ (
    .A(_0325_),
    .B(inst_type[0]),
    .Y(_0476_)
  );
  \$_AND_  _2343_ (
    .A(_0476_),
    .B(_0323_),
    .Y(_0477_)
  );
  \$_OR_  _2344_ (
    .A(_0477_),
    .B(inst_so[7]),
    .Y(_0478_)
  );
  \$_INV_  _2345_ (
    .A(inst_type[2]),
    .Y(_0479_)
  );
  \$_AND_  _2346_ (
    .A(_0479_),
    .B(_0994_),
    .Y(_0480_)
  );
  \$_AND_  _2347_ (
    .A(_0480_),
    .B(_0478_),
    .Y(_0481_)
  );
  \$_OR_  _2348_ (
    .A(_0481_),
    .B(_0475_),
    .Y(inst_src[0])
  );
  \$_AND_  _2349_ (
    .A(inst_src_bin[1]),
    .B(_0470_),
    .Y(_0482_)
  );
  \$_AND_  _2350_ (
    .A(_0482_),
    .B(_0469_),
    .Y(_0483_)
  );
  \$_AND_  _2351_ (
    .A(_0483_),
    .B(inst_src_bin[3]),
    .Y(_0484_)
  );
  \$_AND_  _2352_ (
    .A(_0484_),
    .B(inst_type[2]),
    .Y(_0485_)
  );
  \$_AND_  _2353_ (
    .A(_0480_),
    .B(_0476_),
    .Y(_0486_)
  );
  \$_AND_  _2354_ (
    .A(_0486_),
    .B(_0336_),
    .Y(_0487_)
  );
  \$_OR_  _2355_ (
    .A(_0487_),
    .B(_0485_),
    .Y(inst_src[10])
  );
  \$_AND_  _2356_ (
    .A(inst_src_bin[1]),
    .B(inst_src_bin[0]),
    .Y(_0488_)
  );
  \$_AND_  _2357_ (
    .A(_0488_),
    .B(_0469_),
    .Y(_0489_)
  );
  \$_AND_  _2358_ (
    .A(_0489_),
    .B(inst_src_bin[3]),
    .Y(_0490_)
  );
  \$_AND_  _2359_ (
    .A(_0490_),
    .B(inst_type[2]),
    .Y(_0491_)
  );
  \$_AND_  _2360_ (
    .A(_0486_),
    .B(_0346_),
    .Y(_0492_)
  );
  \$_OR_  _2361_ (
    .A(_0492_),
    .B(_0491_),
    .Y(inst_src[11])
  );
  \$_AND_  _2362_ (
    .A(_0472_),
    .B(inst_src_bin[2]),
    .Y(_0493_)
  );
  \$_AND_  _2363_ (
    .A(_0493_),
    .B(inst_src_bin[3]),
    .Y(_0494_)
  );
  \$_AND_  _2364_ (
    .A(_0494_),
    .B(inst_type[2]),
    .Y(_0495_)
  );
  \$_AND_  _2365_ (
    .A(_0486_),
    .B(_0352_),
    .Y(_0496_)
  );
  \$_OR_  _2366_ (
    .A(_0496_),
    .B(_0495_),
    .Y(inst_src[12])
  );
  \$_AND_  _2367_ (
    .A(_0471_),
    .B(inst_src_bin[0]),
    .Y(_0497_)
  );
  \$_AND_  _2368_ (
    .A(_0497_),
    .B(inst_src_bin[2]),
    .Y(_0498_)
  );
  \$_AND_  _2369_ (
    .A(_0498_),
    .B(inst_src_bin[3]),
    .Y(_0499_)
  );
  \$_AND_  _2370_ (
    .A(_0499_),
    .B(inst_type[2]),
    .Y(_0500_)
  );
  \$_AND_  _2371_ (
    .A(_0486_),
    .B(_0360_),
    .Y(_0501_)
  );
  \$_OR_  _2372_ (
    .A(_0501_),
    .B(_0500_),
    .Y(inst_src[13])
  );
  \$_AND_  _2373_ (
    .A(_0482_),
    .B(inst_src_bin[2]),
    .Y(_0502_)
  );
  \$_AND_  _2374_ (
    .A(_0502_),
    .B(inst_src_bin[3]),
    .Y(_0503_)
  );
  \$_AND_  _2375_ (
    .A(_0503_),
    .B(inst_type[2]),
    .Y(_0504_)
  );
  \$_AND_  _2376_ (
    .A(_0486_),
    .B(_0366_),
    .Y(_0505_)
  );
  \$_OR_  _2377_ (
    .A(_0505_),
    .B(_0504_),
    .Y(inst_src[14])
  );
  \$_INV_  _2378_ (
    .A(_0494_),
    .Y(_0506_)
  );
  \$_INV_  _2379_ (
    .A(_0499_),
    .Y(_0507_)
  );
  \$_AND_  _2380_ (
    .A(_0507_),
    .B(_0506_),
    .Y(_0508_)
  );
  \$_INV_  _2381_ (
    .A(_0502_),
    .Y(_0509_)
  );
  \$_AND_  _2382_ (
    .A(_0497_),
    .B(_0469_),
    .Y(_0510_)
  );
  \$_INV_  _2383_ (
    .A(_0510_),
    .Y(_0511_)
  );
  \$_MUX_  _2384_ (
    .A(_0511_),
    .B(_0509_),
    .S(inst_src_bin[3]),
    .Y(_0512_)
  );
  \$_AND_  _2385_ (
    .A(_0512_),
    .B(_0508_),
    .Y(_0513_)
  );
  \$_INV_  _2386_ (
    .A(_0474_),
    .Y(_0514_)
  );
  \$_AND_  _2387_ (
    .A(_0468_),
    .B(inst_src_bin[2]),
    .Y(_0515_)
  );
  \$_AND_  _2388_ (
    .A(_0515_),
    .B(_0488_),
    .Y(_0516_)
  );
  \$_INV_  _2389_ (
    .A(_0516_),
    .Y(_0517_)
  );
  \$_AND_  _2390_ (
    .A(_0517_),
    .B(inst_type[2]),
    .Y(_0518_)
  );
  \$_AND_  _2391_ (
    .A(_0518_),
    .B(_0514_),
    .Y(_0519_)
  );
  \$_INV_  _2392_ (
    .A(_0484_),
    .Y(_0520_)
  );
  \$_INV_  _2393_ (
    .A(_0490_),
    .Y(_0521_)
  );
  \$_AND_  _2394_ (
    .A(_0521_),
    .B(_0520_),
    .Y(_0522_)
  );
  \$_AND_  _2395_ (
    .A(_0522_),
    .B(_0519_),
    .Y(_0523_)
  );
  \$_AND_  _2396_ (
    .A(_0523_),
    .B(_0513_),
    .Y(_0524_)
  );
  \$_AND_  _2397_ (
    .A(_0510_),
    .B(inst_src_bin[3]),
    .Y(_0525_)
  );
  \$_INV_  _2398_ (
    .A(_0525_),
    .Y(_0526_)
  );
  \$_INV_  _2399_ (
    .A(_0473_),
    .Y(_0527_)
  );
  \$_MUX_  _2400_ (
    .A(_0509_),
    .B(_0527_),
    .S(inst_src_bin[3]),
    .Y(_0528_)
  );
  \$_AND_  _2401_ (
    .A(_0528_),
    .B(_0526_),
    .Y(_0529_)
  );
  \$_AND_  _2402_ (
    .A(_0483_),
    .B(_0468_),
    .Y(_0530_)
  );
  \$_INV_  _2403_ (
    .A(_0530_),
    .Y(_0531_)
  );
  \$_AND_  _2404_ (
    .A(_0489_),
    .B(_0468_),
    .Y(_0532_)
  );
  \$_INV_  _2405_ (
    .A(_0532_),
    .Y(_0533_)
  );
  \$_AND_  _2406_ (
    .A(_0533_),
    .B(_0531_),
    .Y(_0534_)
  );
  \$_AND_  _2407_ (
    .A(_0493_),
    .B(_0468_),
    .Y(_0535_)
  );
  \$_INV_  _2408_ (
    .A(_0535_),
    .Y(_0536_)
  );
  \$_AND_  _2409_ (
    .A(_0498_),
    .B(_0468_),
    .Y(_0537_)
  );
  \$_INV_  _2410_ (
    .A(_0537_),
    .Y(_0538_)
  );
  \$_AND_  _2411_ (
    .A(_0538_),
    .B(_0536_),
    .Y(_0539_)
  );
  \$_AND_  _2412_ (
    .A(_0539_),
    .B(_0534_),
    .Y(_0540_)
  );
  \$_AND_  _2413_ (
    .A(_0540_),
    .B(_0529_),
    .Y(_0541_)
  );
  \$_AND_  _2414_ (
    .A(_0541_),
    .B(_0524_),
    .Y(_0542_)
  );
  \$_AND_  _2415_ (
    .A(_0486_),
    .B(_0440_),
    .Y(_0543_)
  );
  \$_OR_  _2416_ (
    .A(_0543_),
    .B(_0542_),
    .Y(inst_src[15])
  );
  \$_AND_  _2417_ (
    .A(_0510_),
    .B(_0468_),
    .Y(_0544_)
  );
  \$_AND_  _2418_ (
    .A(_0476_),
    .B(_0994_),
    .Y(_0545_)
  );
  \$_AND_  _2419_ (
    .A(_0545_),
    .B(_0445_),
    .Y(_0546_)
  );
  \$_OR_  _2420_ (
    .A(_0546_),
    .B(inst_so[6]),
    .Y(_0547_)
  );
  \$_MUX_  _2421_ (
    .A(_0547_),
    .B(_0544_),
    .S(inst_type[2]),
    .Y(inst_src[1])
  );
  \$_AND_  _2422_ (
    .A(_0530_),
    .B(inst_type[2]),
    .Y(_0548_)
  );
  \$_AND_  _2423_ (
    .A(_0486_),
    .B(_0428_),
    .Y(_0549_)
  );
  \$_OR_  _2424_ (
    .A(_0549_),
    .B(_0548_),
    .Y(inst_src[2])
  );
  \$_AND_  _2425_ (
    .A(_0532_),
    .B(inst_type[2]),
    .Y(_0550_)
  );
  \$_AND_  _2426_ (
    .A(_0486_),
    .B(_0430_),
    .Y(_0551_)
  );
  \$_OR_  _2427_ (
    .A(_0551_),
    .B(_0550_),
    .Y(inst_src[3])
  );
  \$_AND_  _2428_ (
    .A(_0535_),
    .B(inst_type[2]),
    .Y(_0552_)
  );
  \$_AND_  _2429_ (
    .A(_0486_),
    .B(_0433_),
    .Y(_0553_)
  );
  \$_OR_  _2430_ (
    .A(_0553_),
    .B(_0552_),
    .Y(inst_src[4])
  );
  \$_AND_  _2431_ (
    .A(_0537_),
    .B(inst_type[2]),
    .Y(_0554_)
  );
  \$_AND_  _2432_ (
    .A(_0486_),
    .B(_0435_),
    .Y(_0555_)
  );
  \$_OR_  _2433_ (
    .A(_0555_),
    .B(_0554_),
    .Y(inst_src[5])
  );
  \$_AND_  _2434_ (
    .A(_0502_),
    .B(_0468_),
    .Y(_0556_)
  );
  \$_AND_  _2435_ (
    .A(_0556_),
    .B(inst_type[2]),
    .Y(_0557_)
  );
  \$_AND_  _2436_ (
    .A(_0486_),
    .B(_0458_),
    .Y(_0558_)
  );
  \$_OR_  _2437_ (
    .A(_0558_),
    .B(_0557_),
    .Y(inst_src[6])
  );
  \$_AND_  _2438_ (
    .A(_0516_),
    .B(inst_type[2]),
    .Y(_0559_)
  );
  \$_AND_  _2439_ (
    .A(_0486_),
    .B(_0415_),
    .Y(_0560_)
  );
  \$_OR_  _2440_ (
    .A(_0560_),
    .B(_0559_),
    .Y(inst_src[7])
  );
  \$_AND_  _2441_ (
    .A(_0473_),
    .B(inst_src_bin[3]),
    .Y(_0561_)
  );
  \$_AND_  _2442_ (
    .A(_0561_),
    .B(inst_type[2]),
    .Y(_0562_)
  );
  \$_AND_  _2443_ (
    .A(_0486_),
    .B(_0464_),
    .Y(_0563_)
  );
  \$_OR_  _2444_ (
    .A(_0563_),
    .B(_0562_),
    .Y(inst_src[8])
  );
  \$_AND_  _2445_ (
    .A(_0525_),
    .B(inst_type[2]),
    .Y(_0564_)
  );
  \$_AND_  _2446_ (
    .A(_0486_),
    .B(_0423_),
    .Y(_0565_)
  );
  \$_OR_  _2447_ (
    .A(_0565_),
    .B(_0564_),
    .Y(inst_src[9])
  );
  \$_DFF_PP0_  \i_state_reg[0]  /* _2448_ */ (
    .C(mclk),
    .D(_1143_),
    .Q(i_state[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \i_state_reg[1]  /* _2449_ */ (
    .C(mclk),
    .D(_1145_),
    .Q(i_state[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \i_state_reg[2]  /* _2450_ */ (
    .C(mclk),
    .D(_1142_[15]),
    .Q(i_state[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \i_state_reg[3]  /* _2451_ */ (
    .C(mclk),
    .D(_1146_),
    .Q(i_state[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \i_state_reg[4]  /* _2452_ */ (
    .C(mclk),
    .D(_1144_),
    .Q(i_state[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  dbg_halt_st_reg /* _2453_ */ (
    .C(mclk),
    .D(_0000_),
    .Q(dbg_halt_st),
    .R(puc_rst)
  );
  \$_DFF_PP1_  inst_irq_rst_reg /* _2454_ */ (
    .C(mclk),
    .D(_0011_),
    .Q(inst_irq_rst),
    .R(puc_rst)
  );
  \$_DFF_PP1_  \irq_addr_reg[1]  /* _2455_ */ (
    .C(mclk),
    .D(_0019_[0]),
    .Q(irq_addr[1]),
    .R(puc_rst)
  );
  \$_DFF_PP1_  \irq_addr_reg[2]  /* _2456_ */ (
    .C(mclk),
    .D(_0019_[1]),
    .Q(irq_addr[2]),
    .R(puc_rst)
  );
  \$_DFF_PP1_  \irq_addr_reg[3]  /* _2457_ */ (
    .C(mclk),
    .D(_0019_[2]),
    .Q(irq_addr[3]),
    .R(puc_rst)
  );
  \$_DFF_PP1_  \irq_addr_reg[4]  /* _2458_ */ (
    .C(mclk),
    .D(_0019_[3]),
    .Q(irq_addr[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[0]  /* _2459_ */ (
    .C(mclk),
    .D(mab[0]),
    .Q(pc[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[10]  /* _2460_ */ (
    .C(mclk),
    .D(mab[10]),
    .Q(pc[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[11]  /* _2461_ */ (
    .C(mclk),
    .D(mab[11]),
    .Q(pc[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[12]  /* _2462_ */ (
    .C(mclk),
    .D(mab[12]),
    .Q(pc[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[13]  /* _2463_ */ (
    .C(mclk),
    .D(mab[13]),
    .Q(pc[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[14]  /* _2464_ */ (
    .C(mclk),
    .D(mab[14]),
    .Q(pc[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[15]  /* _2465_ */ (
    .C(mclk),
    .D(mab[15]),
    .Q(pc[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[1]  /* _2466_ */ (
    .C(mclk),
    .D(mab[1]),
    .Q(pc[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[2]  /* _2467_ */ (
    .C(mclk),
    .D(mab[2]),
    .Q(pc[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[3]  /* _2468_ */ (
    .C(mclk),
    .D(mab[3]),
    .Q(pc[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[4]  /* _2469_ */ (
    .C(mclk),
    .D(mab[4]),
    .Q(pc[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[5]  /* _2470_ */ (
    .C(mclk),
    .D(mab[5]),
    .Q(pc[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[6]  /* _2471_ */ (
    .C(mclk),
    .D(mab[6]),
    .Q(pc[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[7]  /* _2472_ */ (
    .C(mclk),
    .D(mab[7]),
    .Q(pc[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[8]  /* _2473_ */ (
    .C(mclk),
    .D(mab[8]),
    .Q(pc[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pc_reg[9]  /* _2474_ */ (
    .C(mclk),
    .D(mab[9]),
    .Q(pc[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  pmem_busy_reg /* _2475_ */ (
    .C(mclk),
    .D(fe_pmem_wait),
    .Q(pmem_busy),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[0]  /* _2476_ */ (
    .C(mclk),
    .D(_0014_[0]),
    .Q(inst_sext[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[10]  /* _2477_ */ (
    .C(mclk),
    .D(_0014_[10]),
    .Q(inst_sext[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[11]  /* _2478_ */ (
    .C(mclk),
    .D(_0014_[11]),
    .Q(inst_sext[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[12]  /* _2479_ */ (
    .C(mclk),
    .D(_0014_[12]),
    .Q(inst_sext[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[13]  /* _2480_ */ (
    .C(mclk),
    .D(_0014_[13]),
    .Q(inst_sext[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[14]  /* _2481_ */ (
    .C(mclk),
    .D(_0014_[14]),
    .Q(inst_sext[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[15]  /* _2482_ */ (
    .C(mclk),
    .D(_0014_[15]),
    .Q(inst_sext[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[1]  /* _2483_ */ (
    .C(mclk),
    .D(_0014_[1]),
    .Q(inst_sext[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[2]  /* _2484_ */ (
    .C(mclk),
    .D(_0014_[2]),
    .Q(inst_sext[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[3]  /* _2485_ */ (
    .C(mclk),
    .D(_0014_[3]),
    .Q(inst_sext[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[4]  /* _2486_ */ (
    .C(mclk),
    .D(_0014_[4]),
    .Q(inst_sext[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[5]  /* _2487_ */ (
    .C(mclk),
    .D(_0014_[5]),
    .Q(inst_sext[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[6]  /* _2488_ */ (
    .C(mclk),
    .D(_0014_[6]),
    .Q(inst_sext[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[7]  /* _2489_ */ (
    .C(mclk),
    .D(_0014_[7]),
    .Q(inst_sext[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[8]  /* _2490_ */ (
    .C(mclk),
    .D(_0014_[8]),
    .Q(inst_sext[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sext_reg[9]  /* _2491_ */ (
    .C(mclk),
    .D(_0014_[9]),
    .Q(inst_sext[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[0]  /* _2492_ */ (
    .C(mclk),
    .D(_0010_[0]),
    .Q(inst_dext[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[10]  /* _2493_ */ (
    .C(mclk),
    .D(_0010_[10]),
    .Q(inst_dext[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[11]  /* _2494_ */ (
    .C(mclk),
    .D(_0010_[11]),
    .Q(inst_dext[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[12]  /* _2495_ */ (
    .C(mclk),
    .D(_0010_[12]),
    .Q(inst_dext[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[13]  /* _2496_ */ (
    .C(mclk),
    .D(_0010_[13]),
    .Q(inst_dext[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[14]  /* _2497_ */ (
    .C(mclk),
    .D(_0010_[14]),
    .Q(inst_dext[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[15]  /* _2498_ */ (
    .C(mclk),
    .D(_0010_[15]),
    .Q(inst_dext[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[1]  /* _2499_ */ (
    .C(mclk),
    .D(_0010_[1]),
    .Q(inst_dext[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[2]  /* _2500_ */ (
    .C(mclk),
    .D(_0010_[2]),
    .Q(inst_dext[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[3]  /* _2501_ */ (
    .C(mclk),
    .D(_0010_[3]),
    .Q(inst_dext[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[4]  /* _2502_ */ (
    .C(mclk),
    .D(_0010_[4]),
    .Q(inst_dext[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[5]  /* _2503_ */ (
    .C(mclk),
    .D(_0010_[5]),
    .Q(inst_dext[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[6]  /* _2504_ */ (
    .C(mclk),
    .D(_0010_[6]),
    .Q(inst_dext[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[7]  /* _2505_ */ (
    .C(mclk),
    .D(_0010_[7]),
    .Q(inst_dext[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[8]  /* _2506_ */ (
    .C(mclk),
    .D(_0010_[8]),
    .Q(inst_dext[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dext_reg[9]  /* _2507_ */ (
    .C(mclk),
    .D(_0010_[9]),
    .Q(inst_dext[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_type_reg[0]  /* _2508_ */ (
    .C(mclk),
    .D(_0018_[0]),
    .Q(inst_type[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_type_reg[1]  /* _2509_ */ (
    .C(mclk),
    .D(_0018_[1]),
    .Q(inst_type[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_type_reg[2]  /* _2510_ */ (
    .C(mclk),
    .D(_0018_[2]),
    .Q(inst_type[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[0]  /* _2511_ */ (
    .C(mclk),
    .D(_0015_[0]),
    .Q(inst_so[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[1]  /* _2512_ */ (
    .C(mclk),
    .D(_0015_[1]),
    .Q(inst_so[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[2]  /* _2513_ */ (
    .C(mclk),
    .D(_0015_[2]),
    .Q(inst_so[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[3]  /* _2514_ */ (
    .C(mclk),
    .D(_0015_[3]),
    .Q(inst_so[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[4]  /* _2515_ */ (
    .C(mclk),
    .D(_0015_[4]),
    .Q(inst_so[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[5]  /* _2516_ */ (
    .C(mclk),
    .D(_0015_[5]),
    .Q(inst_so[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[6]  /* _2517_ */ (
    .C(mclk),
    .D(_0015_[6]),
    .Q(inst_so[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_so_reg[7]  /* _2518_ */ (
    .C(mclk),
    .D(_0015_[7]),
    .Q(inst_so[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_jmp_bin_reg[0]  /* _2519_ */ (
    .C(mclk),
    .D(_0012_[0]),
    .Q(inst_jmp_bin[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_jmp_bin_reg[1]  /* _2520_ */ (
    .C(mclk),
    .D(_0012_[1]),
    .Q(inst_jmp_bin[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_jmp_bin_reg[2]  /* _2521_ */ (
    .C(mclk),
    .D(_0012_[2]),
    .Q(inst_jmp_bin[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  inst_mov_reg /* _2522_ */ (
    .C(mclk),
    .D(_0013_),
    .Q(inst_mov),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dest_bin_reg[0]  /* _2523_ */ (
    .C(mclk),
    .D(_0009_[0]),
    .Q(inst_dest_bin[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dest_bin_reg[1]  /* _2524_ */ (
    .C(mclk),
    .D(_0009_[1]),
    .Q(inst_dest_bin[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dest_bin_reg[2]  /* _2525_ */ (
    .C(mclk),
    .D(_0009_[2]),
    .Q(inst_dest_bin[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_dest_bin_reg[3]  /* _2526_ */ (
    .C(mclk),
    .D(_0009_[3]),
    .Q(inst_dest_bin[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_src_bin_reg[0]  /* _2527_ */ (
    .C(mclk),
    .D(_0016_[0]),
    .Q(inst_src_bin[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_src_bin_reg[1]  /* _2528_ */ (
    .C(mclk),
    .D(_0016_[1]),
    .Q(inst_src_bin[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_src_bin_reg[2]  /* _2529_ */ (
    .C(mclk),
    .D(_0016_[2]),
    .Q(inst_src_bin[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_src_bin_reg[3]  /* _2530_ */ (
    .C(mclk),
    .D(_0016_[3]),
    .Q(inst_src_bin[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[0]  /* _2531_ */ (
    .C(mclk),
    .D(_0007_[0]),
    .Q(inst_as[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[1]  /* _2532_ */ (
    .C(mclk),
    .D(_0007_[1]),
    .Q(inst_as[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[2]  /* _2533_ */ (
    .C(mclk),
    .D(_0007_[2]),
    .Q(inst_as[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[3]  /* _2534_ */ (
    .C(mclk),
    .D(_0007_[3]),
    .Q(inst_as[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[4]  /* _2535_ */ (
    .C(mclk),
    .D(_0007_[4]),
    .Q(inst_as[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[5]  /* _2536_ */ (
    .C(mclk),
    .D(_0007_[5]),
    .Q(inst_as[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[6]  /* _2537_ */ (
    .C(mclk),
    .D(_0007_[6]),
    .Q(inst_as[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_as_reg[7]  /* _2538_ */ (
    .C(mclk),
    .D(_0007_[7]),
    .Q(inst_as[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[0]  /* _2539_ */ (
    .C(mclk),
    .D(_0005_[0]),
    .Q(inst_ad[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[1]  /* _2540_ */ (
    .C(mclk),
    .D(_0005_[1]),
    .Q(inst_ad[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[2]  /* _2541_ */ (
    .C(mclk),
    .D(_0005_[2]),
    .Q(inst_ad[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[3]  /* _2542_ */ (
    .C(mclk),
    .D(_0005_[3]),
    .Q(inst_ad[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[4]  /* _2543_ */ (
    .C(mclk),
    .D(_0005_[4]),
    .Q(inst_ad[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[5]  /* _2544_ */ (
    .C(mclk),
    .D(_0005_[5]),
    .Q(inst_ad[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[6]  /* _2545_ */ (
    .C(mclk),
    .D(_0005_[6]),
    .Q(inst_ad[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_ad_reg[7]  /* _2546_ */ (
    .C(mclk),
    .D(_0005_[7]),
    .Q(inst_ad[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  inst_bw_reg /* _2547_ */ (
    .C(mclk),
    .D(_0008_),
    .Q(inst_bw),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sz_reg[0]  /* _2548_ */ (
    .C(mclk),
    .D(_0017_[0]),
    .Q(inst_sz[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_sz_reg[1]  /* _2549_ */ (
    .C(mclk),
    .D(_0017_[1]),
    .Q(inst_sz[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  exec_jmp_reg /* _2550_ */ (
    .C(mclk),
    .D(_0003_),
    .Q(exec_jmp),
    .R(puc_rst)
  );
  \$_DFF_PP0_  exec_dst_wr_reg /* _2551_ */ (
    .C(mclk),
    .D(_0002_),
    .Q(exec_dst_wr),
    .R(puc_rst)
  );
  \$_DFF_PP0_  exec_src_wr_reg /* _2552_ */ (
    .C(mclk),
    .D(_0004_),
    .Q(exec_src_wr),
    .R(puc_rst)
  );
  \$_DFF_PP0_  exec_dext_rdy_reg /* _2553_ */ (
    .C(mclk),
    .D(_0001_),
    .Q(exec_dext_rdy),
    .R(puc_rst)
  );
  \$_DFF_PP1_  \e_state_reg[0]  /* _2554_ */ (
    .C(mclk),
    .D(e_state_nxt[0]),
    .Q(e_state[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \e_state_reg[1]  /* _2555_ */ (
    .C(mclk),
    .D(e_state_nxt[1]),
    .Q(e_state[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \e_state_reg[2]  /* _2556_ */ (
    .C(mclk),
    .D(e_state_nxt[2]),
    .Q(e_state[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \e_state_reg[3]  /* _2557_ */ (
    .C(mclk),
    .D(e_state_nxt[3]),
    .Q(e_state[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[0]  /* _2558_ */ (
    .C(mclk),
    .D(_0006_[0]),
    .Q(inst_alu[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[10]  /* _2559_ */ (
    .C(mclk),
    .D(_0006_[10]),
    .Q(inst_alu[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[11]  /* _2560_ */ (
    .C(mclk),
    .D(_0006_[11]),
    .Q(inst_alu[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[1]  /* _2561_ */ (
    .C(mclk),
    .D(_0006_[1]),
    .Q(inst_alu[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[2]  /* _2562_ */ (
    .C(mclk),
    .D(_0006_[2]),
    .Q(inst_alu[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[3]  /* _2563_ */ (
    .C(mclk),
    .D(_0006_[3]),
    .Q(inst_alu[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[4]  /* _2564_ */ (
    .C(mclk),
    .D(_0006_[4]),
    .Q(inst_alu[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[5]  /* _2565_ */ (
    .C(mclk),
    .D(_0006_[5]),
    .Q(inst_alu[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[6]  /* _2566_ */ (
    .C(mclk),
    .D(_0006_[6]),
    .Q(inst_alu[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[7]  /* _2567_ */ (
    .C(mclk),
    .D(_0006_[7]),
    .Q(inst_alu[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[8]  /* _2568_ */ (
    .C(mclk),
    .D(_0006_[8]),
    .Q(inst_alu[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \inst_alu_reg[9]  /* _2569_ */ (
    .C(mclk),
    .D(_0006_[9]),
    .Q(inst_alu[9]),
    .R(puc_rst)
  );
  assign dest_reg = mdb_in[3:0];
  assign ext_nxt[0] = mdb_in[0];
  assign ir = mdb_in;
  assign irq_acc_all[13:0] = irq_acc;
  assign { irq_addr[15:5], irq_addr[0] } = 12'b111111111110;
  assign irq_num = irq_addr[4:1];
  assign mclk_decode = mclk;
  assign mclk_enable = 1'b1;
  assign mclk_inst_dext = mclk;
  assign mclk_inst_sext = mclk;
  assign mclk_irq_num = mclk;
  assign mclk_pc = mclk;
  assign mclk_wkup = 1'b1;
  assign nmi_acc = irq_acc_all[14];
  assign pc_incr[0] = pc[0];
  assign pc_nxt = mab;
endmodule

module omsp_mem_backbone(dbg_mem_din, dmem_addr, dmem_cen, dmem_din, dmem_wen, eu_mdb_in, fe_mdb_in, fe_pmem_wait, per_addr, per_din, per_we, per_en, pmem_addr, pmem_cen, pmem_din, pmem_wen, dbg_halt_st, dbg_mem_addr, dbg_mem_dout, dbg_mem_en, dbg_mem_wr, dmem_dout, eu_mab, eu_mb_en, eu_mb_wr, eu_mdb_out, fe_mab, fe_mb_en, mclk, per_dout, pmem_dout, puc_rst, scan_enable);
  wire [1:0] _000_;
  wire [1:0] _001_;
  wire [15:0] _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  wire _335_;
  wire _336_;
  wire _337_;
  wire _338_;
  wire _339_;
  wire _340_;
  wire _341_;
  wire _342_;
  wire _343_;
  wire _344_;
  wire _345_;
  input dbg_halt_st;
  input [15:0] dbg_mem_addr;
  output [15:0] dbg_mem_din;
  wire [1:0] dbg_mem_din_sel;
  input [15:0] dbg_mem_dout;
  input dbg_mem_en;
  input [1:0] dbg_mem_wr;
  wire dbg_per_en;
  output [5:0] dmem_addr;
  output dmem_cen;
  output [15:0] dmem_din;
  input [15:0] dmem_dout;
  output [1:0] dmem_wen;
  input [14:0] eu_mab;
  input eu_mb_en;
  input [1:0] eu_mb_wr;
  output [15:0] eu_mdb_in;
  wire [1:0] eu_mdb_in_sel;
  input [15:0] eu_mdb_out;
  input [14:0] fe_mab;
  input fe_mb_en;
  output [15:0] fe_mdb_in;
  wire fe_pmem_cen;
  wire fe_pmem_cen_dly;
  output fe_pmem_wait;
  input mclk;
  wire mclk_bckup;
  output [13:0] per_addr;
  wire [14:0] per_addr_ful;
  wire [7:0] per_addr_mux;
  output [15:0] per_din;
  input [15:0] per_dout;
  wire [15:0] per_dout_val;
  output per_en;
  output [1:0] per_we;
  output [9:0] pmem_addr;
  output pmem_cen;
  output [15:0] pmem_din;
  input [15:0] pmem_dout;
  wire [15:0] pmem_dout_bckup;
  wire pmem_dout_bckup_sel;
  output [1:0] pmem_wen;
  input puc_rst;
  input scan_enable;
  \$_INV_  _346_ (
    .A(dbg_mem_addr[15]),
    .Y(_004_)
  );
  \$_INV_  _347_ (
    .A(dbg_mem_addr[14]),
    .Y(_005_)
  );
  \$_INV_  _348_ (
    .A(dbg_mem_addr[13]),
    .Y(_006_)
  );
  \$_INV_  _349_ (
    .A(dbg_mem_addr[12]),
    .Y(_007_)
  );
  \$_INV_  _350_ (
    .A(dbg_mem_addr[11]),
    .Y(_008_)
  );
  \$_INV_  _351_ (
    .A(dbg_mem_addr[10]),
    .Y(_009_)
  );
  \$_INV_  _352_ (
    .A(dbg_mem_addr[8]),
    .Y(_010_)
  );
  \$_INV_  _353_ (
    .A(dbg_mem_addr[7]),
    .Y(_011_)
  );
  \$_INV_  _354_ (
    .A(dbg_mem_addr[6]),
    .Y(_012_)
  );
  \$_INV_  _355_ (
    .A(dbg_mem_addr[5]),
    .Y(_013_)
  );
  \$_INV_  _356_ (
    .A(dbg_mem_addr[4]),
    .Y(_014_)
  );
  \$_INV_  _357_ (
    .A(dbg_mem_addr[3]),
    .Y(_015_)
  );
  \$_INV_  _358_ (
    .A(dbg_mem_addr[1]),
    .Y(_016_)
  );
  \$_INV_  _359_ (
    .A(dbg_mem_addr[2]),
    .Y(_017_)
  );
  \$_AND_  _360_ (
    .A(_017_),
    .B(_016_),
    .Y(_018_)
  );
  \$_AND_  _361_ (
    .A(_018_),
    .B(_015_),
    .Y(_019_)
  );
  \$_AND_  _362_ (
    .A(_019_),
    .B(_014_),
    .Y(_020_)
  );
  \$_AND_  _363_ (
    .A(_020_),
    .B(_013_),
    .Y(_021_)
  );
  \$_AND_  _364_ (
    .A(_021_),
    .B(_012_),
    .Y(_022_)
  );
  \$_AND_  _365_ (
    .A(_022_),
    .B(_011_),
    .Y(_023_)
  );
  \$_AND_  _366_ (
    .A(_023_),
    .B(_010_),
    .Y(_024_)
  );
  \$_INV_  _367_ (
    .A(_024_),
    .Y(_025_)
  );
  \$_AND_  _368_ (
    .A(_025_),
    .B(dbg_mem_addr[9]),
    .Y(_026_)
  );
  \$_INV_  _369_ (
    .A(_026_),
    .Y(_027_)
  );
  \$_AND_  _370_ (
    .A(_027_),
    .B(_009_),
    .Y(_028_)
  );
  \$_AND_  _371_ (
    .A(_028_),
    .B(_008_),
    .Y(_029_)
  );
  \$_AND_  _372_ (
    .A(_029_),
    .B(_007_),
    .Y(_030_)
  );
  \$_AND_  _373_ (
    .A(_030_),
    .B(_006_),
    .Y(_031_)
  );
  \$_AND_  _374_ (
    .A(_031_),
    .B(_005_),
    .Y(_032_)
  );
  \$_AND_  _375_ (
    .A(_032_),
    .B(_004_),
    .Y(_033_)
  );
  \$_AND_  _376_ (
    .A(_027_),
    .B(dbg_mem_addr[10]),
    .Y(_034_)
  );
  \$_INV_  _377_ (
    .A(dbg_mem_addr[9]),
    .Y(_035_)
  );
  \$_XOR_  _378_ (
    .A(_024_),
    .B(_035_),
    .Y(_036_)
  );
  \$_AND_  _379_ (
    .A(_036_),
    .B(_024_),
    .Y(_037_)
  );
  \$_INV_  _380_ (
    .A(_037_),
    .Y(_038_)
  );
  \$_OR_  _381_ (
    .A(_038_),
    .B(_034_),
    .Y(_039_)
  );
  \$_XOR_  _382_ (
    .A(_028_),
    .B(dbg_mem_addr[11]),
    .Y(_040_)
  );
  \$_INV_  _383_ (
    .A(_040_),
    .Y(_041_)
  );
  \$_OR_  _384_ (
    .A(_041_),
    .B(_039_),
    .Y(_042_)
  );
  \$_XOR_  _385_ (
    .A(_029_),
    .B(dbg_mem_addr[12]),
    .Y(_043_)
  );
  \$_INV_  _386_ (
    .A(_043_),
    .Y(_044_)
  );
  \$_OR_  _387_ (
    .A(_044_),
    .B(_042_),
    .Y(_045_)
  );
  \$_XOR_  _388_ (
    .A(_030_),
    .B(dbg_mem_addr[13]),
    .Y(_046_)
  );
  \$_INV_  _389_ (
    .A(_046_),
    .Y(_047_)
  );
  \$_OR_  _390_ (
    .A(_047_),
    .B(_045_),
    .Y(_048_)
  );
  \$_XOR_  _391_ (
    .A(_031_),
    .B(dbg_mem_addr[14]),
    .Y(_049_)
  );
  \$_INV_  _392_ (
    .A(_049_),
    .Y(_050_)
  );
  \$_OR_  _393_ (
    .A(_050_),
    .B(_048_),
    .Y(_051_)
  );
  \$_INV_  _394_ (
    .A(_033_),
    .Y(_052_)
  );
  \$_OR_  _395_ (
    .A(_052_),
    .B(_051_),
    .Y(_053_)
  );
  \$_AND_  _396_ (
    .A(_053_),
    .B(_033_),
    .Y(_054_)
  );
  \$_AND_  _397_ (
    .A(_010_),
    .B(_011_),
    .Y(_055_)
  );
  \$_INV_  _398_ (
    .A(_055_),
    .Y(_056_)
  );
  \$_AND_  _399_ (
    .A(_009_),
    .B(dbg_mem_addr[9]),
    .Y(_057_)
  );
  \$_AND_  _400_ (
    .A(_057_),
    .B(_056_),
    .Y(_058_)
  );
  \$_OR_  _401_ (
    .A(_058_),
    .B(dbg_mem_addr[10]),
    .Y(_059_)
  );
  \$_OR_  _402_ (
    .A(_059_),
    .B(dbg_mem_addr[11]),
    .Y(_060_)
  );
  \$_OR_  _403_ (
    .A(_060_),
    .B(dbg_mem_addr[12]),
    .Y(_061_)
  );
  \$_OR_  _404_ (
    .A(_061_),
    .B(dbg_mem_addr[13]),
    .Y(_062_)
  );
  \$_OR_  _405_ (
    .A(_062_),
    .B(dbg_mem_addr[14]),
    .Y(_063_)
  );
  \$_AND_  _406_ (
    .A(_063_),
    .B(_004_),
    .Y(_064_)
  );
  \$_INV_  _407_ (
    .A(_064_),
    .Y(_065_)
  );
  \$_AND_  _408_ (
    .A(_004_),
    .B(dbg_mem_en),
    .Y(_066_)
  );
  \$_AND_  _409_ (
    .A(_066_),
    .B(_065_),
    .Y(_067_)
  );
  \$_INV_  _410_ (
    .A(_067_),
    .Y(_068_)
  );
  \$_OR_  _411_ (
    .A(_068_),
    .B(_054_),
    .Y(_069_)
  );
  \$_INV_  _412_ (
    .A(eu_mab[14]),
    .Y(_070_)
  );
  \$_INV_  _413_ (
    .A(eu_mab[13]),
    .Y(_071_)
  );
  \$_INV_  _414_ (
    .A(eu_mab[12]),
    .Y(_072_)
  );
  \$_INV_  _415_ (
    .A(eu_mab[11]),
    .Y(_073_)
  );
  \$_INV_  _416_ (
    .A(eu_mab[10]),
    .Y(_074_)
  );
  \$_INV_  _417_ (
    .A(eu_mab[9]),
    .Y(_075_)
  );
  \$_OR_  _418_ (
    .A(eu_mab[1]),
    .B(eu_mab[0]),
    .Y(_076_)
  );
  \$_OR_  _419_ (
    .A(_076_),
    .B(eu_mab[2]),
    .Y(_077_)
  );
  \$_OR_  _420_ (
    .A(_077_),
    .B(eu_mab[3]),
    .Y(_078_)
  );
  \$_OR_  _421_ (
    .A(_078_),
    .B(eu_mab[4]),
    .Y(_079_)
  );
  \$_OR_  _422_ (
    .A(_079_),
    .B(eu_mab[5]),
    .Y(_080_)
  );
  \$_OR_  _423_ (
    .A(_080_),
    .B(eu_mab[6]),
    .Y(_081_)
  );
  \$_OR_  _424_ (
    .A(_081_),
    .B(eu_mab[7]),
    .Y(_082_)
  );
  \$_AND_  _425_ (
    .A(_082_),
    .B(eu_mab[8]),
    .Y(_083_)
  );
  \$_INV_  _426_ (
    .A(_083_),
    .Y(_084_)
  );
  \$_AND_  _427_ (
    .A(_084_),
    .B(_075_),
    .Y(_085_)
  );
  \$_AND_  _428_ (
    .A(_085_),
    .B(_074_),
    .Y(_086_)
  );
  \$_AND_  _429_ (
    .A(_086_),
    .B(_073_),
    .Y(_087_)
  );
  \$_AND_  _430_ (
    .A(_087_),
    .B(_072_),
    .Y(_088_)
  );
  \$_AND_  _431_ (
    .A(_088_),
    .B(_071_),
    .Y(_089_)
  );
  \$_AND_  _432_ (
    .A(_089_),
    .B(_070_),
    .Y(_090_)
  );
  \$_AND_  _433_ (
    .A(_084_),
    .B(eu_mab[9]),
    .Y(_091_)
  );
  \$_INV_  _434_ (
    .A(eu_mab[8]),
    .Y(_092_)
  );
  \$_XOR_  _435_ (
    .A(_082_),
    .B(_092_),
    .Y(_093_)
  );
  \$_OR_  _436_ (
    .A(_093_),
    .B(_082_),
    .Y(_094_)
  );
  \$_OR_  _437_ (
    .A(_094_),
    .B(_091_),
    .Y(_095_)
  );
  \$_XOR_  _438_ (
    .A(_085_),
    .B(_074_),
    .Y(_096_)
  );
  \$_OR_  _439_ (
    .A(_096_),
    .B(_095_),
    .Y(_097_)
  );
  \$_XOR_  _440_ (
    .A(_086_),
    .B(_073_),
    .Y(_098_)
  );
  \$_OR_  _441_ (
    .A(_098_),
    .B(_097_),
    .Y(_099_)
  );
  \$_XOR_  _442_ (
    .A(_087_),
    .B(_072_),
    .Y(_100_)
  );
  \$_OR_  _443_ (
    .A(_100_),
    .B(_099_),
    .Y(_101_)
  );
  \$_XOR_  _444_ (
    .A(_088_),
    .B(_071_),
    .Y(_102_)
  );
  \$_OR_  _445_ (
    .A(_102_),
    .B(_101_),
    .Y(_103_)
  );
  \$_INV_  _446_ (
    .A(_089_),
    .Y(_104_)
  );
  \$_OR_  _447_ (
    .A(_104_),
    .B(eu_mab[14]),
    .Y(_105_)
  );
  \$_OR_  _448_ (
    .A(_105_),
    .B(_103_),
    .Y(_106_)
  );
  \$_AND_  _449_ (
    .A(_106_),
    .B(_090_),
    .Y(_107_)
  );
  \$_OR_  _450_ (
    .A(eu_mab[7]),
    .B(eu_mab[6]),
    .Y(_108_)
  );
  \$_AND_  _451_ (
    .A(_075_),
    .B(eu_mab[8]),
    .Y(_109_)
  );
  \$_AND_  _452_ (
    .A(_109_),
    .B(_108_),
    .Y(_110_)
  );
  \$_OR_  _453_ (
    .A(_110_),
    .B(eu_mab[9]),
    .Y(_111_)
  );
  \$_OR_  _454_ (
    .A(_111_),
    .B(eu_mab[10]),
    .Y(_112_)
  );
  \$_OR_  _455_ (
    .A(_112_),
    .B(eu_mab[11]),
    .Y(_113_)
  );
  \$_OR_  _456_ (
    .A(_113_),
    .B(eu_mab[12]),
    .Y(_114_)
  );
  \$_OR_  _457_ (
    .A(_114_),
    .B(eu_mab[13]),
    .Y(_115_)
  );
  \$_AND_  _458_ (
    .A(_115_),
    .B(_070_),
    .Y(_116_)
  );
  \$_AND_  _459_ (
    .A(_070_),
    .B(eu_mb_en),
    .Y(_117_)
  );
  \$_INV_  _460_ (
    .A(_117_),
    .Y(_118_)
  );
  \$_OR_  _461_ (
    .A(_118_),
    .B(_116_),
    .Y(_119_)
  );
  \$_OR_  _462_ (
    .A(_119_),
    .B(_107_),
    .Y(_120_)
  );
  \$_AND_  _463_ (
    .A(_120_),
    .B(_069_),
    .Y(dmem_cen)
  );
  \$_INV_  _464_ (
    .A(fe_mb_en),
    .Y(_121_)
  );
  \$_OR_  _465_ (
    .A(fe_mab[1]),
    .B(fe_mab[0]),
    .Y(_122_)
  );
  \$_OR_  _466_ (
    .A(_122_),
    .B(fe_mab[2]),
    .Y(_123_)
  );
  \$_OR_  _467_ (
    .A(_123_),
    .B(fe_mab[3]),
    .Y(_124_)
  );
  \$_OR_  _468_ (
    .A(_124_),
    .B(fe_mab[4]),
    .Y(_125_)
  );
  \$_OR_  _469_ (
    .A(_125_),
    .B(fe_mab[5]),
    .Y(_126_)
  );
  \$_OR_  _470_ (
    .A(_126_),
    .B(fe_mab[6]),
    .Y(_127_)
  );
  \$_OR_  _471_ (
    .A(_127_),
    .B(fe_mab[7]),
    .Y(_128_)
  );
  \$_OR_  _472_ (
    .A(_128_),
    .B(fe_mab[8]),
    .Y(_129_)
  );
  \$_OR_  _473_ (
    .A(_129_),
    .B(fe_mab[9]),
    .Y(_130_)
  );
  \$_AND_  _474_ (
    .A(_130_),
    .B(fe_mab[10]),
    .Y(_131_)
  );
  \$_AND_  _475_ (
    .A(_131_),
    .B(fe_mab[11]),
    .Y(_132_)
  );
  \$_AND_  _476_ (
    .A(_132_),
    .B(fe_mab[12]),
    .Y(_133_)
  );
  \$_AND_  _477_ (
    .A(_133_),
    .B(fe_mab[13]),
    .Y(_134_)
  );
  \$_AND_  _478_ (
    .A(_134_),
    .B(fe_mab[14]),
    .Y(_135_)
  );
  \$_INV_  _479_ (
    .A(_135_),
    .Y(_136_)
  );
  \$_OR_  _480_ (
    .A(_134_),
    .B(fe_mab[14]),
    .Y(_137_)
  );
  \$_INV_  _481_ (
    .A(_137_),
    .Y(_138_)
  );
  \$_OR_  _482_ (
    .A(_133_),
    .B(fe_mab[13]),
    .Y(_139_)
  );
  \$_INV_  _483_ (
    .A(_139_),
    .Y(_140_)
  );
  \$_OR_  _484_ (
    .A(_132_),
    .B(fe_mab[12]),
    .Y(_141_)
  );
  \$_INV_  _485_ (
    .A(_141_),
    .Y(_142_)
  );
  \$_INV_  _486_ (
    .A(fe_mab[11]),
    .Y(_143_)
  );
  \$_INV_  _487_ (
    .A(fe_mab[10]),
    .Y(_144_)
  );
  \$_INV_  _488_ (
    .A(fe_mab[9]),
    .Y(_145_)
  );
  \$_INV_  _489_ (
    .A(fe_mab[8]),
    .Y(_146_)
  );
  \$_INV_  _490_ (
    .A(fe_mab[7]),
    .Y(_147_)
  );
  \$_INV_  _491_ (
    .A(fe_mab[6]),
    .Y(_148_)
  );
  \$_INV_  _492_ (
    .A(fe_mab[5]),
    .Y(_149_)
  );
  \$_INV_  _493_ (
    .A(fe_mab[4]),
    .Y(_150_)
  );
  \$_INV_  _494_ (
    .A(fe_mab[3]),
    .Y(_151_)
  );
  \$_INV_  _495_ (
    .A(fe_mab[2]),
    .Y(_152_)
  );
  \$_INV_  _496_ (
    .A(fe_mab[0]),
    .Y(_153_)
  );
  \$_INV_  _497_ (
    .A(fe_mab[1]),
    .Y(_154_)
  );
  \$_AND_  _498_ (
    .A(_154_),
    .B(_153_),
    .Y(_155_)
  );
  \$_AND_  _499_ (
    .A(_155_),
    .B(_152_),
    .Y(_156_)
  );
  \$_AND_  _500_ (
    .A(_156_),
    .B(_151_),
    .Y(_157_)
  );
  \$_AND_  _501_ (
    .A(_157_),
    .B(_150_),
    .Y(_158_)
  );
  \$_AND_  _502_ (
    .A(_158_),
    .B(_149_),
    .Y(_159_)
  );
  \$_AND_  _503_ (
    .A(_159_),
    .B(_148_),
    .Y(_160_)
  );
  \$_AND_  _504_ (
    .A(_160_),
    .B(_147_),
    .Y(_161_)
  );
  \$_AND_  _505_ (
    .A(_161_),
    .B(_146_),
    .Y(_162_)
  );
  \$_AND_  _506_ (
    .A(_162_),
    .B(_145_),
    .Y(_163_)
  );
  \$_OR_  _507_ (
    .A(_163_),
    .B(_144_),
    .Y(_164_)
  );
  \$_AND_  _508_ (
    .A(_164_),
    .B(_143_),
    .Y(_165_)
  );
  \$_XOR_  _509_ (
    .A(_130_),
    .B(_144_),
    .Y(_166_)
  );
  \$_OR_  _510_ (
    .A(_166_),
    .B(_130_),
    .Y(_167_)
  );
  \$_OR_  _511_ (
    .A(_167_),
    .B(_165_),
    .Y(_168_)
  );
  \$_OR_  _512_ (
    .A(_168_),
    .B(_132_),
    .Y(_169_)
  );
  \$_OR_  _513_ (
    .A(_169_),
    .B(_142_),
    .Y(_170_)
  );
  \$_OR_  _514_ (
    .A(_170_),
    .B(_133_),
    .Y(_171_)
  );
  \$_OR_  _515_ (
    .A(_171_),
    .B(_140_),
    .Y(_172_)
  );
  \$_OR_  _516_ (
    .A(_172_),
    .B(_134_),
    .Y(_173_)
  );
  \$_OR_  _517_ (
    .A(_173_),
    .B(_138_),
    .Y(_174_)
  );
  \$_OR_  _518_ (
    .A(_174_),
    .B(_135_),
    .Y(_175_)
  );
  \$_AND_  _519_ (
    .A(_175_),
    .B(_136_),
    .Y(_176_)
  );
  \$_OR_  _520_ (
    .A(_176_),
    .B(_121_),
    .Y(fe_pmem_cen)
  );
  \$_INV_  _521_ (
    .A(dbg_mem_en),
    .Y(_177_)
  );
  \$_AND_  _522_ (
    .A(_024_),
    .B(_035_),
    .Y(_178_)
  );
  \$_AND_  _523_ (
    .A(_178_),
    .B(_009_),
    .Y(_179_)
  );
  \$_OR_  _524_ (
    .A(_179_),
    .B(_008_),
    .Y(_180_)
  );
  \$_INV_  _525_ (
    .A(_180_),
    .Y(_181_)
  );
  \$_AND_  _526_ (
    .A(_181_),
    .B(dbg_mem_addr[12]),
    .Y(_182_)
  );
  \$_AND_  _527_ (
    .A(_182_),
    .B(dbg_mem_addr[13]),
    .Y(_183_)
  );
  \$_AND_  _528_ (
    .A(_183_),
    .B(dbg_mem_addr[14]),
    .Y(_184_)
  );
  \$_AND_  _529_ (
    .A(_184_),
    .B(dbg_mem_addr[15]),
    .Y(_185_)
  );
  \$_INV_  _530_ (
    .A(_185_),
    .Y(_186_)
  );
  \$_OR_  _531_ (
    .A(_184_),
    .B(dbg_mem_addr[15]),
    .Y(_187_)
  );
  \$_INV_  _532_ (
    .A(_187_),
    .Y(_188_)
  );
  \$_OR_  _533_ (
    .A(_183_),
    .B(dbg_mem_addr[14]),
    .Y(_189_)
  );
  \$_INV_  _534_ (
    .A(_189_),
    .Y(_190_)
  );
  \$_OR_  _535_ (
    .A(_182_),
    .B(dbg_mem_addr[13]),
    .Y(_191_)
  );
  \$_INV_  _536_ (
    .A(_191_),
    .Y(_192_)
  );
  \$_AND_  _537_ (
    .A(_180_),
    .B(_007_),
    .Y(_193_)
  );
  \$_XOR_  _538_ (
    .A(_179_),
    .B(_008_),
    .Y(_194_)
  );
  \$_AND_  _539_ (
    .A(_194_),
    .B(_179_),
    .Y(_195_)
  );
  \$_INV_  _540_ (
    .A(_195_),
    .Y(_196_)
  );
  \$_OR_  _541_ (
    .A(_196_),
    .B(_193_),
    .Y(_197_)
  );
  \$_OR_  _542_ (
    .A(_197_),
    .B(_192_),
    .Y(_198_)
  );
  \$_OR_  _543_ (
    .A(_198_),
    .B(_190_),
    .Y(_199_)
  );
  \$_OR_  _544_ (
    .A(_199_),
    .B(_184_),
    .Y(_200_)
  );
  \$_OR_  _545_ (
    .A(_200_),
    .B(_188_),
    .Y(_201_)
  );
  \$_OR_  _546_ (
    .A(_201_),
    .B(_185_),
    .Y(_202_)
  );
  \$_AND_  _547_ (
    .A(_202_),
    .B(_186_),
    .Y(_203_)
  );
  \$_OR_  _548_ (
    .A(_203_),
    .B(_177_),
    .Y(_204_)
  );
  \$_OR_  _549_ (
    .A(_082_),
    .B(eu_mab[8]),
    .Y(_205_)
  );
  \$_OR_  _550_ (
    .A(_205_),
    .B(eu_mab[9]),
    .Y(_206_)
  );
  \$_AND_  _551_ (
    .A(_206_),
    .B(eu_mab[10]),
    .Y(_207_)
  );
  \$_AND_  _552_ (
    .A(_207_),
    .B(eu_mab[11]),
    .Y(_208_)
  );
  \$_AND_  _553_ (
    .A(_208_),
    .B(eu_mab[12]),
    .Y(_209_)
  );
  \$_AND_  _554_ (
    .A(_209_),
    .B(eu_mab[13]),
    .Y(_210_)
  );
  \$_AND_  _555_ (
    .A(_210_),
    .B(eu_mab[14]),
    .Y(_211_)
  );
  \$_INV_  _556_ (
    .A(_211_),
    .Y(_212_)
  );
  \$_OR_  _557_ (
    .A(_210_),
    .B(eu_mab[14]),
    .Y(_213_)
  );
  \$_INV_  _558_ (
    .A(_213_),
    .Y(_214_)
  );
  \$_OR_  _559_ (
    .A(_209_),
    .B(eu_mab[13]),
    .Y(_215_)
  );
  \$_INV_  _560_ (
    .A(_215_),
    .Y(_216_)
  );
  \$_OR_  _561_ (
    .A(_208_),
    .B(eu_mab[12]),
    .Y(_217_)
  );
  \$_INV_  _562_ (
    .A(_217_),
    .Y(_218_)
  );
  \$_OR_  _563_ (
    .A(_207_),
    .B(eu_mab[11]),
    .Y(_219_)
  );
  \$_INV_  _564_ (
    .A(_219_),
    .Y(_220_)
  );
  \$_XOR_  _565_ (
    .A(_205_),
    .B(_075_),
    .Y(_221_)
  );
  \$_XOR_  _566_ (
    .A(_206_),
    .B(eu_mab[10]),
    .Y(_222_)
  );
  \$_INV_  _567_ (
    .A(_222_),
    .Y(_223_)
  );
  \$_OR_  _568_ (
    .A(_223_),
    .B(_206_),
    .Y(_224_)
  );
  \$_OR_  _569_ (
    .A(_224_),
    .B(_220_),
    .Y(_225_)
  );
  \$_OR_  _570_ (
    .A(_225_),
    .B(_218_),
    .Y(_226_)
  );
  \$_OR_  _571_ (
    .A(_226_),
    .B(_209_),
    .Y(_227_)
  );
  \$_OR_  _572_ (
    .A(_227_),
    .B(_216_),
    .Y(_228_)
  );
  \$_OR_  _573_ (
    .A(_228_),
    .B(_210_),
    .Y(_229_)
  );
  \$_OR_  _574_ (
    .A(_229_),
    .B(_214_),
    .Y(_230_)
  );
  \$_OR_  _575_ (
    .A(_230_),
    .B(_211_),
    .Y(_231_)
  );
  \$_AND_  _576_ (
    .A(_231_),
    .B(_212_),
    .Y(_232_)
  );
  \$_INV_  _577_ (
    .A(eu_mb_wr[1]),
    .Y(_233_)
  );
  \$_INV_  _578_ (
    .A(eu_mb_wr[0]),
    .Y(_234_)
  );
  \$_AND_  _579_ (
    .A(_234_),
    .B(eu_mb_en),
    .Y(_235_)
  );
  \$_AND_  _580_ (
    .A(_235_),
    .B(_233_),
    .Y(_236_)
  );
  \$_INV_  _581_ (
    .A(_236_),
    .Y(_237_)
  );
  \$_OR_  _582_ (
    .A(_237_),
    .B(_232_),
    .Y(_238_)
  );
  \$_AND_  _583_ (
    .A(_238_),
    .B(fe_pmem_cen),
    .Y(_239_)
  );
  \$_AND_  _584_ (
    .A(_239_),
    .B(_204_),
    .Y(pmem_cen)
  );
  \$_INV_  _585_ (
    .A(_210_),
    .Y(_240_)
  );
  \$_INV_  _586_ (
    .A(_209_),
    .Y(_241_)
  );
  \$_INV_  _587_ (
    .A(_082_),
    .Y(_242_)
  );
  \$_AND_  _588_ (
    .A(_093_),
    .B(_242_),
    .Y(_243_)
  );
  \$_AND_  _589_ (
    .A(_221_),
    .B(_243_),
    .Y(_244_)
  );
  \$_AND_  _590_ (
    .A(_222_),
    .B(_244_),
    .Y(_245_)
  );
  \$_AND_  _591_ (
    .A(_245_),
    .B(_219_),
    .Y(_246_)
  );
  \$_AND_  _592_ (
    .A(_246_),
    .B(_217_),
    .Y(_247_)
  );
  \$_AND_  _593_ (
    .A(_247_),
    .B(_241_),
    .Y(_248_)
  );
  \$_AND_  _594_ (
    .A(_248_),
    .B(_215_),
    .Y(_249_)
  );
  \$_AND_  _595_ (
    .A(_249_),
    .B(_240_),
    .Y(_250_)
  );
  \$_AND_  _596_ (
    .A(_250_),
    .B(_213_),
    .Y(_251_)
  );
  \$_AND_  _597_ (
    .A(_251_),
    .B(_212_),
    .Y(_252_)
  );
  \$_OR_  _598_ (
    .A(_252_),
    .B(_211_),
    .Y(_253_)
  );
  \$_AND_  _599_ (
    .A(_236_),
    .B(_253_),
    .Y(_001_[1])
  );
  \$_INV_  _600_ (
    .A(_134_),
    .Y(_254_)
  );
  \$_INV_  _601_ (
    .A(_133_),
    .Y(_255_)
  );
  \$_OR_  _602_ (
    .A(_164_),
    .B(_143_),
    .Y(_256_)
  );
  \$_OR_  _603_ (
    .A(_131_),
    .B(fe_mab[11]),
    .Y(_257_)
  );
  \$_XOR_  _604_ (
    .A(_130_),
    .B(fe_mab[10]),
    .Y(_258_)
  );
  \$_AND_  _605_ (
    .A(_258_),
    .B(_163_),
    .Y(_259_)
  );
  \$_AND_  _606_ (
    .A(_259_),
    .B(_257_),
    .Y(_260_)
  );
  \$_AND_  _607_ (
    .A(_260_),
    .B(_256_),
    .Y(_261_)
  );
  \$_AND_  _608_ (
    .A(_261_),
    .B(_141_),
    .Y(_262_)
  );
  \$_AND_  _609_ (
    .A(_262_),
    .B(_255_),
    .Y(_263_)
  );
  \$_AND_  _610_ (
    .A(_263_),
    .B(_139_),
    .Y(_264_)
  );
  \$_AND_  _611_ (
    .A(_264_),
    .B(_254_),
    .Y(_265_)
  );
  \$_AND_  _612_ (
    .A(_265_),
    .B(_137_),
    .Y(_266_)
  );
  \$_AND_  _613_ (
    .A(_266_),
    .B(_136_),
    .Y(_267_)
  );
  \$_OR_  _614_ (
    .A(_267_),
    .B(_135_),
    .Y(_268_)
  );
  \$_AND_  _615_ (
    .A(_268_),
    .B(fe_mb_en),
    .Y(_269_)
  );
  \$_AND_  _616_ (
    .A(_001_[1]),
    .B(_269_),
    .Y(fe_pmem_wait)
  );
  \$_AND_  _617_ (
    .A(_009_),
    .B(_035_),
    .Y(_270_)
  );
  \$_AND_  _618_ (
    .A(_270_),
    .B(_008_),
    .Y(_271_)
  );
  \$_AND_  _619_ (
    .A(_271_),
    .B(_007_),
    .Y(_272_)
  );
  \$_AND_  _620_ (
    .A(_272_),
    .B(_006_),
    .Y(_273_)
  );
  \$_AND_  _621_ (
    .A(_273_),
    .B(_005_),
    .Y(_274_)
  );
  \$_OR_  _622_ (
    .A(_274_),
    .B(dbg_mem_addr[15]),
    .Y(_275_)
  );
  \$_AND_  _623_ (
    .A(_275_),
    .B(_066_),
    .Y(dbg_per_en)
  );
  \$_INV_  _624_ (
    .A(dbg_mem_wr[0]),
    .Y(pmem_wen[0])
  );
  \$_AND_  _625_ (
    .A(_234_),
    .B(pmem_wen[0]),
    .Y(dmem_wen[0])
  );
  \$_INV_  _626_ (
    .A(dbg_mem_wr[1]),
    .Y(pmem_wen[1])
  );
  \$_AND_  _627_ (
    .A(_233_),
    .B(pmem_wen[1]),
    .Y(dmem_wen[1])
  );
  \$_INV_  _628_ (
    .A(_184_),
    .Y(_276_)
  );
  \$_INV_  _629_ (
    .A(_193_),
    .Y(_277_)
  );
  \$_AND_  _630_ (
    .A(_195_),
    .B(_277_),
    .Y(_278_)
  );
  \$_AND_  _631_ (
    .A(_278_),
    .B(_191_),
    .Y(_279_)
  );
  \$_AND_  _632_ (
    .A(_279_),
    .B(_189_),
    .Y(_280_)
  );
  \$_AND_  _633_ (
    .A(_280_),
    .B(_276_),
    .Y(_281_)
  );
  \$_AND_  _634_ (
    .A(_281_),
    .B(_187_),
    .Y(_282_)
  );
  \$_AND_  _635_ (
    .A(_282_),
    .B(_186_),
    .Y(_283_)
  );
  \$_OR_  _636_ (
    .A(_283_),
    .B(_185_),
    .Y(_284_)
  );
  \$_AND_  _637_ (
    .A(_284_),
    .B(dbg_mem_en),
    .Y(_000_[1])
  );
  \$_INV_  _638_ (
    .A(fe_pmem_cen_dly),
    .Y(_285_)
  );
  \$_INV_  _639_ (
    .A(dbg_halt_st),
    .Y(_286_)
  );
  \$_AND_  _640_ (
    .A(_286_),
    .B(_285_),
    .Y(_287_)
  );
  \$_INV_  _641_ (
    .A(_287_),
    .Y(_288_)
  );
  \$_OR_  _642_ (
    .A(_288_),
    .B(_269_),
    .Y(_289_)
  );
  \$_MUX_  _643_ (
    .A(pmem_dout[0]),
    .B(pmem_dout_bckup[0]),
    .S(_289_),
    .Y(_002_[0])
  );
  \$_MUX_  _644_ (
    .A(pmem_dout[10]),
    .B(pmem_dout_bckup[10]),
    .S(_289_),
    .Y(_002_[10])
  );
  \$_MUX_  _645_ (
    .A(pmem_dout[11]),
    .B(pmem_dout_bckup[11]),
    .S(_289_),
    .Y(_002_[11])
  );
  \$_MUX_  _646_ (
    .A(pmem_dout[12]),
    .B(pmem_dout_bckup[12]),
    .S(_289_),
    .Y(_002_[12])
  );
  \$_MUX_  _647_ (
    .A(pmem_dout[13]),
    .B(pmem_dout_bckup[13]),
    .S(_289_),
    .Y(_002_[13])
  );
  \$_MUX_  _648_ (
    .A(pmem_dout[14]),
    .B(pmem_dout_bckup[14]),
    .S(_289_),
    .Y(_002_[14])
  );
  \$_MUX_  _649_ (
    .A(pmem_dout[15]),
    .B(pmem_dout_bckup[15]),
    .S(_289_),
    .Y(_002_[15])
  );
  \$_MUX_  _650_ (
    .A(pmem_dout[1]),
    .B(pmem_dout_bckup[1]),
    .S(_289_),
    .Y(_002_[1])
  );
  \$_MUX_  _651_ (
    .A(pmem_dout[2]),
    .B(pmem_dout_bckup[2]),
    .S(_289_),
    .Y(_002_[2])
  );
  \$_MUX_  _652_ (
    .A(pmem_dout[3]),
    .B(pmem_dout_bckup[3]),
    .S(_289_),
    .Y(_002_[3])
  );
  \$_MUX_  _653_ (
    .A(pmem_dout[4]),
    .B(pmem_dout_bckup[4]),
    .S(_289_),
    .Y(_002_[4])
  );
  \$_MUX_  _654_ (
    .A(pmem_dout[5]),
    .B(pmem_dout_bckup[5]),
    .S(_289_),
    .Y(_002_[5])
  );
  \$_MUX_  _655_ (
    .A(pmem_dout[6]),
    .B(pmem_dout_bckup[6]),
    .S(_289_),
    .Y(_002_[6])
  );
  \$_MUX_  _656_ (
    .A(pmem_dout[7]),
    .B(pmem_dout_bckup[7]),
    .S(_289_),
    .Y(_002_[7])
  );
  \$_MUX_  _657_ (
    .A(pmem_dout[8]),
    .B(pmem_dout_bckup[8]),
    .S(_289_),
    .Y(_002_[8])
  );
  \$_MUX_  _658_ (
    .A(pmem_dout[9]),
    .B(pmem_dout_bckup[9]),
    .S(_289_),
    .Y(_002_[9])
  );
  \$_INV_  _659_ (
    .A(_289_),
    .Y(_290_)
  );
  \$_OR_  _660_ (
    .A(fe_pmem_cen),
    .B(_285_),
    .Y(_291_)
  );
  \$_AND_  _661_ (
    .A(pmem_dout_bckup_sel),
    .B(_286_),
    .Y(_292_)
  );
  \$_AND_  _662_ (
    .A(_292_),
    .B(_289_),
    .Y(_293_)
  );
  \$_AND_  _663_ (
    .A(_293_),
    .B(_291_),
    .Y(_294_)
  );
  \$_OR_  _664_ (
    .A(_294_),
    .B(_290_),
    .Y(_003_)
  );
  \$_MUX_  _665_ (
    .A(dbg_mem_addr[1]),
    .B(eu_mab[0]),
    .S(_069_),
    .Y(dmem_addr[0])
  );
  \$_MUX_  _666_ (
    .A(dbg_mem_addr[2]),
    .B(eu_mab[1]),
    .S(_069_),
    .Y(dmem_addr[1])
  );
  \$_MUX_  _667_ (
    .A(dbg_mem_addr[3]),
    .B(eu_mab[2]),
    .S(_069_),
    .Y(dmem_addr[2])
  );
  \$_MUX_  _668_ (
    .A(dbg_mem_addr[4]),
    .B(eu_mab[3]),
    .S(_069_),
    .Y(dmem_addr[3])
  );
  \$_MUX_  _669_ (
    .A(dbg_mem_addr[5]),
    .B(eu_mab[4]),
    .S(_069_),
    .Y(dmem_addr[4])
  );
  \$_MUX_  _670_ (
    .A(dbg_mem_addr[6]),
    .B(eu_mab[5]),
    .S(_069_),
    .Y(dmem_addr[5])
  );
  \$_MUX_  _671_ (
    .A(dbg_mem_dout[0]),
    .B(eu_mdb_out[0]),
    .S(_069_),
    .Y(dmem_din[0])
  );
  \$_MUX_  _672_ (
    .A(dbg_mem_dout[10]),
    .B(eu_mdb_out[10]),
    .S(_069_),
    .Y(dmem_din[10])
  );
  \$_MUX_  _673_ (
    .A(dbg_mem_dout[11]),
    .B(eu_mdb_out[11]),
    .S(_069_),
    .Y(dmem_din[11])
  );
  \$_MUX_  _674_ (
    .A(dbg_mem_dout[12]),
    .B(eu_mdb_out[12]),
    .S(_069_),
    .Y(dmem_din[12])
  );
  \$_MUX_  _675_ (
    .A(dbg_mem_dout[13]),
    .B(eu_mdb_out[13]),
    .S(_069_),
    .Y(dmem_din[13])
  );
  \$_MUX_  _676_ (
    .A(dbg_mem_dout[14]),
    .B(eu_mdb_out[14]),
    .S(_069_),
    .Y(dmem_din[14])
  );
  \$_MUX_  _677_ (
    .A(dbg_mem_dout[15]),
    .B(eu_mdb_out[15]),
    .S(_069_),
    .Y(dmem_din[15])
  );
  \$_MUX_  _678_ (
    .A(dbg_mem_dout[1]),
    .B(eu_mdb_out[1]),
    .S(_069_),
    .Y(dmem_din[1])
  );
  \$_MUX_  _679_ (
    .A(dbg_mem_dout[2]),
    .B(eu_mdb_out[2]),
    .S(_069_),
    .Y(dmem_din[2])
  );
  \$_MUX_  _680_ (
    .A(dbg_mem_dout[3]),
    .B(eu_mdb_out[3]),
    .S(_069_),
    .Y(dmem_din[3])
  );
  \$_MUX_  _681_ (
    .A(dbg_mem_dout[4]),
    .B(eu_mdb_out[4]),
    .S(_069_),
    .Y(dmem_din[4])
  );
  \$_MUX_  _682_ (
    .A(dbg_mem_dout[5]),
    .B(eu_mdb_out[5]),
    .S(_069_),
    .Y(dmem_din[5])
  );
  \$_MUX_  _683_ (
    .A(dbg_mem_dout[6]),
    .B(eu_mdb_out[6]),
    .S(_069_),
    .Y(dmem_din[6])
  );
  \$_MUX_  _684_ (
    .A(dbg_mem_dout[7]),
    .B(eu_mdb_out[7]),
    .S(_069_),
    .Y(dmem_din[7])
  );
  \$_MUX_  _685_ (
    .A(dbg_mem_dout[8]),
    .B(eu_mdb_out[8]),
    .S(_069_),
    .Y(dmem_din[8])
  );
  \$_MUX_  _686_ (
    .A(dbg_mem_dout[9]),
    .B(eu_mdb_out[9]),
    .S(_069_),
    .Y(dmem_din[9])
  );
  \$_MUX_  _687_ (
    .A(fe_mab[0]),
    .B(eu_mab[0]),
    .S(_001_[1]),
    .Y(_295_)
  );
  \$_MUX_  _688_ (
    .A(_295_),
    .B(dbg_mem_addr[1]),
    .S(_000_[1]),
    .Y(pmem_addr[0])
  );
  \$_MUX_  _689_ (
    .A(fe_mab[1]),
    .B(eu_mab[1]),
    .S(_001_[1]),
    .Y(_296_)
  );
  \$_MUX_  _690_ (
    .A(_296_),
    .B(dbg_mem_addr[2]),
    .S(_000_[1]),
    .Y(pmem_addr[1])
  );
  \$_MUX_  _691_ (
    .A(fe_mab[2]),
    .B(eu_mab[2]),
    .S(_001_[1]),
    .Y(_297_)
  );
  \$_MUX_  _692_ (
    .A(_297_),
    .B(dbg_mem_addr[3]),
    .S(_000_[1]),
    .Y(pmem_addr[2])
  );
  \$_MUX_  _693_ (
    .A(fe_mab[3]),
    .B(eu_mab[3]),
    .S(_001_[1]),
    .Y(_298_)
  );
  \$_MUX_  _694_ (
    .A(_298_),
    .B(dbg_mem_addr[4]),
    .S(_000_[1]),
    .Y(pmem_addr[3])
  );
  \$_MUX_  _695_ (
    .A(fe_mab[4]),
    .B(eu_mab[4]),
    .S(_001_[1]),
    .Y(_299_)
  );
  \$_MUX_  _696_ (
    .A(_299_),
    .B(dbg_mem_addr[5]),
    .S(_000_[1]),
    .Y(pmem_addr[4])
  );
  \$_MUX_  _697_ (
    .A(fe_mab[5]),
    .B(eu_mab[5]),
    .S(_001_[1]),
    .Y(_300_)
  );
  \$_MUX_  _698_ (
    .A(_300_),
    .B(dbg_mem_addr[6]),
    .S(_000_[1]),
    .Y(pmem_addr[5])
  );
  \$_MUX_  _699_ (
    .A(fe_mab[6]),
    .B(eu_mab[6]),
    .S(_001_[1]),
    .Y(_301_)
  );
  \$_MUX_  _700_ (
    .A(_301_),
    .B(dbg_mem_addr[7]),
    .S(_000_[1]),
    .Y(pmem_addr[6])
  );
  \$_MUX_  _701_ (
    .A(fe_mab[7]),
    .B(eu_mab[7]),
    .S(_001_[1]),
    .Y(_302_)
  );
  \$_MUX_  _702_ (
    .A(_302_),
    .B(dbg_mem_addr[8]),
    .S(_000_[1]),
    .Y(pmem_addr[7])
  );
  \$_MUX_  _703_ (
    .A(fe_mab[8]),
    .B(eu_mab[8]),
    .S(_001_[1]),
    .Y(_303_)
  );
  \$_MUX_  _704_ (
    .A(_303_),
    .B(dbg_mem_addr[9]),
    .S(_000_[1]),
    .Y(pmem_addr[8])
  );
  \$_MUX_  _705_ (
    .A(fe_mab[9]),
    .B(eu_mab[9]),
    .S(_001_[1]),
    .Y(_304_)
  );
  \$_MUX_  _706_ (
    .A(_304_),
    .B(dbg_mem_addr[10]),
    .S(_000_[1]),
    .Y(pmem_addr[9])
  );
  \$_MUX_  _707_ (
    .A(eu_mdb_out[0]),
    .B(dbg_mem_dout[0]),
    .S(dbg_mem_en),
    .Y(per_din[0])
  );
  \$_MUX_  _708_ (
    .A(eu_mdb_out[10]),
    .B(dbg_mem_dout[10]),
    .S(dbg_mem_en),
    .Y(per_din[10])
  );
  \$_MUX_  _709_ (
    .A(eu_mdb_out[11]),
    .B(dbg_mem_dout[11]),
    .S(dbg_mem_en),
    .Y(per_din[11])
  );
  \$_MUX_  _710_ (
    .A(eu_mdb_out[12]),
    .B(dbg_mem_dout[12]),
    .S(dbg_mem_en),
    .Y(per_din[12])
  );
  \$_MUX_  _711_ (
    .A(eu_mdb_out[13]),
    .B(dbg_mem_dout[13]),
    .S(dbg_mem_en),
    .Y(per_din[13])
  );
  \$_MUX_  _712_ (
    .A(eu_mdb_out[14]),
    .B(dbg_mem_dout[14]),
    .S(dbg_mem_en),
    .Y(per_din[14])
  );
  \$_MUX_  _713_ (
    .A(eu_mdb_out[15]),
    .B(dbg_mem_dout[15]),
    .S(dbg_mem_en),
    .Y(per_din[15])
  );
  \$_MUX_  _714_ (
    .A(eu_mdb_out[1]),
    .B(dbg_mem_dout[1]),
    .S(dbg_mem_en),
    .Y(per_din[1])
  );
  \$_MUX_  _715_ (
    .A(eu_mdb_out[2]),
    .B(dbg_mem_dout[2]),
    .S(dbg_mem_en),
    .Y(per_din[2])
  );
  \$_MUX_  _716_ (
    .A(eu_mdb_out[3]),
    .B(dbg_mem_dout[3]),
    .S(dbg_mem_en),
    .Y(per_din[3])
  );
  \$_MUX_  _717_ (
    .A(eu_mdb_out[4]),
    .B(dbg_mem_dout[4]),
    .S(dbg_mem_en),
    .Y(per_din[4])
  );
  \$_MUX_  _718_ (
    .A(eu_mdb_out[5]),
    .B(dbg_mem_dout[5]),
    .S(dbg_mem_en),
    .Y(per_din[5])
  );
  \$_MUX_  _719_ (
    .A(eu_mdb_out[6]),
    .B(dbg_mem_dout[6]),
    .S(dbg_mem_en),
    .Y(per_din[6])
  );
  \$_MUX_  _720_ (
    .A(eu_mdb_out[7]),
    .B(dbg_mem_dout[7]),
    .S(dbg_mem_en),
    .Y(per_din[7])
  );
  \$_MUX_  _721_ (
    .A(eu_mdb_out[8]),
    .B(dbg_mem_dout[8]),
    .S(dbg_mem_en),
    .Y(per_din[8])
  );
  \$_MUX_  _722_ (
    .A(eu_mdb_out[9]),
    .B(dbg_mem_dout[9]),
    .S(dbg_mem_en),
    .Y(per_din[9])
  );
  \$_MUX_  _723_ (
    .A(eu_mb_wr[0]),
    .B(dbg_mem_wr[0]),
    .S(dbg_mem_en),
    .Y(per_we[0])
  );
  \$_MUX_  _724_ (
    .A(eu_mb_wr[1]),
    .B(dbg_mem_wr[1]),
    .S(dbg_mem_en),
    .Y(per_we[1])
  );
  \$_AND_  _725_ (
    .A(dbg_per_en),
    .B(dbg_mem_en),
    .Y(_305_)
  );
  \$_AND_  _726_ (
    .A(_075_),
    .B(_092_),
    .Y(_306_)
  );
  \$_AND_  _727_ (
    .A(_306_),
    .B(_074_),
    .Y(_307_)
  );
  \$_AND_  _728_ (
    .A(_307_),
    .B(_073_),
    .Y(_308_)
  );
  \$_AND_  _729_ (
    .A(_308_),
    .B(_072_),
    .Y(_309_)
  );
  \$_AND_  _730_ (
    .A(_309_),
    .B(_071_),
    .Y(_310_)
  );
  \$_OR_  _731_ (
    .A(_310_),
    .B(eu_mab[14]),
    .Y(_311_)
  );
  \$_AND_  _732_ (
    .A(_117_),
    .B(_177_),
    .Y(_312_)
  );
  \$_AND_  _733_ (
    .A(_312_),
    .B(_311_),
    .Y(_313_)
  );
  \$_OR_  _734_ (
    .A(_313_),
    .B(_305_),
    .Y(per_en)
  );
  \$_MUX_  _735_ (
    .A(eu_mab[0]),
    .B(dbg_mem_addr[1]),
    .S(dbg_mem_en),
    .Y(per_addr[0])
  );
  \$_MUX_  _736_ (
    .A(eu_mab[1]),
    .B(dbg_mem_addr[2]),
    .S(dbg_mem_en),
    .Y(per_addr[1])
  );
  \$_MUX_  _737_ (
    .A(eu_mab[2]),
    .B(dbg_mem_addr[3]),
    .S(dbg_mem_en),
    .Y(per_addr[2])
  );
  \$_MUX_  _738_ (
    .A(eu_mab[3]),
    .B(dbg_mem_addr[4]),
    .S(dbg_mem_en),
    .Y(per_addr[3])
  );
  \$_MUX_  _739_ (
    .A(eu_mab[4]),
    .B(dbg_mem_addr[5]),
    .S(dbg_mem_en),
    .Y(per_addr[4])
  );
  \$_MUX_  _740_ (
    .A(eu_mab[5]),
    .B(dbg_mem_addr[6]),
    .S(dbg_mem_en),
    .Y(per_addr[5])
  );
  \$_MUX_  _741_ (
    .A(eu_mab[6]),
    .B(dbg_mem_addr[7]),
    .S(dbg_mem_en),
    .Y(per_addr[6])
  );
  \$_MUX_  _742_ (
    .A(eu_mab[7]),
    .B(dbg_mem_addr[8]),
    .S(dbg_mem_en),
    .Y(per_addr[7])
  );
  \$_MUX_  _743_ (
    .A(pmem_dout[0]),
    .B(pmem_dout_bckup[0]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[0])
  );
  \$_MUX_  _744_ (
    .A(pmem_dout[10]),
    .B(pmem_dout_bckup[10]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[10])
  );
  \$_MUX_  _745_ (
    .A(pmem_dout[11]),
    .B(pmem_dout_bckup[11]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[11])
  );
  \$_MUX_  _746_ (
    .A(pmem_dout[12]),
    .B(pmem_dout_bckup[12]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[12])
  );
  \$_MUX_  _747_ (
    .A(pmem_dout[13]),
    .B(pmem_dout_bckup[13]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[13])
  );
  \$_MUX_  _748_ (
    .A(pmem_dout[14]),
    .B(pmem_dout_bckup[14]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[14])
  );
  \$_MUX_  _749_ (
    .A(pmem_dout[15]),
    .B(pmem_dout_bckup[15]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[15])
  );
  \$_MUX_  _750_ (
    .A(pmem_dout[1]),
    .B(pmem_dout_bckup[1]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[1])
  );
  \$_MUX_  _751_ (
    .A(pmem_dout[2]),
    .B(pmem_dout_bckup[2]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[2])
  );
  \$_MUX_  _752_ (
    .A(pmem_dout[3]),
    .B(pmem_dout_bckup[3]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[3])
  );
  \$_MUX_  _753_ (
    .A(pmem_dout[4]),
    .B(pmem_dout_bckup[4]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[4])
  );
  \$_MUX_  _754_ (
    .A(pmem_dout[5]),
    .B(pmem_dout_bckup[5]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[5])
  );
  \$_MUX_  _755_ (
    .A(pmem_dout[6]),
    .B(pmem_dout_bckup[6]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[6])
  );
  \$_MUX_  _756_ (
    .A(pmem_dout[7]),
    .B(pmem_dout_bckup[7]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[7])
  );
  \$_MUX_  _757_ (
    .A(pmem_dout[8]),
    .B(pmem_dout_bckup[8]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[8])
  );
  \$_MUX_  _758_ (
    .A(pmem_dout[9]),
    .B(pmem_dout_bckup[9]),
    .S(pmem_dout_bckup_sel),
    .Y(fe_mdb_in[9])
  );
  \$_MUX_  _759_ (
    .A(dmem_dout[0]),
    .B(per_dout_val[0]),
    .S(eu_mdb_in_sel[0]),
    .Y(_314_)
  );
  \$_MUX_  _760_ (
    .A(_314_),
    .B(pmem_dout[0]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[0])
  );
  \$_MUX_  _761_ (
    .A(dmem_dout[10]),
    .B(per_dout_val[10]),
    .S(eu_mdb_in_sel[0]),
    .Y(_315_)
  );
  \$_MUX_  _762_ (
    .A(_315_),
    .B(pmem_dout[10]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[10])
  );
  \$_MUX_  _763_ (
    .A(dmem_dout[11]),
    .B(per_dout_val[11]),
    .S(eu_mdb_in_sel[0]),
    .Y(_316_)
  );
  \$_MUX_  _764_ (
    .A(_316_),
    .B(pmem_dout[11]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[11])
  );
  \$_MUX_  _765_ (
    .A(dmem_dout[12]),
    .B(per_dout_val[12]),
    .S(eu_mdb_in_sel[0]),
    .Y(_317_)
  );
  \$_MUX_  _766_ (
    .A(_317_),
    .B(pmem_dout[12]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[12])
  );
  \$_MUX_  _767_ (
    .A(dmem_dout[13]),
    .B(per_dout_val[13]),
    .S(eu_mdb_in_sel[0]),
    .Y(_318_)
  );
  \$_MUX_  _768_ (
    .A(_318_),
    .B(pmem_dout[13]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[13])
  );
  \$_MUX_  _769_ (
    .A(dmem_dout[14]),
    .B(per_dout_val[14]),
    .S(eu_mdb_in_sel[0]),
    .Y(_319_)
  );
  \$_MUX_  _770_ (
    .A(_319_),
    .B(pmem_dout[14]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[14])
  );
  \$_MUX_  _771_ (
    .A(dmem_dout[15]),
    .B(per_dout_val[15]),
    .S(eu_mdb_in_sel[0]),
    .Y(_320_)
  );
  \$_MUX_  _772_ (
    .A(_320_),
    .B(pmem_dout[15]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[15])
  );
  \$_MUX_  _773_ (
    .A(dmem_dout[1]),
    .B(per_dout_val[1]),
    .S(eu_mdb_in_sel[0]),
    .Y(_321_)
  );
  \$_MUX_  _774_ (
    .A(_321_),
    .B(pmem_dout[1]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[1])
  );
  \$_MUX_  _775_ (
    .A(dmem_dout[2]),
    .B(per_dout_val[2]),
    .S(eu_mdb_in_sel[0]),
    .Y(_322_)
  );
  \$_MUX_  _776_ (
    .A(_322_),
    .B(pmem_dout[2]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[2])
  );
  \$_MUX_  _777_ (
    .A(dmem_dout[3]),
    .B(per_dout_val[3]),
    .S(eu_mdb_in_sel[0]),
    .Y(_323_)
  );
  \$_MUX_  _778_ (
    .A(_323_),
    .B(pmem_dout[3]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[3])
  );
  \$_MUX_  _779_ (
    .A(dmem_dout[4]),
    .B(per_dout_val[4]),
    .S(eu_mdb_in_sel[0]),
    .Y(_324_)
  );
  \$_MUX_  _780_ (
    .A(_324_),
    .B(pmem_dout[4]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[4])
  );
  \$_MUX_  _781_ (
    .A(dmem_dout[5]),
    .B(per_dout_val[5]),
    .S(eu_mdb_in_sel[0]),
    .Y(_325_)
  );
  \$_MUX_  _782_ (
    .A(_325_),
    .B(pmem_dout[5]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[5])
  );
  \$_MUX_  _783_ (
    .A(dmem_dout[6]),
    .B(per_dout_val[6]),
    .S(eu_mdb_in_sel[0]),
    .Y(_326_)
  );
  \$_MUX_  _784_ (
    .A(_326_),
    .B(pmem_dout[6]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[6])
  );
  \$_MUX_  _785_ (
    .A(dmem_dout[7]),
    .B(per_dout_val[7]),
    .S(eu_mdb_in_sel[0]),
    .Y(_327_)
  );
  \$_MUX_  _786_ (
    .A(_327_),
    .B(pmem_dout[7]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[7])
  );
  \$_MUX_  _787_ (
    .A(dmem_dout[8]),
    .B(per_dout_val[8]),
    .S(eu_mdb_in_sel[0]),
    .Y(_328_)
  );
  \$_MUX_  _788_ (
    .A(_328_),
    .B(pmem_dout[8]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[8])
  );
  \$_MUX_  _789_ (
    .A(dmem_dout[9]),
    .B(per_dout_val[9]),
    .S(eu_mdb_in_sel[0]),
    .Y(_329_)
  );
  \$_MUX_  _790_ (
    .A(_329_),
    .B(pmem_dout[9]),
    .S(eu_mdb_in_sel[1]),
    .Y(eu_mdb_in[9])
  );
  \$_MUX_  _791_ (
    .A(dmem_dout[0]),
    .B(per_dout_val[0]),
    .S(dbg_mem_din_sel[0]),
    .Y(_330_)
  );
  \$_MUX_  _792_ (
    .A(_330_),
    .B(pmem_dout[0]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[0])
  );
  \$_MUX_  _793_ (
    .A(dmem_dout[10]),
    .B(per_dout_val[10]),
    .S(dbg_mem_din_sel[0]),
    .Y(_331_)
  );
  \$_MUX_  _794_ (
    .A(_331_),
    .B(pmem_dout[10]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[10])
  );
  \$_MUX_  _795_ (
    .A(dmem_dout[11]),
    .B(per_dout_val[11]),
    .S(dbg_mem_din_sel[0]),
    .Y(_332_)
  );
  \$_MUX_  _796_ (
    .A(_332_),
    .B(pmem_dout[11]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[11])
  );
  \$_MUX_  _797_ (
    .A(dmem_dout[12]),
    .B(per_dout_val[12]),
    .S(dbg_mem_din_sel[0]),
    .Y(_333_)
  );
  \$_MUX_  _798_ (
    .A(_333_),
    .B(pmem_dout[12]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[12])
  );
  \$_MUX_  _799_ (
    .A(dmem_dout[13]),
    .B(per_dout_val[13]),
    .S(dbg_mem_din_sel[0]),
    .Y(_334_)
  );
  \$_MUX_  _800_ (
    .A(_334_),
    .B(pmem_dout[13]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[13])
  );
  \$_MUX_  _801_ (
    .A(dmem_dout[14]),
    .B(per_dout_val[14]),
    .S(dbg_mem_din_sel[0]),
    .Y(_335_)
  );
  \$_MUX_  _802_ (
    .A(_335_),
    .B(pmem_dout[14]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[14])
  );
  \$_MUX_  _803_ (
    .A(dmem_dout[15]),
    .B(per_dout_val[15]),
    .S(dbg_mem_din_sel[0]),
    .Y(_336_)
  );
  \$_MUX_  _804_ (
    .A(_336_),
    .B(pmem_dout[15]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[15])
  );
  \$_MUX_  _805_ (
    .A(dmem_dout[1]),
    .B(per_dout_val[1]),
    .S(dbg_mem_din_sel[0]),
    .Y(_337_)
  );
  \$_MUX_  _806_ (
    .A(_337_),
    .B(pmem_dout[1]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[1])
  );
  \$_MUX_  _807_ (
    .A(dmem_dout[2]),
    .B(per_dout_val[2]),
    .S(dbg_mem_din_sel[0]),
    .Y(_338_)
  );
  \$_MUX_  _808_ (
    .A(_338_),
    .B(pmem_dout[2]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[2])
  );
  \$_MUX_  _809_ (
    .A(dmem_dout[3]),
    .B(per_dout_val[3]),
    .S(dbg_mem_din_sel[0]),
    .Y(_339_)
  );
  \$_MUX_  _810_ (
    .A(_339_),
    .B(pmem_dout[3]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[3])
  );
  \$_MUX_  _811_ (
    .A(dmem_dout[4]),
    .B(per_dout_val[4]),
    .S(dbg_mem_din_sel[0]),
    .Y(_340_)
  );
  \$_MUX_  _812_ (
    .A(_340_),
    .B(pmem_dout[4]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[4])
  );
  \$_MUX_  _813_ (
    .A(dmem_dout[5]),
    .B(per_dout_val[5]),
    .S(dbg_mem_din_sel[0]),
    .Y(_341_)
  );
  \$_MUX_  _814_ (
    .A(_341_),
    .B(pmem_dout[5]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[5])
  );
  \$_MUX_  _815_ (
    .A(dmem_dout[6]),
    .B(per_dout_val[6]),
    .S(dbg_mem_din_sel[0]),
    .Y(_342_)
  );
  \$_MUX_  _816_ (
    .A(_342_),
    .B(pmem_dout[6]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[6])
  );
  \$_MUX_  _817_ (
    .A(dmem_dout[7]),
    .B(per_dout_val[7]),
    .S(dbg_mem_din_sel[0]),
    .Y(_343_)
  );
  \$_MUX_  _818_ (
    .A(_343_),
    .B(pmem_dout[7]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[7])
  );
  \$_MUX_  _819_ (
    .A(dmem_dout[8]),
    .B(per_dout_val[8]),
    .S(dbg_mem_din_sel[0]),
    .Y(_344_)
  );
  \$_MUX_  _820_ (
    .A(_344_),
    .B(pmem_dout[8]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[8])
  );
  \$_MUX_  _821_ (
    .A(dmem_dout[9]),
    .B(per_dout_val[9]),
    .S(dbg_mem_din_sel[0]),
    .Y(_345_)
  );
  \$_MUX_  _822_ (
    .A(_345_),
    .B(pmem_dout[9]),
    .S(dbg_mem_din_sel[1]),
    .Y(dbg_mem_din[9])
  );
  \$_DFF_PP0_  \per_dout_val_reg[0]  /* _823_ */ (
    .C(mclk),
    .D(per_dout[0]),
    .Q(per_dout_val[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[10]  /* _824_ */ (
    .C(mclk),
    .D(per_dout[10]),
    .Q(per_dout_val[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[11]  /* _825_ */ (
    .C(mclk),
    .D(per_dout[11]),
    .Q(per_dout_val[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[12]  /* _826_ */ (
    .C(mclk),
    .D(per_dout[12]),
    .Q(per_dout_val[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[13]  /* _827_ */ (
    .C(mclk),
    .D(per_dout[13]),
    .Q(per_dout_val[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[14]  /* _828_ */ (
    .C(mclk),
    .D(per_dout[14]),
    .Q(per_dout_val[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[15]  /* _829_ */ (
    .C(mclk),
    .D(per_dout[15]),
    .Q(per_dout_val[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[1]  /* _830_ */ (
    .C(mclk),
    .D(per_dout[1]),
    .Q(per_dout_val[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[2]  /* _831_ */ (
    .C(mclk),
    .D(per_dout[2]),
    .Q(per_dout_val[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[3]  /* _832_ */ (
    .C(mclk),
    .D(per_dout[3]),
    .Q(per_dout_val[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[4]  /* _833_ */ (
    .C(mclk),
    .D(per_dout[4]),
    .Q(per_dout_val[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[5]  /* _834_ */ (
    .C(mclk),
    .D(per_dout[5]),
    .Q(per_dout_val[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[6]  /* _835_ */ (
    .C(mclk),
    .D(per_dout[6]),
    .Q(per_dout_val[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[7]  /* _836_ */ (
    .C(mclk),
    .D(per_dout[7]),
    .Q(per_dout_val[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[8]  /* _837_ */ (
    .C(mclk),
    .D(per_dout[8]),
    .Q(per_dout_val[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \per_dout_val_reg[9]  /* _838_ */ (
    .C(mclk),
    .D(per_dout[9]),
    .Q(per_dout_val[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  fe_pmem_cen_dly_reg /* _839_ */ (
    .C(mclk),
    .D(fe_pmem_cen),
    .Q(fe_pmem_cen_dly),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[0]  /* _840_ */ (
    .C(mclk),
    .D(_002_[0]),
    .Q(pmem_dout_bckup[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[10]  /* _841_ */ (
    .C(mclk),
    .D(_002_[10]),
    .Q(pmem_dout_bckup[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[11]  /* _842_ */ (
    .C(mclk),
    .D(_002_[11]),
    .Q(pmem_dout_bckup[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[12]  /* _843_ */ (
    .C(mclk),
    .D(_002_[12]),
    .Q(pmem_dout_bckup[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[13]  /* _844_ */ (
    .C(mclk),
    .D(_002_[13]),
    .Q(pmem_dout_bckup[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[14]  /* _845_ */ (
    .C(mclk),
    .D(_002_[14]),
    .Q(pmem_dout_bckup[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[15]  /* _846_ */ (
    .C(mclk),
    .D(_002_[15]),
    .Q(pmem_dout_bckup[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[1]  /* _847_ */ (
    .C(mclk),
    .D(_002_[1]),
    .Q(pmem_dout_bckup[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[2]  /* _848_ */ (
    .C(mclk),
    .D(_002_[2]),
    .Q(pmem_dout_bckup[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[3]  /* _849_ */ (
    .C(mclk),
    .D(_002_[3]),
    .Q(pmem_dout_bckup[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[4]  /* _850_ */ (
    .C(mclk),
    .D(_002_[4]),
    .Q(pmem_dout_bckup[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[5]  /* _851_ */ (
    .C(mclk),
    .D(_002_[5]),
    .Q(pmem_dout_bckup[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[6]  /* _852_ */ (
    .C(mclk),
    .D(_002_[6]),
    .Q(pmem_dout_bckup[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[7]  /* _853_ */ (
    .C(mclk),
    .D(_002_[7]),
    .Q(pmem_dout_bckup[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[8]  /* _854_ */ (
    .C(mclk),
    .D(_002_[8]),
    .Q(pmem_dout_bckup[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \pmem_dout_bckup_reg[9]  /* _855_ */ (
    .C(mclk),
    .D(_002_[9]),
    .Q(pmem_dout_bckup[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  pmem_dout_bckup_sel_reg /* _856_ */ (
    .C(mclk),
    .D(_003_),
    .Q(pmem_dout_bckup_sel),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \eu_mdb_in_sel_reg[0]  /* _857_ */ (
    .C(mclk),
    .D(per_en),
    .Q(eu_mdb_in_sel[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \eu_mdb_in_sel_reg[1]  /* _858_ */ (
    .C(mclk),
    .D(_001_[1]),
    .Q(eu_mdb_in_sel[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \dbg_mem_din_sel_reg[0]  /* _859_ */ (
    .C(mclk),
    .D(dbg_per_en),
    .Q(dbg_mem_din_sel[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \dbg_mem_din_sel_reg[1]  /* _860_ */ (
    .C(mclk),
    .D(_000_[1]),
    .Q(dbg_mem_din_sel[1]),
    .R(puc_rst)
  );
  assign mclk_bckup = mclk;
  assign per_addr[13:8] = 6'b000000;
  assign per_addr_ful = { 7'b0000000, per_addr[7:0] };
  assign per_addr_mux = per_addr[7:0];
  assign pmem_din = dbg_mem_dout;
endmodule

module omsp_multiplier(per_dout, mclk, per_addr, per_din, per_en, per_we, puc_rst, scan_enable);
  wire _0000_;
  wire [15:0] _0001_;
  wire [15:0] _0002_;
  wire [15:0] _0003_;
  wire [15:0] _0004_;
  wire _0005_;
  wire [1:0] _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire acc_sel;
  wire [1:0] cycle;
  wire early_read;
  input mclk;
  wire mclk_op1;
  wire mclk_op2;
  wire mclk_reshi;
  wire mclk_reslo;
  wire [15:0] op1;
  wire [15:0] op1_rd;
  wire [16:0] op1_xp;
  wire [15:0] op2;
  wire [8:0] op2_hi_xp;
  wire [8:0] op2_lo_xp;
  wire [15:0] op2_rd;
  wire op2_wr;
  wire [8:0] op2_xp;
  input [13:0] per_addr;
  input [15:0] per_din;
  output [15:0] per_dout;
  input per_en;
  input [1:0] per_we;
  wire [25:0] product;
  input puc_rst;
  wire [3:0] reg_addr;
  wire [15:0] reg_wr;
  wire [15:0] reshi;
  wire [15:0] reslo;
  wire [31:0] result;
  input scan_enable;
  wire sign_sel;
  wire [15:0] sumext;
  wire [1:0] sumext_s;
  \$_INV_  _0572_ (
    .A(per_addr[0]),
    .Y(_0007_)
  );
  \$_INV_  _0573_ (
    .A(per_addr[1]),
    .Y(_0008_)
  );
  \$_AND_  _0574_ (
    .A(_0008_),
    .B(_0007_),
    .Y(_0009_)
  );
  \$_AND_  _0575_ (
    .A(_0009_),
    .B(per_addr[2]),
    .Y(_0010_)
  );
  \$_OR_  _0576_ (
    .A(per_we[1]),
    .B(per_we[0]),
    .Y(_0011_)
  );
  \$_INV_  _0577_ (
    .A(per_addr[12]),
    .Y(_0012_)
  );
  \$_AND_  _0578_ (
    .A(per_addr[3]),
    .B(_0012_),
    .Y(_0013_)
  );
  \$_AND_  _0579_ (
    .A(per_addr[7]),
    .B(per_addr[4]),
    .Y(_0014_)
  );
  \$_AND_  _0580_ (
    .A(_0014_),
    .B(_0013_),
    .Y(_0015_)
  );
  \$_OR_  _0581_ (
    .A(per_addr[9]),
    .B(per_addr[8]),
    .Y(_0016_)
  );
  \$_OR_  _0582_ (
    .A(per_addr[11]),
    .B(per_addr[10]),
    .Y(_0017_)
  );
  \$_OR_  _0583_ (
    .A(_0017_),
    .B(_0016_),
    .Y(_0018_)
  );
  \$_INV_  _0584_ (
    .A(_0018_),
    .Y(_0019_)
  );
  \$_INV_  _0585_ (
    .A(per_addr[13]),
    .Y(_0020_)
  );
  \$_AND_  _0586_ (
    .A(_0020_),
    .B(per_en),
    .Y(_0021_)
  );
  \$_OR_  _0587_ (
    .A(per_addr[6]),
    .B(per_addr[5]),
    .Y(_0022_)
  );
  \$_INV_  _0588_ (
    .A(_0022_),
    .Y(_0023_)
  );
  \$_AND_  _0589_ (
    .A(_0023_),
    .B(_0021_),
    .Y(_0024_)
  );
  \$_AND_  _0590_ (
    .A(_0024_),
    .B(_0019_),
    .Y(_0025_)
  );
  \$_AND_  _0591_ (
    .A(_0025_),
    .B(_0015_),
    .Y(_0026_)
  );
  \$_AND_  _0592_ (
    .A(_0026_),
    .B(_0011_),
    .Y(_0027_)
  );
  \$_AND_  _0593_ (
    .A(_0027_),
    .B(_0010_),
    .Y(op2_wr)
  );
  \$_AND_  _0594_ (
    .A(sign_sel),
    .B(op1[15]),
    .Y(op1_xp[16])
  );
  \$_INV_  _0595_ (
    .A(cycle[1]),
    .Y(_0028_)
  );
  \$_AND_  _0596_ (
    .A(product[23]),
    .B(sign_sel),
    .Y(_0029_)
  );
  \$_MUX_  _0597_ (
    .A(_0029_),
    .B(product[23]),
    .S(cycle[0]),
    .Y(_0030_)
  );
  \$_XOR_  _0598_ (
    .A(_0030_),
    .B(reshi[15]),
    .Y(_0031_)
  );
  \$_INV_  _0599_ (
    .A(product[22]),
    .Y(_0032_)
  );
  \$_INV_  _0600_ (
    .A(_0029_),
    .Y(_0033_)
  );
  \$_MUX_  _0601_ (
    .A(_0033_),
    .B(_0032_),
    .S(cycle[0]),
    .Y(_0034_)
  );
  \$_INV_  _0602_ (
    .A(_0034_),
    .Y(_0035_)
  );
  \$_AND_  _0603_ (
    .A(_0035_),
    .B(reshi[14]),
    .Y(_0036_)
  );
  \$_XOR_  _0604_ (
    .A(_0034_),
    .B(reshi[14]),
    .Y(_0037_)
  );
  \$_INV_  _0605_ (
    .A(_0037_),
    .Y(_0038_)
  );
  \$_INV_  _0606_ (
    .A(product[21]),
    .Y(_0039_)
  );
  \$_MUX_  _0607_ (
    .A(_0033_),
    .B(_0039_),
    .S(cycle[0]),
    .Y(_0040_)
  );
  \$_INV_  _0608_ (
    .A(_0040_),
    .Y(_0041_)
  );
  \$_AND_  _0609_ (
    .A(_0041_),
    .B(reshi[13]),
    .Y(_0042_)
  );
  \$_XOR_  _0610_ (
    .A(_0040_),
    .B(reshi[13]),
    .Y(_0043_)
  );
  \$_INV_  _0611_ (
    .A(_0043_),
    .Y(_0044_)
  );
  \$_INV_  _0612_ (
    .A(product[20]),
    .Y(_0045_)
  );
  \$_MUX_  _0613_ (
    .A(_0033_),
    .B(_0045_),
    .S(cycle[0]),
    .Y(_0046_)
  );
  \$_INV_  _0614_ (
    .A(_0046_),
    .Y(_0047_)
  );
  \$_AND_  _0615_ (
    .A(_0047_),
    .B(reshi[12]),
    .Y(_0048_)
  );
  \$_XOR_  _0616_ (
    .A(_0046_),
    .B(reshi[12]),
    .Y(_0049_)
  );
  \$_INV_  _0617_ (
    .A(_0049_),
    .Y(_0050_)
  );
  \$_INV_  _0618_ (
    .A(product[19]),
    .Y(_0051_)
  );
  \$_MUX_  _0619_ (
    .A(_0033_),
    .B(_0051_),
    .S(cycle[0]),
    .Y(_0052_)
  );
  \$_INV_  _0620_ (
    .A(_0052_),
    .Y(_0053_)
  );
  \$_AND_  _0621_ (
    .A(_0053_),
    .B(reshi[11]),
    .Y(_0054_)
  );
  \$_XOR_  _0622_ (
    .A(_0052_),
    .B(reshi[11]),
    .Y(_0055_)
  );
  \$_INV_  _0623_ (
    .A(_0055_),
    .Y(_0056_)
  );
  \$_INV_  _0624_ (
    .A(product[18]),
    .Y(_0057_)
  );
  \$_MUX_  _0625_ (
    .A(_0033_),
    .B(_0057_),
    .S(cycle[0]),
    .Y(_0058_)
  );
  \$_INV_  _0626_ (
    .A(_0058_),
    .Y(_0059_)
  );
  \$_AND_  _0627_ (
    .A(_0059_),
    .B(reshi[10]),
    .Y(_0060_)
  );
  \$_XOR_  _0628_ (
    .A(_0058_),
    .B(reshi[10]),
    .Y(_0061_)
  );
  \$_INV_  _0629_ (
    .A(_0061_),
    .Y(_0062_)
  );
  \$_INV_  _0630_ (
    .A(product[17]),
    .Y(_0063_)
  );
  \$_MUX_  _0631_ (
    .A(_0033_),
    .B(_0063_),
    .S(cycle[0]),
    .Y(_0064_)
  );
  \$_INV_  _0632_ (
    .A(_0064_),
    .Y(_0065_)
  );
  \$_AND_  _0633_ (
    .A(_0065_),
    .B(reshi[9]),
    .Y(_0066_)
  );
  \$_XOR_  _0634_ (
    .A(_0064_),
    .B(reshi[9]),
    .Y(_0067_)
  );
  \$_INV_  _0635_ (
    .A(_0067_),
    .Y(_0068_)
  );
  \$_INV_  _0636_ (
    .A(product[16]),
    .Y(_0069_)
  );
  \$_MUX_  _0637_ (
    .A(_0033_),
    .B(_0069_),
    .S(cycle[0]),
    .Y(_0070_)
  );
  \$_INV_  _0638_ (
    .A(_0070_),
    .Y(_0071_)
  );
  \$_AND_  _0639_ (
    .A(_0071_),
    .B(reshi[8]),
    .Y(_0072_)
  );
  \$_XOR_  _0640_ (
    .A(_0070_),
    .B(reshi[8]),
    .Y(_0073_)
  );
  \$_INV_  _0641_ (
    .A(_0073_),
    .Y(_0074_)
  );
  \$_MUX_  _0642_ (
    .A(product[23]),
    .B(product[15]),
    .S(cycle[0]),
    .Y(_0075_)
  );
  \$_AND_  _0643_ (
    .A(_0075_),
    .B(reshi[7]),
    .Y(_0076_)
  );
  \$_XOR_  _0644_ (
    .A(_0075_),
    .B(reshi[7]),
    .Y(_0077_)
  );
  \$_INV_  _0645_ (
    .A(product[14]),
    .Y(_0078_)
  );
  \$_MUX_  _0646_ (
    .A(_0032_),
    .B(_0078_),
    .S(cycle[0]),
    .Y(_0079_)
  );
  \$_INV_  _0647_ (
    .A(_0079_),
    .Y(_0080_)
  );
  \$_AND_  _0648_ (
    .A(_0080_),
    .B(reshi[6]),
    .Y(_0081_)
  );
  \$_XOR_  _0649_ (
    .A(_0079_),
    .B(reshi[6]),
    .Y(_0082_)
  );
  \$_INV_  _0650_ (
    .A(_0082_),
    .Y(_0083_)
  );
  \$_INV_  _0651_ (
    .A(product[13]),
    .Y(_0084_)
  );
  \$_MUX_  _0652_ (
    .A(_0039_),
    .B(_0084_),
    .S(cycle[0]),
    .Y(_0085_)
  );
  \$_INV_  _0653_ (
    .A(_0085_),
    .Y(_0086_)
  );
  \$_AND_  _0654_ (
    .A(_0086_),
    .B(reshi[5]),
    .Y(_0087_)
  );
  \$_XOR_  _0655_ (
    .A(_0085_),
    .B(reshi[5]),
    .Y(_0088_)
  );
  \$_INV_  _0656_ (
    .A(_0088_),
    .Y(_0089_)
  );
  \$_INV_  _0657_ (
    .A(product[12]),
    .Y(_0090_)
  );
  \$_MUX_  _0658_ (
    .A(_0045_),
    .B(_0090_),
    .S(cycle[0]),
    .Y(_0091_)
  );
  \$_INV_  _0659_ (
    .A(_0091_),
    .Y(_0092_)
  );
  \$_AND_  _0660_ (
    .A(_0092_),
    .B(reshi[4]),
    .Y(_0093_)
  );
  \$_XOR_  _0661_ (
    .A(_0091_),
    .B(reshi[4]),
    .Y(_0094_)
  );
  \$_INV_  _0662_ (
    .A(_0094_),
    .Y(_0095_)
  );
  \$_INV_  _0663_ (
    .A(product[11]),
    .Y(_0096_)
  );
  \$_MUX_  _0664_ (
    .A(_0051_),
    .B(_0096_),
    .S(cycle[0]),
    .Y(_0097_)
  );
  \$_INV_  _0665_ (
    .A(_0097_),
    .Y(_0098_)
  );
  \$_AND_  _0666_ (
    .A(_0098_),
    .B(reshi[3]),
    .Y(_0099_)
  );
  \$_XOR_  _0667_ (
    .A(_0097_),
    .B(reshi[3]),
    .Y(_0100_)
  );
  \$_INV_  _0668_ (
    .A(_0100_),
    .Y(_0101_)
  );
  \$_INV_  _0669_ (
    .A(product[10]),
    .Y(_0102_)
  );
  \$_MUX_  _0670_ (
    .A(_0057_),
    .B(_0102_),
    .S(cycle[0]),
    .Y(_0103_)
  );
  \$_INV_  _0671_ (
    .A(_0103_),
    .Y(_0104_)
  );
  \$_AND_  _0672_ (
    .A(_0104_),
    .B(reshi[2]),
    .Y(_0105_)
  );
  \$_XOR_  _0673_ (
    .A(_0103_),
    .B(reshi[2]),
    .Y(_0106_)
  );
  \$_INV_  _0674_ (
    .A(_0106_),
    .Y(_0107_)
  );
  \$_INV_  _0675_ (
    .A(product[9]),
    .Y(_0108_)
  );
  \$_MUX_  _0676_ (
    .A(_0063_),
    .B(_0108_),
    .S(cycle[0]),
    .Y(_0109_)
  );
  \$_INV_  _0677_ (
    .A(_0109_),
    .Y(_0110_)
  );
  \$_AND_  _0678_ (
    .A(_0110_),
    .B(reshi[1]),
    .Y(_0111_)
  );
  \$_XOR_  _0679_ (
    .A(_0109_),
    .B(reshi[1]),
    .Y(_0112_)
  );
  \$_INV_  _0680_ (
    .A(_0112_),
    .Y(_0113_)
  );
  \$_INV_  _0681_ (
    .A(product[8]),
    .Y(_0114_)
  );
  \$_MUX_  _0682_ (
    .A(_0069_),
    .B(_0114_),
    .S(cycle[0]),
    .Y(_0115_)
  );
  \$_INV_  _0683_ (
    .A(_0115_),
    .Y(_0116_)
  );
  \$_AND_  _0684_ (
    .A(_0116_),
    .B(reshi[0]),
    .Y(_0117_)
  );
  \$_XOR_  _0685_ (
    .A(_0115_),
    .B(reshi[0]),
    .Y(_0118_)
  );
  \$_INV_  _0686_ (
    .A(_0118_),
    .Y(_0119_)
  );
  \$_MUX_  _0687_ (
    .A(product[15]),
    .B(product[7]),
    .S(cycle[0]),
    .Y(_0120_)
  );
  \$_AND_  _0688_ (
    .A(_0120_),
    .B(reslo[15]),
    .Y(_0121_)
  );
  \$_XOR_  _0689_ (
    .A(_0120_),
    .B(reslo[15]),
    .Y(_0122_)
  );
  \$_INV_  _0690_ (
    .A(product[6]),
    .Y(_0123_)
  );
  \$_MUX_  _0691_ (
    .A(_0078_),
    .B(_0123_),
    .S(cycle[0]),
    .Y(_0124_)
  );
  \$_INV_  _0692_ (
    .A(_0124_),
    .Y(_0125_)
  );
  \$_AND_  _0693_ (
    .A(_0125_),
    .B(reslo[14]),
    .Y(_0126_)
  );
  \$_XOR_  _0694_ (
    .A(_0124_),
    .B(reslo[14]),
    .Y(_0127_)
  );
  \$_INV_  _0695_ (
    .A(_0127_),
    .Y(_0128_)
  );
  \$_INV_  _0696_ (
    .A(product[5]),
    .Y(_0129_)
  );
  \$_MUX_  _0697_ (
    .A(_0084_),
    .B(_0129_),
    .S(cycle[0]),
    .Y(_0130_)
  );
  \$_INV_  _0698_ (
    .A(_0130_),
    .Y(_0131_)
  );
  \$_AND_  _0699_ (
    .A(_0131_),
    .B(reslo[13]),
    .Y(_0132_)
  );
  \$_XOR_  _0700_ (
    .A(_0130_),
    .B(reslo[13]),
    .Y(_0133_)
  );
  \$_INV_  _0701_ (
    .A(_0133_),
    .Y(_0134_)
  );
  \$_INV_  _0702_ (
    .A(product[4]),
    .Y(_0135_)
  );
  \$_MUX_  _0703_ (
    .A(_0090_),
    .B(_0135_),
    .S(cycle[0]),
    .Y(_0136_)
  );
  \$_INV_  _0704_ (
    .A(_0136_),
    .Y(_0137_)
  );
  \$_AND_  _0705_ (
    .A(_0137_),
    .B(reslo[12]),
    .Y(_0138_)
  );
  \$_XOR_  _0706_ (
    .A(_0136_),
    .B(reslo[12]),
    .Y(_0139_)
  );
  \$_INV_  _0707_ (
    .A(_0139_),
    .Y(_0140_)
  );
  \$_INV_  _0708_ (
    .A(product[3]),
    .Y(_0141_)
  );
  \$_MUX_  _0709_ (
    .A(_0096_),
    .B(_0141_),
    .S(cycle[0]),
    .Y(_0142_)
  );
  \$_INV_  _0710_ (
    .A(_0142_),
    .Y(_0143_)
  );
  \$_AND_  _0711_ (
    .A(_0143_),
    .B(reslo[11]),
    .Y(_0144_)
  );
  \$_XOR_  _0712_ (
    .A(_0142_),
    .B(reslo[11]),
    .Y(_0145_)
  );
  \$_INV_  _0713_ (
    .A(_0145_),
    .Y(_0146_)
  );
  \$_INV_  _0714_ (
    .A(product[2]),
    .Y(_0147_)
  );
  \$_MUX_  _0715_ (
    .A(_0102_),
    .B(_0147_),
    .S(cycle[0]),
    .Y(_0148_)
  );
  \$_INV_  _0716_ (
    .A(_0148_),
    .Y(_0149_)
  );
  \$_AND_  _0717_ (
    .A(_0149_),
    .B(reslo[10]),
    .Y(_0150_)
  );
  \$_XOR_  _0718_ (
    .A(_0148_),
    .B(reslo[10]),
    .Y(_0151_)
  );
  \$_INV_  _0719_ (
    .A(_0151_),
    .Y(_0152_)
  );
  \$_INV_  _0720_ (
    .A(cycle[0]),
    .Y(_0153_)
  );
  \$_INV_  _0721_ (
    .A(product[1]),
    .Y(_0154_)
  );
  \$_MUX_  _0722_ (
    .A(_0154_),
    .B(_0108_),
    .S(_0153_),
    .Y(_0155_)
  );
  \$_INV_  _0723_ (
    .A(_0155_),
    .Y(_0156_)
  );
  \$_AND_  _0724_ (
    .A(_0156_),
    .B(reslo[9]),
    .Y(_0157_)
  );
  \$_XOR_  _0725_ (
    .A(_0155_),
    .B(reslo[9]),
    .Y(_0158_)
  );
  \$_INV_  _0726_ (
    .A(_0158_),
    .Y(_0159_)
  );
  \$_INV_  _0727_ (
    .A(product[0]),
    .Y(_0160_)
  );
  \$_MUX_  _0728_ (
    .A(_0114_),
    .B(_0160_),
    .S(cycle[0]),
    .Y(_0161_)
  );
  \$_INV_  _0729_ (
    .A(_0161_),
    .Y(_0162_)
  );
  \$_AND_  _0730_ (
    .A(_0162_),
    .B(reslo[8]),
    .Y(_0163_)
  );
  \$_XOR_  _0731_ (
    .A(_0161_),
    .B(reslo[8]),
    .Y(_0164_)
  );
  \$_INV_  _0732_ (
    .A(_0164_),
    .Y(_0165_)
  );
  \$_AND_  _0733_ (
    .A(product[7]),
    .B(_0153_),
    .Y(_0166_)
  );
  \$_AND_  _0734_ (
    .A(_0166_),
    .B(reslo[7]),
    .Y(_0167_)
  );
  \$_XOR_  _0735_ (
    .A(_0166_),
    .B(reslo[7]),
    .Y(_0168_)
  );
  \$_AND_  _0736_ (
    .A(product[6]),
    .B(_0153_),
    .Y(_0169_)
  );
  \$_AND_  _0737_ (
    .A(_0169_),
    .B(reslo[6]),
    .Y(_0170_)
  );
  \$_XOR_  _0738_ (
    .A(_0169_),
    .B(reslo[6]),
    .Y(_0171_)
  );
  \$_AND_  _0739_ (
    .A(product[5]),
    .B(_0153_),
    .Y(_0172_)
  );
  \$_AND_  _0740_ (
    .A(_0172_),
    .B(reslo[5]),
    .Y(_0173_)
  );
  \$_XOR_  _0741_ (
    .A(_0172_),
    .B(reslo[5]),
    .Y(_0174_)
  );
  \$_AND_  _0742_ (
    .A(product[4]),
    .B(_0153_),
    .Y(_0175_)
  );
  \$_AND_  _0743_ (
    .A(_0175_),
    .B(reslo[4]),
    .Y(_0176_)
  );
  \$_XOR_  _0744_ (
    .A(_0175_),
    .B(reslo[4]),
    .Y(_0177_)
  );
  \$_AND_  _0745_ (
    .A(product[3]),
    .B(_0153_),
    .Y(_0178_)
  );
  \$_AND_  _0746_ (
    .A(_0178_),
    .B(reslo[3]),
    .Y(_0179_)
  );
  \$_XOR_  _0747_ (
    .A(_0178_),
    .B(reslo[3]),
    .Y(_0180_)
  );
  \$_AND_  _0748_ (
    .A(product[2]),
    .B(_0153_),
    .Y(_0181_)
  );
  \$_AND_  _0749_ (
    .A(_0181_),
    .B(reslo[2]),
    .Y(_0182_)
  );
  \$_XOR_  _0750_ (
    .A(_0181_),
    .B(reslo[2]),
    .Y(_0183_)
  );
  \$_AND_  _0751_ (
    .A(product[1]),
    .B(_0153_),
    .Y(_0184_)
  );
  \$_AND_  _0752_ (
    .A(_0184_),
    .B(reslo[1]),
    .Y(_0185_)
  );
  \$_XOR_  _0753_ (
    .A(_0184_),
    .B(reslo[1]),
    .Y(_0186_)
  );
  \$_AND_  _0754_ (
    .A(product[0]),
    .B(_0153_),
    .Y(_0187_)
  );
  \$_AND_  _0755_ (
    .A(_0187_),
    .B(reslo[0]),
    .Y(_0188_)
  );
  \$_AND_  _0756_ (
    .A(_0188_),
    .B(_0186_),
    .Y(_0189_)
  );
  \$_OR_  _0757_ (
    .A(_0189_),
    .B(_0185_),
    .Y(_0190_)
  );
  \$_AND_  _0758_ (
    .A(_0190_),
    .B(_0183_),
    .Y(_0191_)
  );
  \$_OR_  _0759_ (
    .A(_0191_),
    .B(_0182_),
    .Y(_0192_)
  );
  \$_AND_  _0760_ (
    .A(_0192_),
    .B(_0180_),
    .Y(_0193_)
  );
  \$_OR_  _0761_ (
    .A(_0193_),
    .B(_0179_),
    .Y(_0194_)
  );
  \$_AND_  _0762_ (
    .A(_0194_),
    .B(_0177_),
    .Y(_0195_)
  );
  \$_OR_  _0763_ (
    .A(_0195_),
    .B(_0176_),
    .Y(_0196_)
  );
  \$_AND_  _0764_ (
    .A(_0196_),
    .B(_0174_),
    .Y(_0197_)
  );
  \$_OR_  _0765_ (
    .A(_0197_),
    .B(_0173_),
    .Y(_0198_)
  );
  \$_AND_  _0766_ (
    .A(_0198_),
    .B(_0171_),
    .Y(_0199_)
  );
  \$_OR_  _0767_ (
    .A(_0199_),
    .B(_0170_),
    .Y(_0200_)
  );
  \$_AND_  _0768_ (
    .A(_0200_),
    .B(_0168_),
    .Y(_0201_)
  );
  \$_OR_  _0769_ (
    .A(_0201_),
    .B(_0167_),
    .Y(_0202_)
  );
  \$_AND_  _0770_ (
    .A(_0202_),
    .B(_0165_),
    .Y(_0203_)
  );
  \$_OR_  _0771_ (
    .A(_0203_),
    .B(_0163_),
    .Y(_0204_)
  );
  \$_AND_  _0772_ (
    .A(_0204_),
    .B(_0159_),
    .Y(_0205_)
  );
  \$_OR_  _0773_ (
    .A(_0205_),
    .B(_0157_),
    .Y(_0206_)
  );
  \$_AND_  _0774_ (
    .A(_0206_),
    .B(_0152_),
    .Y(_0207_)
  );
  \$_OR_  _0775_ (
    .A(_0207_),
    .B(_0150_),
    .Y(_0208_)
  );
  \$_AND_  _0776_ (
    .A(_0208_),
    .B(_0146_),
    .Y(_0209_)
  );
  \$_OR_  _0777_ (
    .A(_0209_),
    .B(_0144_),
    .Y(_0210_)
  );
  \$_AND_  _0778_ (
    .A(_0210_),
    .B(_0140_),
    .Y(_0211_)
  );
  \$_OR_  _0779_ (
    .A(_0211_),
    .B(_0138_),
    .Y(_0212_)
  );
  \$_AND_  _0780_ (
    .A(_0212_),
    .B(_0134_),
    .Y(_0213_)
  );
  \$_OR_  _0781_ (
    .A(_0213_),
    .B(_0132_),
    .Y(_0214_)
  );
  \$_AND_  _0782_ (
    .A(_0214_),
    .B(_0128_),
    .Y(_0215_)
  );
  \$_OR_  _0783_ (
    .A(_0215_),
    .B(_0126_),
    .Y(_0216_)
  );
  \$_AND_  _0784_ (
    .A(_0216_),
    .B(_0122_),
    .Y(_0217_)
  );
  \$_OR_  _0785_ (
    .A(_0217_),
    .B(_0121_),
    .Y(_0218_)
  );
  \$_AND_  _0786_ (
    .A(_0218_),
    .B(_0119_),
    .Y(_0219_)
  );
  \$_OR_  _0787_ (
    .A(_0219_),
    .B(_0117_),
    .Y(_0220_)
  );
  \$_AND_  _0788_ (
    .A(_0220_),
    .B(_0113_),
    .Y(_0221_)
  );
  \$_OR_  _0789_ (
    .A(_0221_),
    .B(_0111_),
    .Y(_0222_)
  );
  \$_AND_  _0790_ (
    .A(_0222_),
    .B(_0107_),
    .Y(_0223_)
  );
  \$_OR_  _0791_ (
    .A(_0223_),
    .B(_0105_),
    .Y(_0224_)
  );
  \$_AND_  _0792_ (
    .A(_0224_),
    .B(_0101_),
    .Y(_0225_)
  );
  \$_OR_  _0793_ (
    .A(_0225_),
    .B(_0099_),
    .Y(_0226_)
  );
  \$_AND_  _0794_ (
    .A(_0226_),
    .B(_0095_),
    .Y(_0227_)
  );
  \$_OR_  _0795_ (
    .A(_0227_),
    .B(_0093_),
    .Y(_0228_)
  );
  \$_AND_  _0796_ (
    .A(_0228_),
    .B(_0089_),
    .Y(_0229_)
  );
  \$_OR_  _0797_ (
    .A(_0229_),
    .B(_0087_),
    .Y(_0230_)
  );
  \$_AND_  _0798_ (
    .A(_0230_),
    .B(_0083_),
    .Y(_0231_)
  );
  \$_OR_  _0799_ (
    .A(_0231_),
    .B(_0081_),
    .Y(_0232_)
  );
  \$_AND_  _0800_ (
    .A(_0232_),
    .B(_0077_),
    .Y(_0233_)
  );
  \$_OR_  _0801_ (
    .A(_0233_),
    .B(_0076_),
    .Y(_0234_)
  );
  \$_AND_  _0802_ (
    .A(_0234_),
    .B(_0074_),
    .Y(_0235_)
  );
  \$_OR_  _0803_ (
    .A(_0235_),
    .B(_0072_),
    .Y(_0236_)
  );
  \$_AND_  _0804_ (
    .A(_0236_),
    .B(_0068_),
    .Y(_0237_)
  );
  \$_OR_  _0805_ (
    .A(_0237_),
    .B(_0066_),
    .Y(_0238_)
  );
  \$_AND_  _0806_ (
    .A(_0238_),
    .B(_0062_),
    .Y(_0239_)
  );
  \$_OR_  _0807_ (
    .A(_0239_),
    .B(_0060_),
    .Y(_0240_)
  );
  \$_AND_  _0808_ (
    .A(_0240_),
    .B(_0056_),
    .Y(_0241_)
  );
  \$_OR_  _0809_ (
    .A(_0241_),
    .B(_0054_),
    .Y(_0242_)
  );
  \$_AND_  _0810_ (
    .A(_0242_),
    .B(_0050_),
    .Y(_0243_)
  );
  \$_OR_  _0811_ (
    .A(_0243_),
    .B(_0048_),
    .Y(_0244_)
  );
  \$_AND_  _0812_ (
    .A(_0244_),
    .B(_0044_),
    .Y(_0245_)
  );
  \$_OR_  _0813_ (
    .A(_0245_),
    .B(_0042_),
    .Y(_0246_)
  );
  \$_AND_  _0814_ (
    .A(_0246_),
    .B(_0038_),
    .Y(_0247_)
  );
  \$_OR_  _0815_ (
    .A(_0247_),
    .B(_0036_),
    .Y(_0248_)
  );
  \$_AND_  _0816_ (
    .A(_0248_),
    .B(_0031_),
    .Y(_0249_)
  );
  \$_AND_  _0817_ (
    .A(_0030_),
    .B(reshi[15]),
    .Y(_0250_)
  );
  \$_OR_  _0818_ (
    .A(_0250_),
    .B(sumext[0]),
    .Y(_0251_)
  );
  \$_OR_  _0819_ (
    .A(_0251_),
    .B(_0249_),
    .Y(_0252_)
  );
  \$_XOR_  _0820_ (
    .A(_0248_),
    .B(_0031_),
    .Y(_0253_)
  );
  \$_MUX_  _0821_ (
    .A(_0252_),
    .B(_0253_),
    .S(sign_sel),
    .Y(_0254_)
  );
  \$_MUX_  _0822_ (
    .A(_0254_),
    .B(sumext[0]),
    .S(_0028_),
    .Y(_0255_)
  );
  \$_INV_  _0823_ (
    .A(_0011_),
    .Y(_0256_)
  );
  \$_AND_  _0824_ (
    .A(_0026_),
    .B(_0256_),
    .Y(_0257_)
  );
  \$_AND_  _0825_ (
    .A(per_addr[1]),
    .B(per_addr[0]),
    .Y(_0258_)
  );
  \$_AND_  _0826_ (
    .A(_0258_),
    .B(per_addr[2]),
    .Y(_0259_)
  );
  \$_AND_  _0827_ (
    .A(_0259_),
    .B(_0257_),
    .Y(_0260_)
  );
  \$_AND_  _0828_ (
    .A(_0260_),
    .B(_0255_),
    .Y(_0261_)
  );
  \$_XOR_  _0829_ (
    .A(_0218_),
    .B(_0119_),
    .Y(_0262_)
  );
  \$_MUX_  _0830_ (
    .A(_0262_),
    .B(reshi[0]),
    .S(_0028_),
    .Y(_0263_)
  );
  \$_AND_  _0831_ (
    .A(per_addr[1]),
    .B(_0007_),
    .Y(_0264_)
  );
  \$_AND_  _0832_ (
    .A(_0264_),
    .B(per_addr[2]),
    .Y(_0265_)
  );
  \$_AND_  _0833_ (
    .A(_0265_),
    .B(_0257_),
    .Y(_0266_)
  );
  \$_AND_  _0834_ (
    .A(_0266_),
    .B(_0263_),
    .Y(_0267_)
  );
  \$_INV_  _0835_ (
    .A(per_addr[2]),
    .Y(_0268_)
  );
  \$_AND_  _0836_ (
    .A(_0009_),
    .B(_0268_),
    .Y(_0269_)
  );
  \$_AND_  _0837_ (
    .A(_0269_),
    .B(_0257_),
    .Y(_0270_)
  );
  \$_AND_  _0838_ (
    .A(_0008_),
    .B(per_addr[0]),
    .Y(_0271_)
  );
  \$_AND_  _0839_ (
    .A(_0271_),
    .B(_0268_),
    .Y(_0272_)
  );
  \$_AND_  _0840_ (
    .A(_0272_),
    .B(_0257_),
    .Y(_0273_)
  );
  \$_OR_  _0841_ (
    .A(_0273_),
    .B(_0270_),
    .Y(_0274_)
  );
  \$_AND_  _0842_ (
    .A(_0264_),
    .B(_0268_),
    .Y(_0275_)
  );
  \$_AND_  _0843_ (
    .A(_0275_),
    .B(_0257_),
    .Y(_0276_)
  );
  \$_AND_  _0844_ (
    .A(_0258_),
    .B(_0268_),
    .Y(_0277_)
  );
  \$_AND_  _0845_ (
    .A(_0277_),
    .B(_0257_),
    .Y(_0278_)
  );
  \$_OR_  _0846_ (
    .A(_0278_),
    .B(_0276_),
    .Y(_0279_)
  );
  \$_OR_  _0847_ (
    .A(_0279_),
    .B(_0274_),
    .Y(_0280_)
  );
  \$_AND_  _0848_ (
    .A(_0280_),
    .B(op1[0]),
    .Y(_0281_)
  );
  \$_AND_  _0849_ (
    .A(_0257_),
    .B(_0010_),
    .Y(_0282_)
  );
  \$_AND_  _0850_ (
    .A(_0282_),
    .B(op2[0]),
    .Y(_0283_)
  );
  \$_XOR_  _0851_ (
    .A(_0187_),
    .B(reslo[0]),
    .Y(_0284_)
  );
  \$_MUX_  _0852_ (
    .A(_0284_),
    .B(reslo[0]),
    .S(_0028_),
    .Y(_0285_)
  );
  \$_AND_  _0853_ (
    .A(_0271_),
    .B(per_addr[2]),
    .Y(_0286_)
  );
  \$_AND_  _0854_ (
    .A(_0286_),
    .B(_0257_),
    .Y(_0287_)
  );
  \$_AND_  _0855_ (
    .A(_0287_),
    .B(_0285_),
    .Y(_0288_)
  );
  \$_OR_  _0856_ (
    .A(_0288_),
    .B(_0283_),
    .Y(_0289_)
  );
  \$_OR_  _0857_ (
    .A(_0289_),
    .B(_0281_),
    .Y(_0290_)
  );
  \$_OR_  _0858_ (
    .A(_0290_),
    .B(_0267_),
    .Y(_0291_)
  );
  \$_OR_  _0859_ (
    .A(_0291_),
    .B(_0261_),
    .Y(per_dout[0])
  );
  \$_AND_  _0860_ (
    .A(_0253_),
    .B(sign_sel),
    .Y(_0292_)
  );
  \$_MUX_  _0861_ (
    .A(_0292_),
    .B(sumext[15]),
    .S(_0028_),
    .Y(_0293_)
  );
  \$_AND_  _0862_ (
    .A(_0293_),
    .B(_0260_),
    .Y(_0294_)
  );
  \$_XOR_  _0863_ (
    .A(_0238_),
    .B(_0062_),
    .Y(_0295_)
  );
  \$_MUX_  _0864_ (
    .A(_0295_),
    .B(reshi[10]),
    .S(_0028_),
    .Y(_0296_)
  );
  \$_AND_  _0865_ (
    .A(_0296_),
    .B(_0266_),
    .Y(_0297_)
  );
  \$_XOR_  _0866_ (
    .A(_0206_),
    .B(_0152_),
    .Y(_0298_)
  );
  \$_MUX_  _0867_ (
    .A(_0298_),
    .B(reslo[10]),
    .S(_0028_),
    .Y(_0299_)
  );
  \$_AND_  _0868_ (
    .A(_0299_),
    .B(_0287_),
    .Y(_0300_)
  );
  \$_AND_  _0869_ (
    .A(_0280_),
    .B(op1[10]),
    .Y(_0301_)
  );
  \$_AND_  _0870_ (
    .A(_0282_),
    .B(op2[10]),
    .Y(_0302_)
  );
  \$_OR_  _0871_ (
    .A(_0302_),
    .B(_0301_),
    .Y(_0303_)
  );
  \$_OR_  _0872_ (
    .A(_0303_),
    .B(_0300_),
    .Y(_0304_)
  );
  \$_OR_  _0873_ (
    .A(_0304_),
    .B(_0297_),
    .Y(_0305_)
  );
  \$_OR_  _0874_ (
    .A(_0305_),
    .B(_0294_),
    .Y(per_dout[10])
  );
  \$_XOR_  _0875_ (
    .A(_0240_),
    .B(_0056_),
    .Y(_0306_)
  );
  \$_MUX_  _0876_ (
    .A(_0306_),
    .B(reshi[11]),
    .S(_0028_),
    .Y(_0307_)
  );
  \$_AND_  _0877_ (
    .A(_0307_),
    .B(_0266_),
    .Y(_0308_)
  );
  \$_XOR_  _0878_ (
    .A(_0208_),
    .B(_0146_),
    .Y(_0309_)
  );
  \$_MUX_  _0879_ (
    .A(_0309_),
    .B(reslo[11]),
    .S(_0028_),
    .Y(_0310_)
  );
  \$_AND_  _0880_ (
    .A(_0310_),
    .B(_0287_),
    .Y(_0311_)
  );
  \$_AND_  _0881_ (
    .A(_0280_),
    .B(op1[11]),
    .Y(_0312_)
  );
  \$_AND_  _0882_ (
    .A(_0282_),
    .B(op2[11]),
    .Y(_0313_)
  );
  \$_OR_  _0883_ (
    .A(_0313_),
    .B(_0312_),
    .Y(_0314_)
  );
  \$_OR_  _0884_ (
    .A(_0314_),
    .B(_0311_),
    .Y(_0315_)
  );
  \$_OR_  _0885_ (
    .A(_0315_),
    .B(_0308_),
    .Y(_0316_)
  );
  \$_OR_  _0886_ (
    .A(_0316_),
    .B(_0294_),
    .Y(per_dout[11])
  );
  \$_XOR_  _0887_ (
    .A(_0242_),
    .B(_0050_),
    .Y(_0317_)
  );
  \$_MUX_  _0888_ (
    .A(_0317_),
    .B(reshi[12]),
    .S(_0028_),
    .Y(_0318_)
  );
  \$_AND_  _0889_ (
    .A(_0318_),
    .B(_0266_),
    .Y(_0319_)
  );
  \$_XOR_  _0890_ (
    .A(_0210_),
    .B(_0140_),
    .Y(_0320_)
  );
  \$_MUX_  _0891_ (
    .A(_0320_),
    .B(reslo[12]),
    .S(_0028_),
    .Y(_0321_)
  );
  \$_AND_  _0892_ (
    .A(_0321_),
    .B(_0287_),
    .Y(_0322_)
  );
  \$_AND_  _0893_ (
    .A(_0280_),
    .B(op1[12]),
    .Y(_0323_)
  );
  \$_AND_  _0894_ (
    .A(_0282_),
    .B(op2[12]),
    .Y(_0324_)
  );
  \$_OR_  _0895_ (
    .A(_0324_),
    .B(_0323_),
    .Y(_0325_)
  );
  \$_OR_  _0896_ (
    .A(_0325_),
    .B(_0322_),
    .Y(_0326_)
  );
  \$_OR_  _0897_ (
    .A(_0326_),
    .B(_0319_),
    .Y(_0327_)
  );
  \$_OR_  _0898_ (
    .A(_0327_),
    .B(_0294_),
    .Y(per_dout[12])
  );
  \$_XOR_  _0899_ (
    .A(_0244_),
    .B(_0044_),
    .Y(_0328_)
  );
  \$_MUX_  _0900_ (
    .A(_0328_),
    .B(reshi[13]),
    .S(_0028_),
    .Y(_0329_)
  );
  \$_AND_  _0901_ (
    .A(_0329_),
    .B(_0266_),
    .Y(_0330_)
  );
  \$_XOR_  _0902_ (
    .A(_0212_),
    .B(_0134_),
    .Y(_0331_)
  );
  \$_MUX_  _0903_ (
    .A(_0331_),
    .B(reslo[13]),
    .S(_0028_),
    .Y(_0332_)
  );
  \$_AND_  _0904_ (
    .A(_0332_),
    .B(_0287_),
    .Y(_0333_)
  );
  \$_AND_  _0905_ (
    .A(_0280_),
    .B(op1[13]),
    .Y(_0334_)
  );
  \$_AND_  _0906_ (
    .A(_0282_),
    .B(op2[13]),
    .Y(_0335_)
  );
  \$_OR_  _0907_ (
    .A(_0335_),
    .B(_0334_),
    .Y(_0336_)
  );
  \$_OR_  _0908_ (
    .A(_0336_),
    .B(_0333_),
    .Y(_0337_)
  );
  \$_OR_  _0909_ (
    .A(_0337_),
    .B(_0330_),
    .Y(_0338_)
  );
  \$_OR_  _0910_ (
    .A(_0338_),
    .B(_0294_),
    .Y(per_dout[13])
  );
  \$_XOR_  _0911_ (
    .A(_0246_),
    .B(_0038_),
    .Y(_0339_)
  );
  \$_MUX_  _0912_ (
    .A(_0339_),
    .B(reshi[14]),
    .S(_0028_),
    .Y(_0340_)
  );
  \$_AND_  _0913_ (
    .A(_0340_),
    .B(_0266_),
    .Y(_0341_)
  );
  \$_XOR_  _0914_ (
    .A(_0214_),
    .B(_0128_),
    .Y(_0342_)
  );
  \$_MUX_  _0915_ (
    .A(_0342_),
    .B(reslo[14]),
    .S(_0028_),
    .Y(_0343_)
  );
  \$_AND_  _0916_ (
    .A(_0343_),
    .B(_0287_),
    .Y(_0344_)
  );
  \$_AND_  _0917_ (
    .A(_0280_),
    .B(op1[14]),
    .Y(_0345_)
  );
  \$_AND_  _0918_ (
    .A(_0282_),
    .B(op2[14]),
    .Y(_0346_)
  );
  \$_OR_  _0919_ (
    .A(_0346_),
    .B(_0345_),
    .Y(_0347_)
  );
  \$_OR_  _0920_ (
    .A(_0347_),
    .B(_0344_),
    .Y(_0348_)
  );
  \$_OR_  _0921_ (
    .A(_0348_),
    .B(_0341_),
    .Y(_0349_)
  );
  \$_OR_  _0922_ (
    .A(_0349_),
    .B(_0294_),
    .Y(per_dout[14])
  );
  \$_MUX_  _0923_ (
    .A(_0253_),
    .B(reshi[15]),
    .S(_0028_),
    .Y(_0350_)
  );
  \$_AND_  _0924_ (
    .A(_0350_),
    .B(_0266_),
    .Y(_0351_)
  );
  \$_XOR_  _0925_ (
    .A(_0216_),
    .B(_0122_),
    .Y(_0352_)
  );
  \$_MUX_  _0926_ (
    .A(_0352_),
    .B(reslo[15]),
    .S(_0028_),
    .Y(_0353_)
  );
  \$_AND_  _0927_ (
    .A(_0353_),
    .B(_0287_),
    .Y(_0354_)
  );
  \$_AND_  _0928_ (
    .A(_0280_),
    .B(op1[15]),
    .Y(_0355_)
  );
  \$_AND_  _0929_ (
    .A(_0282_),
    .B(op2[15]),
    .Y(_0356_)
  );
  \$_OR_  _0930_ (
    .A(_0356_),
    .B(_0355_),
    .Y(_0357_)
  );
  \$_OR_  _0931_ (
    .A(_0357_),
    .B(_0354_),
    .Y(_0358_)
  );
  \$_OR_  _0932_ (
    .A(_0358_),
    .B(_0351_),
    .Y(_0359_)
  );
  \$_OR_  _0933_ (
    .A(_0359_),
    .B(_0294_),
    .Y(per_dout[15])
  );
  \$_XOR_  _0934_ (
    .A(_0220_),
    .B(_0113_),
    .Y(_0360_)
  );
  \$_MUX_  _0935_ (
    .A(_0360_),
    .B(reshi[1]),
    .S(_0028_),
    .Y(_0361_)
  );
  \$_AND_  _0936_ (
    .A(_0361_),
    .B(_0266_),
    .Y(_0362_)
  );
  \$_AND_  _0937_ (
    .A(_0280_),
    .B(op1[1]),
    .Y(_0363_)
  );
  \$_AND_  _0938_ (
    .A(_0282_),
    .B(op2[1]),
    .Y(_0364_)
  );
  \$_XOR_  _0939_ (
    .A(_0188_),
    .B(_0186_),
    .Y(_0365_)
  );
  \$_MUX_  _0940_ (
    .A(_0365_),
    .B(reslo[1]),
    .S(_0028_),
    .Y(_0366_)
  );
  \$_AND_  _0941_ (
    .A(_0366_),
    .B(_0287_),
    .Y(_0367_)
  );
  \$_OR_  _0942_ (
    .A(_0367_),
    .B(_0364_),
    .Y(_0368_)
  );
  \$_OR_  _0943_ (
    .A(_0368_),
    .B(_0363_),
    .Y(_0369_)
  );
  \$_OR_  _0944_ (
    .A(_0369_),
    .B(_0362_),
    .Y(_0370_)
  );
  \$_OR_  _0945_ (
    .A(_0370_),
    .B(_0294_),
    .Y(per_dout[1])
  );
  \$_XOR_  _0946_ (
    .A(_0222_),
    .B(_0107_),
    .Y(_0371_)
  );
  \$_MUX_  _0947_ (
    .A(_0371_),
    .B(reshi[2]),
    .S(_0028_),
    .Y(_0372_)
  );
  \$_AND_  _0948_ (
    .A(_0372_),
    .B(_0266_),
    .Y(_0373_)
  );
  \$_XOR_  _0949_ (
    .A(_0190_),
    .B(_0183_),
    .Y(_0374_)
  );
  \$_MUX_  _0950_ (
    .A(_0374_),
    .B(reslo[2]),
    .S(_0028_),
    .Y(_0375_)
  );
  \$_AND_  _0951_ (
    .A(_0375_),
    .B(_0287_),
    .Y(_0376_)
  );
  \$_AND_  _0952_ (
    .A(_0280_),
    .B(op1[2]),
    .Y(_0377_)
  );
  \$_AND_  _0953_ (
    .A(_0282_),
    .B(op2[2]),
    .Y(_0378_)
  );
  \$_OR_  _0954_ (
    .A(_0378_),
    .B(_0377_),
    .Y(_0379_)
  );
  \$_OR_  _0955_ (
    .A(_0379_),
    .B(_0376_),
    .Y(_0380_)
  );
  \$_OR_  _0956_ (
    .A(_0380_),
    .B(_0373_),
    .Y(_0381_)
  );
  \$_OR_  _0957_ (
    .A(_0381_),
    .B(_0294_),
    .Y(per_dout[2])
  );
  \$_XOR_  _0958_ (
    .A(_0224_),
    .B(_0101_),
    .Y(_0382_)
  );
  \$_MUX_  _0959_ (
    .A(_0382_),
    .B(reshi[3]),
    .S(_0028_),
    .Y(_0383_)
  );
  \$_AND_  _0960_ (
    .A(_0383_),
    .B(_0266_),
    .Y(_0384_)
  );
  \$_XOR_  _0961_ (
    .A(_0192_),
    .B(_0180_),
    .Y(_0385_)
  );
  \$_MUX_  _0962_ (
    .A(_0385_),
    .B(reslo[3]),
    .S(_0028_),
    .Y(_0386_)
  );
  \$_AND_  _0963_ (
    .A(_0386_),
    .B(_0287_),
    .Y(_0387_)
  );
  \$_AND_  _0964_ (
    .A(_0280_),
    .B(op1[3]),
    .Y(_0388_)
  );
  \$_AND_  _0965_ (
    .A(_0282_),
    .B(op2[3]),
    .Y(_0389_)
  );
  \$_OR_  _0966_ (
    .A(_0389_),
    .B(_0388_),
    .Y(_0390_)
  );
  \$_OR_  _0967_ (
    .A(_0390_),
    .B(_0387_),
    .Y(_0391_)
  );
  \$_OR_  _0968_ (
    .A(_0391_),
    .B(_0384_),
    .Y(_0392_)
  );
  \$_OR_  _0969_ (
    .A(_0392_),
    .B(_0294_),
    .Y(per_dout[3])
  );
  \$_XOR_  _0970_ (
    .A(_0226_),
    .B(_0095_),
    .Y(_0393_)
  );
  \$_MUX_  _0971_ (
    .A(_0393_),
    .B(reshi[4]),
    .S(_0028_),
    .Y(_0394_)
  );
  \$_AND_  _0972_ (
    .A(_0394_),
    .B(_0266_),
    .Y(_0395_)
  );
  \$_XOR_  _0973_ (
    .A(_0194_),
    .B(_0177_),
    .Y(_0396_)
  );
  \$_MUX_  _0974_ (
    .A(_0396_),
    .B(reslo[4]),
    .S(_0028_),
    .Y(_0397_)
  );
  \$_AND_  _0975_ (
    .A(_0397_),
    .B(_0287_),
    .Y(_0398_)
  );
  \$_AND_  _0976_ (
    .A(_0280_),
    .B(op1[4]),
    .Y(_0399_)
  );
  \$_AND_  _0977_ (
    .A(_0282_),
    .B(op2[4]),
    .Y(_0400_)
  );
  \$_OR_  _0978_ (
    .A(_0400_),
    .B(_0399_),
    .Y(_0401_)
  );
  \$_OR_  _0979_ (
    .A(_0401_),
    .B(_0398_),
    .Y(_0402_)
  );
  \$_OR_  _0980_ (
    .A(_0402_),
    .B(_0395_),
    .Y(_0403_)
  );
  \$_OR_  _0981_ (
    .A(_0403_),
    .B(_0294_),
    .Y(per_dout[4])
  );
  \$_XOR_  _0982_ (
    .A(_0228_),
    .B(_0089_),
    .Y(_0404_)
  );
  \$_MUX_  _0983_ (
    .A(_0404_),
    .B(reshi[5]),
    .S(_0028_),
    .Y(_0405_)
  );
  \$_AND_  _0984_ (
    .A(_0405_),
    .B(_0266_),
    .Y(_0406_)
  );
  \$_XOR_  _0985_ (
    .A(_0196_),
    .B(_0174_),
    .Y(_0407_)
  );
  \$_MUX_  _0986_ (
    .A(_0407_),
    .B(reslo[5]),
    .S(_0028_),
    .Y(_0408_)
  );
  \$_AND_  _0987_ (
    .A(_0408_),
    .B(_0287_),
    .Y(_0409_)
  );
  \$_AND_  _0988_ (
    .A(_0280_),
    .B(op1[5]),
    .Y(_0410_)
  );
  \$_AND_  _0989_ (
    .A(_0282_),
    .B(op2[5]),
    .Y(_0411_)
  );
  \$_OR_  _0990_ (
    .A(_0411_),
    .B(_0410_),
    .Y(_0412_)
  );
  \$_OR_  _0991_ (
    .A(_0412_),
    .B(_0409_),
    .Y(_0413_)
  );
  \$_OR_  _0992_ (
    .A(_0413_),
    .B(_0406_),
    .Y(_0414_)
  );
  \$_OR_  _0993_ (
    .A(_0414_),
    .B(_0294_),
    .Y(per_dout[5])
  );
  \$_XOR_  _0994_ (
    .A(_0230_),
    .B(_0083_),
    .Y(_0415_)
  );
  \$_MUX_  _0995_ (
    .A(_0415_),
    .B(reshi[6]),
    .S(_0028_),
    .Y(_0416_)
  );
  \$_AND_  _0996_ (
    .A(_0416_),
    .B(_0266_),
    .Y(_0417_)
  );
  \$_XOR_  _0997_ (
    .A(_0198_),
    .B(_0171_),
    .Y(_0418_)
  );
  \$_MUX_  _0998_ (
    .A(_0418_),
    .B(reslo[6]),
    .S(_0028_),
    .Y(_0419_)
  );
  \$_AND_  _0999_ (
    .A(_0419_),
    .B(_0287_),
    .Y(_0420_)
  );
  \$_AND_  _1000_ (
    .A(_0280_),
    .B(op1[6]),
    .Y(_0421_)
  );
  \$_AND_  _1001_ (
    .A(_0282_),
    .B(op2[6]),
    .Y(_0422_)
  );
  \$_OR_  _1002_ (
    .A(_0422_),
    .B(_0421_),
    .Y(_0423_)
  );
  \$_OR_  _1003_ (
    .A(_0423_),
    .B(_0420_),
    .Y(_0424_)
  );
  \$_OR_  _1004_ (
    .A(_0424_),
    .B(_0417_),
    .Y(_0425_)
  );
  \$_OR_  _1005_ (
    .A(_0425_),
    .B(_0294_),
    .Y(per_dout[6])
  );
  \$_XOR_  _1006_ (
    .A(_0232_),
    .B(_0077_),
    .Y(_0426_)
  );
  \$_MUX_  _1007_ (
    .A(_0426_),
    .B(reshi[7]),
    .S(_0028_),
    .Y(_0427_)
  );
  \$_AND_  _1008_ (
    .A(_0427_),
    .B(_0266_),
    .Y(_0428_)
  );
  \$_XOR_  _1009_ (
    .A(_0200_),
    .B(_0168_),
    .Y(_0429_)
  );
  \$_MUX_  _1010_ (
    .A(_0429_),
    .B(reslo[7]),
    .S(_0028_),
    .Y(_0430_)
  );
  \$_AND_  _1011_ (
    .A(_0430_),
    .B(_0287_),
    .Y(_0431_)
  );
  \$_AND_  _1012_ (
    .A(_0280_),
    .B(op1[7]),
    .Y(_0432_)
  );
  \$_AND_  _1013_ (
    .A(_0282_),
    .B(op2[7]),
    .Y(_0433_)
  );
  \$_OR_  _1014_ (
    .A(_0433_),
    .B(_0432_),
    .Y(_0434_)
  );
  \$_OR_  _1015_ (
    .A(_0434_),
    .B(_0431_),
    .Y(_0435_)
  );
  \$_OR_  _1016_ (
    .A(_0435_),
    .B(_0428_),
    .Y(_0436_)
  );
  \$_OR_  _1017_ (
    .A(_0436_),
    .B(_0294_),
    .Y(per_dout[7])
  );
  \$_XOR_  _1018_ (
    .A(_0234_),
    .B(_0074_),
    .Y(_0437_)
  );
  \$_MUX_  _1019_ (
    .A(_0437_),
    .B(reshi[8]),
    .S(_0028_),
    .Y(_0438_)
  );
  \$_AND_  _1020_ (
    .A(_0438_),
    .B(_0266_),
    .Y(_0439_)
  );
  \$_XOR_  _1021_ (
    .A(_0202_),
    .B(_0165_),
    .Y(_0440_)
  );
  \$_MUX_  _1022_ (
    .A(_0440_),
    .B(reslo[8]),
    .S(_0028_),
    .Y(_0441_)
  );
  \$_AND_  _1023_ (
    .A(_0441_),
    .B(_0287_),
    .Y(_0442_)
  );
  \$_AND_  _1024_ (
    .A(_0280_),
    .B(op1[8]),
    .Y(_0443_)
  );
  \$_AND_  _1025_ (
    .A(_0282_),
    .B(op2[8]),
    .Y(_0444_)
  );
  \$_OR_  _1026_ (
    .A(_0444_),
    .B(_0443_),
    .Y(_0445_)
  );
  \$_OR_  _1027_ (
    .A(_0445_),
    .B(_0442_),
    .Y(_0446_)
  );
  \$_OR_  _1028_ (
    .A(_0446_),
    .B(_0439_),
    .Y(_0447_)
  );
  \$_OR_  _1029_ (
    .A(_0447_),
    .B(_0294_),
    .Y(per_dout[8])
  );
  \$_XOR_  _1030_ (
    .A(_0236_),
    .B(_0068_),
    .Y(_0448_)
  );
  \$_MUX_  _1031_ (
    .A(_0448_),
    .B(reshi[9]),
    .S(_0028_),
    .Y(_0449_)
  );
  \$_AND_  _1032_ (
    .A(_0449_),
    .B(_0266_),
    .Y(_0450_)
  );
  \$_XOR_  _1033_ (
    .A(_0204_),
    .B(_0159_),
    .Y(_0451_)
  );
  \$_MUX_  _1034_ (
    .A(_0451_),
    .B(reslo[9]),
    .S(_0028_),
    .Y(_0452_)
  );
  \$_AND_  _1035_ (
    .A(_0452_),
    .B(_0287_),
    .Y(_0453_)
  );
  \$_AND_  _1036_ (
    .A(_0280_),
    .B(op1[9]),
    .Y(_0454_)
  );
  \$_AND_  _1037_ (
    .A(_0282_),
    .B(op2[9]),
    .Y(_0455_)
  );
  \$_OR_  _1038_ (
    .A(_0455_),
    .B(_0454_),
    .Y(_0456_)
  );
  \$_OR_  _1039_ (
    .A(_0456_),
    .B(_0453_),
    .Y(_0457_)
  );
  \$_OR_  _1040_ (
    .A(_0457_),
    .B(_0450_),
    .Y(_0458_)
  );
  \$_OR_  _1041_ (
    .A(_0458_),
    .B(_0294_),
    .Y(per_dout[9])
  );
  \$_INV_  _1042_ (
    .A(_0027_),
    .Y(_0459_)
  );
  \$_INV_  _1043_ (
    .A(_0269_),
    .Y(_0460_)
  );
  \$_OR_  _1044_ (
    .A(_0460_),
    .B(_0459_),
    .Y(_0461_)
  );
  \$_AND_  _1045_ (
    .A(_0272_),
    .B(_0027_),
    .Y(_0462_)
  );
  \$_INV_  _1046_ (
    .A(_0462_),
    .Y(_0463_)
  );
  \$_AND_  _1047_ (
    .A(_0463_),
    .B(_0461_),
    .Y(_0464_)
  );
  \$_AND_  _1048_ (
    .A(_0275_),
    .B(_0027_),
    .Y(_0465_)
  );
  \$_AND_  _1049_ (
    .A(_0277_),
    .B(_0027_),
    .Y(_0466_)
  );
  \$_OR_  _1050_ (
    .A(_0466_),
    .B(_0465_),
    .Y(_0467_)
  );
  \$_INV_  _1051_ (
    .A(_0467_),
    .Y(_0468_)
  );
  \$_AND_  _1052_ (
    .A(_0468_),
    .B(_0464_),
    .Y(_0469_)
  );
  \$_MUX_  _1053_ (
    .A(per_din[0]),
    .B(op1[0]),
    .S(_0469_),
    .Y(_0001_[0])
  );
  \$_MUX_  _1054_ (
    .A(per_din[10]),
    .B(op1[10]),
    .S(_0469_),
    .Y(_0001_[10])
  );
  \$_MUX_  _1055_ (
    .A(per_din[11]),
    .B(op1[11]),
    .S(_0469_),
    .Y(_0001_[11])
  );
  \$_MUX_  _1056_ (
    .A(per_din[12]),
    .B(op1[12]),
    .S(_0469_),
    .Y(_0001_[12])
  );
  \$_MUX_  _1057_ (
    .A(per_din[13]),
    .B(op1[13]),
    .S(_0469_),
    .Y(_0001_[13])
  );
  \$_MUX_  _1058_ (
    .A(per_din[14]),
    .B(op1[14]),
    .S(_0469_),
    .Y(_0001_[14])
  );
  \$_MUX_  _1059_ (
    .A(per_din[15]),
    .B(op1[15]),
    .S(_0469_),
    .Y(_0001_[15])
  );
  \$_MUX_  _1060_ (
    .A(per_din[1]),
    .B(op1[1]),
    .S(_0469_),
    .Y(_0001_[1])
  );
  \$_MUX_  _1061_ (
    .A(per_din[2]),
    .B(op1[2]),
    .S(_0469_),
    .Y(_0001_[2])
  );
  \$_MUX_  _1062_ (
    .A(per_din[3]),
    .B(op1[3]),
    .S(_0469_),
    .Y(_0001_[3])
  );
  \$_MUX_  _1063_ (
    .A(per_din[4]),
    .B(op1[4]),
    .S(_0469_),
    .Y(_0001_[4])
  );
  \$_MUX_  _1064_ (
    .A(per_din[5]),
    .B(op1[5]),
    .S(_0469_),
    .Y(_0001_[5])
  );
  \$_MUX_  _1065_ (
    .A(per_din[6]),
    .B(op1[6]),
    .S(_0469_),
    .Y(_0001_[6])
  );
  \$_MUX_  _1066_ (
    .A(per_din[7]),
    .B(op1[7]),
    .S(_0469_),
    .Y(_0001_[7])
  );
  \$_MUX_  _1067_ (
    .A(per_din[8]),
    .B(op1[8]),
    .S(_0469_),
    .Y(_0001_[8])
  );
  \$_MUX_  _1068_ (
    .A(per_din[9]),
    .B(op1[9]),
    .S(_0469_),
    .Y(_0001_[9])
  );
  \$_MUX_  _1069_ (
    .A(op2[0]),
    .B(per_din[0]),
    .S(op2_wr),
    .Y(_0002_[0])
  );
  \$_MUX_  _1070_ (
    .A(op2[10]),
    .B(per_din[10]),
    .S(op2_wr),
    .Y(_0002_[10])
  );
  \$_MUX_  _1071_ (
    .A(op2[11]),
    .B(per_din[11]),
    .S(op2_wr),
    .Y(_0002_[11])
  );
  \$_MUX_  _1072_ (
    .A(op2[12]),
    .B(per_din[12]),
    .S(op2_wr),
    .Y(_0002_[12])
  );
  \$_MUX_  _1073_ (
    .A(op2[13]),
    .B(per_din[13]),
    .S(op2_wr),
    .Y(_0002_[13])
  );
  \$_MUX_  _1074_ (
    .A(op2[14]),
    .B(per_din[14]),
    .S(op2_wr),
    .Y(_0002_[14])
  );
  \$_MUX_  _1075_ (
    .A(op2[15]),
    .B(per_din[15]),
    .S(op2_wr),
    .Y(_0002_[15])
  );
  \$_MUX_  _1076_ (
    .A(op2[1]),
    .B(per_din[1]),
    .S(op2_wr),
    .Y(_0002_[1])
  );
  \$_MUX_  _1077_ (
    .A(op2[2]),
    .B(per_din[2]),
    .S(op2_wr),
    .Y(_0002_[2])
  );
  \$_MUX_  _1078_ (
    .A(op2[3]),
    .B(per_din[3]),
    .S(op2_wr),
    .Y(_0002_[3])
  );
  \$_MUX_  _1079_ (
    .A(op2[4]),
    .B(per_din[4]),
    .S(op2_wr),
    .Y(_0002_[4])
  );
  \$_MUX_  _1080_ (
    .A(op2[5]),
    .B(per_din[5]),
    .S(op2_wr),
    .Y(_0002_[5])
  );
  \$_MUX_  _1081_ (
    .A(op2[6]),
    .B(per_din[6]),
    .S(op2_wr),
    .Y(_0002_[6])
  );
  \$_MUX_  _1082_ (
    .A(op2[7]),
    .B(per_din[7]),
    .S(op2_wr),
    .Y(_0002_[7])
  );
  \$_MUX_  _1083_ (
    .A(op2[8]),
    .B(per_din[8]),
    .S(op2_wr),
    .Y(_0002_[8])
  );
  \$_MUX_  _1084_ (
    .A(op2[9]),
    .B(per_din[9]),
    .S(op2_wr),
    .Y(_0002_[9])
  );
  \$_INV_  _1085_ (
    .A(op2_wr),
    .Y(_0470_)
  );
  \$_OR_  _1086_ (
    .A(_0470_),
    .B(acc_sel),
    .Y(_0471_)
  );
  \$_AND_  _1087_ (
    .A(_0286_),
    .B(_0027_),
    .Y(_0472_)
  );
  \$_INV_  _1088_ (
    .A(_0472_),
    .Y(_0473_)
  );
  \$_AND_  _1089_ (
    .A(_0028_),
    .B(_0153_),
    .Y(_0474_)
  );
  \$_AND_  _1090_ (
    .A(_0285_),
    .B(_0473_),
    .Y(_0475_)
  );
  \$_AND_  _1091_ (
    .A(_0475_),
    .B(_0471_),
    .Y(_0476_)
  );
  \$_AND_  _1092_ (
    .A(_0472_),
    .B(per_din[0]),
    .Y(_0477_)
  );
  \$_OR_  _1093_ (
    .A(_0477_),
    .B(_0476_),
    .Y(_0004_[0])
  );
  \$_MUX_  _1094_ (
    .A(_0298_),
    .B(reslo[10]),
    .S(_0474_),
    .Y(_0478_)
  );
  \$_AND_  _1095_ (
    .A(_0473_),
    .B(_0471_),
    .Y(_0479_)
  );
  \$_AND_  _1096_ (
    .A(_0479_),
    .B(_0478_),
    .Y(_0480_)
  );
  \$_AND_  _1097_ (
    .A(_0472_),
    .B(per_din[10]),
    .Y(_0481_)
  );
  \$_OR_  _1098_ (
    .A(_0481_),
    .B(_0480_),
    .Y(_0004_[10])
  );
  \$_MUX_  _1099_ (
    .A(_0309_),
    .B(reslo[11]),
    .S(_0474_),
    .Y(_0482_)
  );
  \$_AND_  _1100_ (
    .A(_0482_),
    .B(_0479_),
    .Y(_0483_)
  );
  \$_AND_  _1101_ (
    .A(_0472_),
    .B(per_din[11]),
    .Y(_0484_)
  );
  \$_OR_  _1102_ (
    .A(_0484_),
    .B(_0483_),
    .Y(_0004_[11])
  );
  \$_MUX_  _1103_ (
    .A(_0320_),
    .B(reslo[12]),
    .S(_0474_),
    .Y(_0485_)
  );
  \$_AND_  _1104_ (
    .A(_0485_),
    .B(_0479_),
    .Y(_0486_)
  );
  \$_AND_  _1105_ (
    .A(_0472_),
    .B(per_din[12]),
    .Y(_0487_)
  );
  \$_OR_  _1106_ (
    .A(_0487_),
    .B(_0486_),
    .Y(_0004_[12])
  );
  \$_MUX_  _1107_ (
    .A(_0331_),
    .B(reslo[13]),
    .S(_0474_),
    .Y(_0488_)
  );
  \$_AND_  _1108_ (
    .A(_0488_),
    .B(_0479_),
    .Y(_0489_)
  );
  \$_AND_  _1109_ (
    .A(_0472_),
    .B(per_din[13]),
    .Y(_0490_)
  );
  \$_OR_  _1110_ (
    .A(_0490_),
    .B(_0489_),
    .Y(_0004_[13])
  );
  \$_MUX_  _1111_ (
    .A(_0342_),
    .B(reslo[14]),
    .S(_0474_),
    .Y(_0491_)
  );
  \$_AND_  _1112_ (
    .A(_0491_),
    .B(_0479_),
    .Y(_0492_)
  );
  \$_AND_  _1113_ (
    .A(_0472_),
    .B(per_din[14]),
    .Y(_0493_)
  );
  \$_OR_  _1114_ (
    .A(_0493_),
    .B(_0492_),
    .Y(_0004_[14])
  );
  \$_MUX_  _1115_ (
    .A(_0352_),
    .B(reslo[15]),
    .S(_0474_),
    .Y(_0494_)
  );
  \$_AND_  _1116_ (
    .A(_0494_),
    .B(_0479_),
    .Y(_0495_)
  );
  \$_AND_  _1117_ (
    .A(_0472_),
    .B(per_din[15]),
    .Y(_0496_)
  );
  \$_OR_  _1118_ (
    .A(_0496_),
    .B(_0495_),
    .Y(_0004_[15])
  );
  \$_AND_  _1119_ (
    .A(_0366_),
    .B(_0479_),
    .Y(_0497_)
  );
  \$_AND_  _1120_ (
    .A(_0472_),
    .B(per_din[1]),
    .Y(_0498_)
  );
  \$_OR_  _1121_ (
    .A(_0498_),
    .B(_0497_),
    .Y(_0004_[1])
  );
  \$_AND_  _1122_ (
    .A(_0375_),
    .B(_0479_),
    .Y(_0499_)
  );
  \$_AND_  _1123_ (
    .A(_0472_),
    .B(per_din[2]),
    .Y(_0500_)
  );
  \$_OR_  _1124_ (
    .A(_0500_),
    .B(_0499_),
    .Y(_0004_[2])
  );
  \$_AND_  _1125_ (
    .A(_0386_),
    .B(_0479_),
    .Y(_0501_)
  );
  \$_AND_  _1126_ (
    .A(_0472_),
    .B(per_din[3]),
    .Y(_0502_)
  );
  \$_OR_  _1127_ (
    .A(_0502_),
    .B(_0501_),
    .Y(_0004_[3])
  );
  \$_AND_  _1128_ (
    .A(_0397_),
    .B(_0479_),
    .Y(_0503_)
  );
  \$_AND_  _1129_ (
    .A(_0472_),
    .B(per_din[4]),
    .Y(_0504_)
  );
  \$_OR_  _1130_ (
    .A(_0504_),
    .B(_0503_),
    .Y(_0004_[4])
  );
  \$_AND_  _1131_ (
    .A(_0408_),
    .B(_0479_),
    .Y(_0505_)
  );
  \$_AND_  _1132_ (
    .A(_0472_),
    .B(per_din[5]),
    .Y(_0506_)
  );
  \$_OR_  _1133_ (
    .A(_0506_),
    .B(_0505_),
    .Y(_0004_[5])
  );
  \$_AND_  _1134_ (
    .A(_0419_),
    .B(_0479_),
    .Y(_0507_)
  );
  \$_AND_  _1135_ (
    .A(_0472_),
    .B(per_din[6]),
    .Y(_0508_)
  );
  \$_OR_  _1136_ (
    .A(_0508_),
    .B(_0507_),
    .Y(_0004_[6])
  );
  \$_AND_  _1137_ (
    .A(_0430_),
    .B(_0479_),
    .Y(_0509_)
  );
  \$_AND_  _1138_ (
    .A(_0472_),
    .B(per_din[7]),
    .Y(_0510_)
  );
  \$_OR_  _1139_ (
    .A(_0510_),
    .B(_0509_),
    .Y(_0004_[7])
  );
  \$_MUX_  _1140_ (
    .A(_0440_),
    .B(reslo[8]),
    .S(_0474_),
    .Y(_0511_)
  );
  \$_AND_  _1141_ (
    .A(_0511_),
    .B(_0479_),
    .Y(_0512_)
  );
  \$_AND_  _1142_ (
    .A(_0472_),
    .B(per_din[8]),
    .Y(_0513_)
  );
  \$_OR_  _1143_ (
    .A(_0513_),
    .B(_0512_),
    .Y(_0004_[8])
  );
  \$_MUX_  _1144_ (
    .A(_0451_),
    .B(reslo[9]),
    .S(_0474_),
    .Y(_0514_)
  );
  \$_AND_  _1145_ (
    .A(_0514_),
    .B(_0479_),
    .Y(_0515_)
  );
  \$_AND_  _1146_ (
    .A(_0472_),
    .B(per_din[9]),
    .Y(_0516_)
  );
  \$_OR_  _1147_ (
    .A(_0516_),
    .B(_0515_),
    .Y(_0004_[9])
  );
  \$_MUX_  _1148_ (
    .A(_0262_),
    .B(reshi[0]),
    .S(_0474_),
    .Y(_0517_)
  );
  \$_AND_  _1149_ (
    .A(_0265_),
    .B(_0027_),
    .Y(_0518_)
  );
  \$_INV_  _1150_ (
    .A(_0518_),
    .Y(_0519_)
  );
  \$_AND_  _1151_ (
    .A(_0519_),
    .B(_0471_),
    .Y(_0520_)
  );
  \$_AND_  _1152_ (
    .A(_0520_),
    .B(_0517_),
    .Y(_0521_)
  );
  \$_AND_  _1153_ (
    .A(_0518_),
    .B(per_din[0]),
    .Y(_0522_)
  );
  \$_OR_  _1154_ (
    .A(_0522_),
    .B(_0521_),
    .Y(_0003_[0])
  );
  \$_MUX_  _1155_ (
    .A(_0295_),
    .B(reshi[10]),
    .S(_0474_),
    .Y(_0523_)
  );
  \$_AND_  _1156_ (
    .A(_0523_),
    .B(_0520_),
    .Y(_0524_)
  );
  \$_AND_  _1157_ (
    .A(_0518_),
    .B(per_din[10]),
    .Y(_0525_)
  );
  \$_OR_  _1158_ (
    .A(_0525_),
    .B(_0524_),
    .Y(_0003_[10])
  );
  \$_MUX_  _1159_ (
    .A(_0306_),
    .B(reshi[11]),
    .S(_0474_),
    .Y(_0526_)
  );
  \$_AND_  _1160_ (
    .A(_0526_),
    .B(_0520_),
    .Y(_0527_)
  );
  \$_AND_  _1161_ (
    .A(_0518_),
    .B(per_din[11]),
    .Y(_0528_)
  );
  \$_OR_  _1162_ (
    .A(_0528_),
    .B(_0527_),
    .Y(_0003_[11])
  );
  \$_MUX_  _1163_ (
    .A(_0317_),
    .B(reshi[12]),
    .S(_0474_),
    .Y(_0529_)
  );
  \$_AND_  _1164_ (
    .A(_0529_),
    .B(_0520_),
    .Y(_0530_)
  );
  \$_AND_  _1165_ (
    .A(_0518_),
    .B(per_din[12]),
    .Y(_0531_)
  );
  \$_OR_  _1166_ (
    .A(_0531_),
    .B(_0530_),
    .Y(_0003_[12])
  );
  \$_MUX_  _1167_ (
    .A(_0328_),
    .B(reshi[13]),
    .S(_0474_),
    .Y(_0532_)
  );
  \$_AND_  _1168_ (
    .A(_0532_),
    .B(_0520_),
    .Y(_0533_)
  );
  \$_AND_  _1169_ (
    .A(_0518_),
    .B(per_din[13]),
    .Y(_0534_)
  );
  \$_OR_  _1170_ (
    .A(_0534_),
    .B(_0533_),
    .Y(_0003_[13])
  );
  \$_MUX_  _1171_ (
    .A(_0339_),
    .B(reshi[14]),
    .S(_0474_),
    .Y(_0535_)
  );
  \$_AND_  _1172_ (
    .A(_0535_),
    .B(_0520_),
    .Y(_0536_)
  );
  \$_AND_  _1173_ (
    .A(_0518_),
    .B(per_din[14]),
    .Y(_0537_)
  );
  \$_OR_  _1174_ (
    .A(_0537_),
    .B(_0536_),
    .Y(_0003_[14])
  );
  \$_MUX_  _1175_ (
    .A(_0253_),
    .B(reshi[15]),
    .S(_0474_),
    .Y(_0538_)
  );
  \$_AND_  _1176_ (
    .A(_0538_),
    .B(_0520_),
    .Y(_0539_)
  );
  \$_AND_  _1177_ (
    .A(_0518_),
    .B(per_din[15]),
    .Y(_0540_)
  );
  \$_OR_  _1178_ (
    .A(_0540_),
    .B(_0539_),
    .Y(_0003_[15])
  );
  \$_MUX_  _1179_ (
    .A(_0360_),
    .B(reshi[1]),
    .S(_0474_),
    .Y(_0541_)
  );
  \$_AND_  _1180_ (
    .A(_0541_),
    .B(_0520_),
    .Y(_0542_)
  );
  \$_AND_  _1181_ (
    .A(_0518_),
    .B(per_din[1]),
    .Y(_0543_)
  );
  \$_OR_  _1182_ (
    .A(_0543_),
    .B(_0542_),
    .Y(_0003_[1])
  );
  \$_MUX_  _1183_ (
    .A(_0371_),
    .B(reshi[2]),
    .S(_0474_),
    .Y(_0544_)
  );
  \$_AND_  _1184_ (
    .A(_0544_),
    .B(_0520_),
    .Y(_0545_)
  );
  \$_AND_  _1185_ (
    .A(_0518_),
    .B(per_din[2]),
    .Y(_0546_)
  );
  \$_OR_  _1186_ (
    .A(_0546_),
    .B(_0545_),
    .Y(_0003_[2])
  );
  \$_MUX_  _1187_ (
    .A(_0382_),
    .B(reshi[3]),
    .S(_0474_),
    .Y(_0547_)
  );
  \$_AND_  _1188_ (
    .A(_0547_),
    .B(_0520_),
    .Y(_0548_)
  );
  \$_AND_  _1189_ (
    .A(_0518_),
    .B(per_din[3]),
    .Y(_0549_)
  );
  \$_OR_  _1190_ (
    .A(_0549_),
    .B(_0548_),
    .Y(_0003_[3])
  );
  \$_MUX_  _1191_ (
    .A(_0393_),
    .B(reshi[4]),
    .S(_0474_),
    .Y(_0550_)
  );
  \$_AND_  _1192_ (
    .A(_0550_),
    .B(_0520_),
    .Y(_0551_)
  );
  \$_AND_  _1193_ (
    .A(_0518_),
    .B(per_din[4]),
    .Y(_0552_)
  );
  \$_OR_  _1194_ (
    .A(_0552_),
    .B(_0551_),
    .Y(_0003_[4])
  );
  \$_MUX_  _1195_ (
    .A(_0404_),
    .B(reshi[5]),
    .S(_0474_),
    .Y(_0553_)
  );
  \$_AND_  _1196_ (
    .A(_0553_),
    .B(_0520_),
    .Y(_0554_)
  );
  \$_AND_  _1197_ (
    .A(_0518_),
    .B(per_din[5]),
    .Y(_0555_)
  );
  \$_OR_  _1198_ (
    .A(_0555_),
    .B(_0554_),
    .Y(_0003_[5])
  );
  \$_MUX_  _1199_ (
    .A(_0415_),
    .B(reshi[6]),
    .S(_0474_),
    .Y(_0556_)
  );
  \$_AND_  _1200_ (
    .A(_0556_),
    .B(_0520_),
    .Y(_0557_)
  );
  \$_AND_  _1201_ (
    .A(_0518_),
    .B(per_din[6]),
    .Y(_0558_)
  );
  \$_OR_  _1202_ (
    .A(_0558_),
    .B(_0557_),
    .Y(_0003_[6])
  );
  \$_MUX_  _1203_ (
    .A(_0426_),
    .B(reshi[7]),
    .S(_0474_),
    .Y(_0559_)
  );
  \$_AND_  _1204_ (
    .A(_0559_),
    .B(_0520_),
    .Y(_0560_)
  );
  \$_AND_  _1205_ (
    .A(_0518_),
    .B(per_din[7]),
    .Y(_0561_)
  );
  \$_OR_  _1206_ (
    .A(_0561_),
    .B(_0560_),
    .Y(_0003_[7])
  );
  \$_MUX_  _1207_ (
    .A(_0437_),
    .B(reshi[8]),
    .S(_0474_),
    .Y(_0562_)
  );
  \$_AND_  _1208_ (
    .A(_0562_),
    .B(_0520_),
    .Y(_0563_)
  );
  \$_AND_  _1209_ (
    .A(_0518_),
    .B(per_din[8]),
    .Y(_0564_)
  );
  \$_OR_  _1210_ (
    .A(_0564_),
    .B(_0563_),
    .Y(_0003_[8])
  );
  \$_MUX_  _1211_ (
    .A(_0448_),
    .B(reshi[9]),
    .S(_0474_),
    .Y(_0565_)
  );
  \$_AND_  _1212_ (
    .A(_0565_),
    .B(_0520_),
    .Y(_0566_)
  );
  \$_AND_  _1213_ (
    .A(_0518_),
    .B(per_din[9]),
    .Y(_0567_)
  );
  \$_OR_  _1214_ (
    .A(_0567_),
    .B(_0566_),
    .Y(_0003_[9])
  );
  \$_MUX_  _1215_ (
    .A(_0254_),
    .B(sumext[0]),
    .S(_0474_),
    .Y(_0568_)
  );
  \$_AND_  _1216_ (
    .A(_0568_),
    .B(_0470_),
    .Y(_0006_[0])
  );
  \$_MUX_  _1217_ (
    .A(_0292_),
    .B(sumext[15]),
    .S(_0474_),
    .Y(_0569_)
  );
  \$_AND_  _1218_ (
    .A(_0569_),
    .B(_0470_),
    .Y(_0006_[1])
  );
  \$_OR_  _1219_ (
    .A(_0466_),
    .B(_0462_),
    .Y(_0570_)
  );
  \$_MUX_  _1220_ (
    .A(_0570_),
    .B(sign_sel),
    .S(_0469_),
    .Y(_0005_)
  );
  \$_MUX_  _1221_ (
    .A(_0467_),
    .B(acc_sel),
    .S(_0469_),
    .Y(_0000_)
  );
  \$_MUX_  _1222_ (
    .A(op2[0]),
    .B(op2[8]),
    .S(cycle[0]),
    .Y(op2_xp[0])
  );
  \$_MUX_  _1223_ (
    .A(op2[1]),
    .B(op2[9]),
    .S(cycle[0]),
    .Y(op2_xp[1])
  );
  \$_MUX_  _1224_ (
    .A(op2[2]),
    .B(op2[10]),
    .S(cycle[0]),
    .Y(op2_xp[2])
  );
  \$_MUX_  _1225_ (
    .A(op2[3]),
    .B(op2[11]),
    .S(cycle[0]),
    .Y(op2_xp[3])
  );
  \$_MUX_  _1226_ (
    .A(op2[4]),
    .B(op2[12]),
    .S(cycle[0]),
    .Y(op2_xp[4])
  );
  \$_MUX_  _1227_ (
    .A(op2[5]),
    .B(op2[13]),
    .S(cycle[0]),
    .Y(op2_xp[5])
  );
  \$_MUX_  _1228_ (
    .A(op2[6]),
    .B(op2[14]),
    .S(cycle[0]),
    .Y(op2_xp[6])
  );
  \$_MUX_  _1229_ (
    .A(op2[7]),
    .B(op2[15]),
    .S(cycle[0]),
    .Y(op2_xp[7])
  );
  \$_AND_  _1230_ (
    .A(cycle[0]),
    .B(op2[15]),
    .Y(_0571_)
  );
  \$_AND_  _1231_ (
    .A(_0571_),
    .B(sign_sel),
    .Y(op2_xp[8])
  );
  \$mul  #(
    .A_SIGNED(1),
    .A_WIDTH(17),
    .B_SIGNED(1),
    .B_WIDTH(9),
    .Y_WIDTH(26)
  ) _1232_ (
    .A({ op1_xp[16], op1 }),
    .B(op2_xp),
    .Y(product)
  );
  \$_DFF_PP0_  \op1_reg[0]  /* _1233_ */ (
    .C(mclk),
    .D(_0001_[0]),
    .Q(op1[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[10]  /* _1234_ */ (
    .C(mclk),
    .D(_0001_[10]),
    .Q(op1[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[11]  /* _1235_ */ (
    .C(mclk),
    .D(_0001_[11]),
    .Q(op1[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[12]  /* _1236_ */ (
    .C(mclk),
    .D(_0001_[12]),
    .Q(op1[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[13]  /* _1237_ */ (
    .C(mclk),
    .D(_0001_[13]),
    .Q(op1[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[14]  /* _1238_ */ (
    .C(mclk),
    .D(_0001_[14]),
    .Q(op1[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[15]  /* _1239_ */ (
    .C(mclk),
    .D(_0001_[15]),
    .Q(op1[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[1]  /* _1240_ */ (
    .C(mclk),
    .D(_0001_[1]),
    .Q(op1[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[2]  /* _1241_ */ (
    .C(mclk),
    .D(_0001_[2]),
    .Q(op1[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[3]  /* _1242_ */ (
    .C(mclk),
    .D(_0001_[3]),
    .Q(op1[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[4]  /* _1243_ */ (
    .C(mclk),
    .D(_0001_[4]),
    .Q(op1[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[5]  /* _1244_ */ (
    .C(mclk),
    .D(_0001_[5]),
    .Q(op1[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[6]  /* _1245_ */ (
    .C(mclk),
    .D(_0001_[6]),
    .Q(op1[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[7]  /* _1246_ */ (
    .C(mclk),
    .D(_0001_[7]),
    .Q(op1[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[8]  /* _1247_ */ (
    .C(mclk),
    .D(_0001_[8]),
    .Q(op1[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op1_reg[9]  /* _1248_ */ (
    .C(mclk),
    .D(_0001_[9]),
    .Q(op1[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[0]  /* _1249_ */ (
    .C(mclk),
    .D(_0002_[0]),
    .Q(op2[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[10]  /* _1250_ */ (
    .C(mclk),
    .D(_0002_[10]),
    .Q(op2[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[11]  /* _1251_ */ (
    .C(mclk),
    .D(_0002_[11]),
    .Q(op2[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[12]  /* _1252_ */ (
    .C(mclk),
    .D(_0002_[12]),
    .Q(op2[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[13]  /* _1253_ */ (
    .C(mclk),
    .D(_0002_[13]),
    .Q(op2[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[14]  /* _1254_ */ (
    .C(mclk),
    .D(_0002_[14]),
    .Q(op2[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[15]  /* _1255_ */ (
    .C(mclk),
    .D(_0002_[15]),
    .Q(op2[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[1]  /* _1256_ */ (
    .C(mclk),
    .D(_0002_[1]),
    .Q(op2[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[2]  /* _1257_ */ (
    .C(mclk),
    .D(_0002_[2]),
    .Q(op2[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[3]  /* _1258_ */ (
    .C(mclk),
    .D(_0002_[3]),
    .Q(op2[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[4]  /* _1259_ */ (
    .C(mclk),
    .D(_0002_[4]),
    .Q(op2[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[5]  /* _1260_ */ (
    .C(mclk),
    .D(_0002_[5]),
    .Q(op2[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[6]  /* _1261_ */ (
    .C(mclk),
    .D(_0002_[6]),
    .Q(op2[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[7]  /* _1262_ */ (
    .C(mclk),
    .D(_0002_[7]),
    .Q(op2[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[8]  /* _1263_ */ (
    .C(mclk),
    .D(_0002_[8]),
    .Q(op2[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \op2_reg[9]  /* _1264_ */ (
    .C(mclk),
    .D(_0002_[9]),
    .Q(op2[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[0]  /* _1265_ */ (
    .C(mclk),
    .D(_0004_[0]),
    .Q(reslo[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[10]  /* _1266_ */ (
    .C(mclk),
    .D(_0004_[10]),
    .Q(reslo[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[11]  /* _1267_ */ (
    .C(mclk),
    .D(_0004_[11]),
    .Q(reslo[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[12]  /* _1268_ */ (
    .C(mclk),
    .D(_0004_[12]),
    .Q(reslo[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[13]  /* _1269_ */ (
    .C(mclk),
    .D(_0004_[13]),
    .Q(reslo[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[14]  /* _1270_ */ (
    .C(mclk),
    .D(_0004_[14]),
    .Q(reslo[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[15]  /* _1271_ */ (
    .C(mclk),
    .D(_0004_[15]),
    .Q(reslo[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[1]  /* _1272_ */ (
    .C(mclk),
    .D(_0004_[1]),
    .Q(reslo[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[2]  /* _1273_ */ (
    .C(mclk),
    .D(_0004_[2]),
    .Q(reslo[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[3]  /* _1274_ */ (
    .C(mclk),
    .D(_0004_[3]),
    .Q(reslo[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[4]  /* _1275_ */ (
    .C(mclk),
    .D(_0004_[4]),
    .Q(reslo[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[5]  /* _1276_ */ (
    .C(mclk),
    .D(_0004_[5]),
    .Q(reslo[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[6]  /* _1277_ */ (
    .C(mclk),
    .D(_0004_[6]),
    .Q(reslo[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[7]  /* _1278_ */ (
    .C(mclk),
    .D(_0004_[7]),
    .Q(reslo[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[8]  /* _1279_ */ (
    .C(mclk),
    .D(_0004_[8]),
    .Q(reslo[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reslo_reg[9]  /* _1280_ */ (
    .C(mclk),
    .D(_0004_[9]),
    .Q(reslo[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[0]  /* _1281_ */ (
    .C(mclk),
    .D(_0003_[0]),
    .Q(reshi[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[10]  /* _1282_ */ (
    .C(mclk),
    .D(_0003_[10]),
    .Q(reshi[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[11]  /* _1283_ */ (
    .C(mclk),
    .D(_0003_[11]),
    .Q(reshi[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[12]  /* _1284_ */ (
    .C(mclk),
    .D(_0003_[12]),
    .Q(reshi[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[13]  /* _1285_ */ (
    .C(mclk),
    .D(_0003_[13]),
    .Q(reshi[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[14]  /* _1286_ */ (
    .C(mclk),
    .D(_0003_[14]),
    .Q(reshi[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[15]  /* _1287_ */ (
    .C(mclk),
    .D(_0003_[15]),
    .Q(reshi[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[1]  /* _1288_ */ (
    .C(mclk),
    .D(_0003_[1]),
    .Q(reshi[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[2]  /* _1289_ */ (
    .C(mclk),
    .D(_0003_[2]),
    .Q(reshi[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[3]  /* _1290_ */ (
    .C(mclk),
    .D(_0003_[3]),
    .Q(reshi[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[4]  /* _1291_ */ (
    .C(mclk),
    .D(_0003_[4]),
    .Q(reshi[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[5]  /* _1292_ */ (
    .C(mclk),
    .D(_0003_[5]),
    .Q(reshi[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[6]  /* _1293_ */ (
    .C(mclk),
    .D(_0003_[6]),
    .Q(reshi[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[7]  /* _1294_ */ (
    .C(mclk),
    .D(_0003_[7]),
    .Q(reshi[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[8]  /* _1295_ */ (
    .C(mclk),
    .D(_0003_[8]),
    .Q(reshi[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \reshi_reg[9]  /* _1296_ */ (
    .C(mclk),
    .D(_0003_[9]),
    .Q(reshi[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \sumext_reg[0]  /* _1297_ */ (
    .C(mclk),
    .D(_0006_[0]),
    .Q(sumext[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \sumext_reg[15]  /* _1298_ */ (
    .C(mclk),
    .D(_0006_[1]),
    .Q(sumext[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  sign_sel_reg /* _1299_ */ (
    .C(mclk),
    .D(_0005_),
    .Q(sign_sel),
    .R(puc_rst)
  );
  \$_DFF_PP0_  acc_sel_reg /* _1300_ */ (
    .C(mclk),
    .D(_0000_),
    .Q(acc_sel),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \cycle_reg[0]  /* _1301_ */ (
    .C(mclk),
    .D(op2_wr),
    .Q(cycle[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \cycle_reg[1]  /* _1302_ */ (
    .C(mclk),
    .D(cycle[0]),
    .Q(cycle[1]),
    .R(puc_rst)
  );
  assign early_read = cycle[1];
  assign mclk_op1 = mclk;
  assign mclk_op2 = mclk;
  assign mclk_reshi = mclk;
  assign mclk_reslo = mclk;
  assign op1_rd = op1;
  assign op1_xp[15:0] = op1;
  assign op2_hi_xp[7:0] = op2[15:8];
  assign op2_lo_xp = { 1'b0, op2[7:0] };
  assign op2_rd = op2;
  assign reg_addr = { per_addr[2:0], 1'b0 };
  assign { reg_wr[15], reg_wr[13], reg_wr[11], reg_wr[9:7], reg_wr[5], reg_wr[3], reg_wr[1] } = { 4'b0000, op2_wr, 4'b0000 };
  assign result = { reshi, reslo };
  assign sumext[14:1] = { sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15], sumext[15] };
  assign sumext_s = { sumext[15], sumext[0] };
endmodule

module omsp_register_file(cpuoff, gie, oscoff, pc_sw, pc_sw_wr, reg_dest, reg_src, scg0, scg1, status, alu_stat, alu_stat_wr, inst_bw, inst_dest, inst_src, mclk, pc, puc_rst, reg_dest_val, reg_dest_wr, reg_pc_call, reg_sp_val, reg_sp_wr, reg_sr_wr, reg_sr_clr, reg_incr, scan_enable);
  wire [15:0] _0000_;
  wire [15:0] _0001_;
  wire [15:0] _0002_;
  wire [15:0] _0003_;
  wire [15:0] _0004_;
  wire [15:0] _0005_;
  wire [15:0] _0006_;
  wire [15:0] _0007_;
  wire [15:0] _0008_;
  wire [15:0] _0009_;
  wire [15:0] _0010_;
  wire [15:0] _0011_;
  wire [15:0] _0012_;
  wire [15:0] _0013_;
  wire [15:0] _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  input [3:0] alu_stat;
  input [3:0] alu_stat_wr;
  output cpuoff;
  output gie;
  input inst_bw;
  input [15:0] inst_dest;
  input [15:0] inst_src;
  input mclk;
  wire mclk_r1;
  wire mclk_r10;
  wire mclk_r11;
  wire mclk_r12;
  wire mclk_r13;
  wire mclk_r14;
  wire mclk_r15;
  wire mclk_r2;
  wire mclk_r3;
  wire mclk_r4;
  wire mclk_r5;
  wire mclk_r6;
  wire mclk_r7;
  wire mclk_r8;
  wire mclk_r9;
  output oscoff;
  input [15:0] pc;
  output [15:0] pc_sw;
  output pc_sw_wr;
  input puc_rst;
  wire [15:0] r0;
  wire [15:0] r1;
  wire [15:0] r10;
  wire [15:0] r11;
  wire [15:0] r12;
  wire [15:0] r13;
  wire [15:0] r14;
  wire [15:0] r15;
  wire [15:0] r2;
  wire [15:0] r3;
  wire [15:0] r4;
  wire [15:0] r5;
  wire [15:0] r6;
  wire [15:0] r7;
  wire [15:0] r8;
  wire [15:0] r9;
  output [15:0] reg_dest;
  input [15:0] reg_dest_val;
  wire [15:0] reg_dest_val_in;
  input reg_dest_wr;
  input reg_incr;
  input reg_pc_call;
  input [15:0] reg_sp_val;
  input reg_sp_wr;
  input reg_sr_clr;
  input reg_sr_wr;
  output [15:0] reg_src;
  input scan_enable;
  output scg0;
  output scg1;
  output [3:0] status;
  \$_OR_  _1299_ (
    .A(inst_src[2]),
    .B(reg_sr_clr),
    .Y(_0912_)
  );
  \$_AND_  _1300_ (
    .A(_0912_),
    .B(r2[0]),
    .Y(_0913_)
  );
  \$_INV_  _1301_ (
    .A(reg_sr_clr),
    .Y(_0914_)
  );
  \$_AND_  _1302_ (
    .A(inst_src[0]),
    .B(_0914_),
    .Y(_0915_)
  );
  \$_AND_  _1303_ (
    .A(_0915_),
    .B(pc[0]),
    .Y(_0916_)
  );
  \$_AND_  _1304_ (
    .A(inst_src[1]),
    .B(_0914_),
    .Y(_0917_)
  );
  \$_AND_  _1305_ (
    .A(_0917_),
    .B(r1[0]),
    .Y(_0918_)
  );
  \$_OR_  _1306_ (
    .A(_0918_),
    .B(_0916_),
    .Y(_0919_)
  );
  \$_AND_  _1307_ (
    .A(inst_src[3]),
    .B(_0914_),
    .Y(_0920_)
  );
  \$_AND_  _1308_ (
    .A(_0920_),
    .B(r3[0]),
    .Y(_0921_)
  );
  \$_AND_  _1309_ (
    .A(inst_src[4]),
    .B(_0914_),
    .Y(_0922_)
  );
  \$_AND_  _1310_ (
    .A(_0922_),
    .B(r4[0]),
    .Y(_0923_)
  );
  \$_OR_  _1311_ (
    .A(_0923_),
    .B(_0921_),
    .Y(_0924_)
  );
  \$_OR_  _1312_ (
    .A(_0924_),
    .B(_0919_),
    .Y(_0925_)
  );
  \$_OR_  _1313_ (
    .A(_0925_),
    .B(_0913_),
    .Y(_0926_)
  );
  \$_AND_  _1314_ (
    .A(inst_src[15]),
    .B(_0914_),
    .Y(_0927_)
  );
  \$_AND_  _1315_ (
    .A(_0927_),
    .B(r15[0]),
    .Y(_0928_)
  );
  \$_AND_  _1316_ (
    .A(inst_src[13]),
    .B(_0914_),
    .Y(_0929_)
  );
  \$_AND_  _1317_ (
    .A(_0929_),
    .B(r13[0]),
    .Y(_0930_)
  );
  \$_AND_  _1318_ (
    .A(inst_src[14]),
    .B(_0914_),
    .Y(_0931_)
  );
  \$_AND_  _1319_ (
    .A(_0931_),
    .B(r14[0]),
    .Y(_0932_)
  );
  \$_OR_  _1320_ (
    .A(_0932_),
    .B(_0930_),
    .Y(_0933_)
  );
  \$_OR_  _1321_ (
    .A(_0933_),
    .B(_0928_),
    .Y(_0934_)
  );
  \$_AND_  _1322_ (
    .A(inst_src[9]),
    .B(_0914_),
    .Y(_0935_)
  );
  \$_AND_  _1323_ (
    .A(_0935_),
    .B(r9[0]),
    .Y(_0936_)
  );
  \$_AND_  _1324_ (
    .A(inst_src[10]),
    .B(_0914_),
    .Y(_0937_)
  );
  \$_AND_  _1325_ (
    .A(_0937_),
    .B(r10[0]),
    .Y(_0938_)
  );
  \$_OR_  _1326_ (
    .A(_0938_),
    .B(_0936_),
    .Y(_0939_)
  );
  \$_AND_  _1327_ (
    .A(inst_src[11]),
    .B(_0914_),
    .Y(_0940_)
  );
  \$_AND_  _1328_ (
    .A(_0940_),
    .B(r11[0]),
    .Y(_0941_)
  );
  \$_AND_  _1329_ (
    .A(inst_src[12]),
    .B(_0914_),
    .Y(_0942_)
  );
  \$_AND_  _1330_ (
    .A(_0942_),
    .B(r12[0]),
    .Y(_0943_)
  );
  \$_OR_  _1331_ (
    .A(_0943_),
    .B(_0941_),
    .Y(_0944_)
  );
  \$_OR_  _1332_ (
    .A(_0944_),
    .B(_0939_),
    .Y(_0945_)
  );
  \$_AND_  _1333_ (
    .A(inst_src[5]),
    .B(_0914_),
    .Y(_0946_)
  );
  \$_AND_  _1334_ (
    .A(_0946_),
    .B(r5[0]),
    .Y(_0947_)
  );
  \$_AND_  _1335_ (
    .A(inst_src[6]),
    .B(_0914_),
    .Y(_0948_)
  );
  \$_AND_  _1336_ (
    .A(_0948_),
    .B(r6[0]),
    .Y(_0949_)
  );
  \$_OR_  _1337_ (
    .A(_0949_),
    .B(_0947_),
    .Y(_0950_)
  );
  \$_AND_  _1338_ (
    .A(inst_src[7]),
    .B(_0914_),
    .Y(_0951_)
  );
  \$_AND_  _1339_ (
    .A(_0951_),
    .B(r7[0]),
    .Y(_0952_)
  );
  \$_AND_  _1340_ (
    .A(inst_src[8]),
    .B(_0914_),
    .Y(_0953_)
  );
  \$_AND_  _1341_ (
    .A(_0953_),
    .B(r8[0]),
    .Y(_0954_)
  );
  \$_OR_  _1342_ (
    .A(_0954_),
    .B(_0952_),
    .Y(_0955_)
  );
  \$_OR_  _1343_ (
    .A(_0955_),
    .B(_0950_),
    .Y(_0956_)
  );
  \$_OR_  _1344_ (
    .A(_0956_),
    .B(_0945_),
    .Y(_0957_)
  );
  \$_OR_  _1345_ (
    .A(_0957_),
    .B(_0934_),
    .Y(_0958_)
  );
  \$_OR_  _1346_ (
    .A(_0958_),
    .B(_0926_),
    .Y(reg_src[0])
  );
  \$_AND_  _1347_ (
    .A(_0912_),
    .B(r2[15]),
    .Y(_0959_)
  );
  \$_AND_  _1348_ (
    .A(_0915_),
    .B(pc[10]),
    .Y(_0960_)
  );
  \$_AND_  _1349_ (
    .A(_0917_),
    .B(r1[10]),
    .Y(_0961_)
  );
  \$_OR_  _1350_ (
    .A(_0961_),
    .B(_0960_),
    .Y(_0962_)
  );
  \$_AND_  _1351_ (
    .A(_0920_),
    .B(r3[10]),
    .Y(_0963_)
  );
  \$_AND_  _1352_ (
    .A(_0922_),
    .B(r4[10]),
    .Y(_0964_)
  );
  \$_OR_  _1353_ (
    .A(_0964_),
    .B(_0963_),
    .Y(_0965_)
  );
  \$_OR_  _1354_ (
    .A(_0965_),
    .B(_0962_),
    .Y(_0966_)
  );
  \$_OR_  _1355_ (
    .A(_0966_),
    .B(_0959_),
    .Y(_0967_)
  );
  \$_AND_  _1356_ (
    .A(_0927_),
    .B(r15[10]),
    .Y(_0968_)
  );
  \$_AND_  _1357_ (
    .A(_0929_),
    .B(r13[10]),
    .Y(_0969_)
  );
  \$_AND_  _1358_ (
    .A(_0931_),
    .B(r14[10]),
    .Y(_0970_)
  );
  \$_OR_  _1359_ (
    .A(_0970_),
    .B(_0969_),
    .Y(_0971_)
  );
  \$_OR_  _1360_ (
    .A(_0971_),
    .B(_0968_),
    .Y(_0972_)
  );
  \$_AND_  _1361_ (
    .A(_0935_),
    .B(r9[10]),
    .Y(_0973_)
  );
  \$_AND_  _1362_ (
    .A(_0937_),
    .B(r10[10]),
    .Y(_0974_)
  );
  \$_OR_  _1363_ (
    .A(_0974_),
    .B(_0973_),
    .Y(_0975_)
  );
  \$_AND_  _1364_ (
    .A(_0940_),
    .B(r11[10]),
    .Y(_0976_)
  );
  \$_AND_  _1365_ (
    .A(_0942_),
    .B(r12[10]),
    .Y(_0977_)
  );
  \$_OR_  _1366_ (
    .A(_0977_),
    .B(_0976_),
    .Y(_0978_)
  );
  \$_OR_  _1367_ (
    .A(_0978_),
    .B(_0975_),
    .Y(_0979_)
  );
  \$_AND_  _1368_ (
    .A(_0946_),
    .B(r5[10]),
    .Y(_0980_)
  );
  \$_AND_  _1369_ (
    .A(_0948_),
    .B(r6[10]),
    .Y(_0981_)
  );
  \$_OR_  _1370_ (
    .A(_0981_),
    .B(_0980_),
    .Y(_0982_)
  );
  \$_AND_  _1371_ (
    .A(_0951_),
    .B(r7[10]),
    .Y(_0983_)
  );
  \$_AND_  _1372_ (
    .A(_0953_),
    .B(r8[10]),
    .Y(_0984_)
  );
  \$_OR_  _1373_ (
    .A(_0984_),
    .B(_0983_),
    .Y(_0985_)
  );
  \$_OR_  _1374_ (
    .A(_0985_),
    .B(_0982_),
    .Y(_0986_)
  );
  \$_OR_  _1375_ (
    .A(_0986_),
    .B(_0979_),
    .Y(_0987_)
  );
  \$_OR_  _1376_ (
    .A(_0987_),
    .B(_0972_),
    .Y(_0988_)
  );
  \$_OR_  _1377_ (
    .A(_0988_),
    .B(_0967_),
    .Y(reg_src[10])
  );
  \$_AND_  _1378_ (
    .A(_0915_),
    .B(pc[11]),
    .Y(_0989_)
  );
  \$_AND_  _1379_ (
    .A(_0917_),
    .B(r1[11]),
    .Y(_0990_)
  );
  \$_OR_  _1380_ (
    .A(_0990_),
    .B(_0989_),
    .Y(_0991_)
  );
  \$_AND_  _1381_ (
    .A(_0920_),
    .B(r3[11]),
    .Y(_0992_)
  );
  \$_AND_  _1382_ (
    .A(_0922_),
    .B(r4[11]),
    .Y(_0993_)
  );
  \$_OR_  _1383_ (
    .A(_0993_),
    .B(_0992_),
    .Y(_0994_)
  );
  \$_OR_  _1384_ (
    .A(_0994_),
    .B(_0991_),
    .Y(_0995_)
  );
  \$_OR_  _1385_ (
    .A(_0995_),
    .B(_0959_),
    .Y(_0996_)
  );
  \$_AND_  _1386_ (
    .A(_0927_),
    .B(r15[11]),
    .Y(_0997_)
  );
  \$_AND_  _1387_ (
    .A(_0929_),
    .B(r13[11]),
    .Y(_0998_)
  );
  \$_AND_  _1388_ (
    .A(_0931_),
    .B(r14[11]),
    .Y(_0999_)
  );
  \$_OR_  _1389_ (
    .A(_0999_),
    .B(_0998_),
    .Y(_1000_)
  );
  \$_OR_  _1390_ (
    .A(_1000_),
    .B(_0997_),
    .Y(_1001_)
  );
  \$_AND_  _1391_ (
    .A(_0935_),
    .B(r9[11]),
    .Y(_1002_)
  );
  \$_AND_  _1392_ (
    .A(_0937_),
    .B(r10[11]),
    .Y(_1003_)
  );
  \$_OR_  _1393_ (
    .A(_1003_),
    .B(_1002_),
    .Y(_1004_)
  );
  \$_AND_  _1394_ (
    .A(_0940_),
    .B(r11[11]),
    .Y(_1005_)
  );
  \$_AND_  _1395_ (
    .A(_0942_),
    .B(r12[11]),
    .Y(_1006_)
  );
  \$_OR_  _1396_ (
    .A(_1006_),
    .B(_1005_),
    .Y(_1007_)
  );
  \$_OR_  _1397_ (
    .A(_1007_),
    .B(_1004_),
    .Y(_1008_)
  );
  \$_AND_  _1398_ (
    .A(_0946_),
    .B(r5[11]),
    .Y(_1009_)
  );
  \$_AND_  _1399_ (
    .A(_0948_),
    .B(r6[11]),
    .Y(_1010_)
  );
  \$_OR_  _1400_ (
    .A(_1010_),
    .B(_1009_),
    .Y(_1011_)
  );
  \$_AND_  _1401_ (
    .A(_0951_),
    .B(r7[11]),
    .Y(_1012_)
  );
  \$_AND_  _1402_ (
    .A(_0953_),
    .B(r8[11]),
    .Y(_1013_)
  );
  \$_OR_  _1403_ (
    .A(_1013_),
    .B(_1012_),
    .Y(_1014_)
  );
  \$_OR_  _1404_ (
    .A(_1014_),
    .B(_1011_),
    .Y(_1015_)
  );
  \$_OR_  _1405_ (
    .A(_1015_),
    .B(_1008_),
    .Y(_1016_)
  );
  \$_OR_  _1406_ (
    .A(_1016_),
    .B(_1001_),
    .Y(_1017_)
  );
  \$_OR_  _1407_ (
    .A(_1017_),
    .B(_0996_),
    .Y(reg_src[11])
  );
  \$_AND_  _1408_ (
    .A(_0915_),
    .B(pc[12]),
    .Y(_1018_)
  );
  \$_AND_  _1409_ (
    .A(_0917_),
    .B(r1[12]),
    .Y(_1019_)
  );
  \$_OR_  _1410_ (
    .A(_1019_),
    .B(_1018_),
    .Y(_1020_)
  );
  \$_AND_  _1411_ (
    .A(_0920_),
    .B(r3[12]),
    .Y(_1021_)
  );
  \$_AND_  _1412_ (
    .A(_0922_),
    .B(r4[12]),
    .Y(_1022_)
  );
  \$_OR_  _1413_ (
    .A(_1022_),
    .B(_1021_),
    .Y(_1023_)
  );
  \$_OR_  _1414_ (
    .A(_1023_),
    .B(_1020_),
    .Y(_1024_)
  );
  \$_OR_  _1415_ (
    .A(_1024_),
    .B(_0959_),
    .Y(_1025_)
  );
  \$_AND_  _1416_ (
    .A(_0927_),
    .B(r15[12]),
    .Y(_1026_)
  );
  \$_AND_  _1417_ (
    .A(_0929_),
    .B(r13[12]),
    .Y(_1027_)
  );
  \$_AND_  _1418_ (
    .A(_0931_),
    .B(r14[12]),
    .Y(_1028_)
  );
  \$_OR_  _1419_ (
    .A(_1028_),
    .B(_1027_),
    .Y(_1029_)
  );
  \$_OR_  _1420_ (
    .A(_1029_),
    .B(_1026_),
    .Y(_1030_)
  );
  \$_AND_  _1421_ (
    .A(_0935_),
    .B(r9[12]),
    .Y(_1031_)
  );
  \$_AND_  _1422_ (
    .A(_0937_),
    .B(r10[12]),
    .Y(_1032_)
  );
  \$_OR_  _1423_ (
    .A(_1032_),
    .B(_1031_),
    .Y(_1033_)
  );
  \$_AND_  _1424_ (
    .A(_0940_),
    .B(r11[12]),
    .Y(_1034_)
  );
  \$_AND_  _1425_ (
    .A(_0942_),
    .B(r12[12]),
    .Y(_1035_)
  );
  \$_OR_  _1426_ (
    .A(_1035_),
    .B(_1034_),
    .Y(_1036_)
  );
  \$_OR_  _1427_ (
    .A(_1036_),
    .B(_1033_),
    .Y(_1037_)
  );
  \$_AND_  _1428_ (
    .A(_0946_),
    .B(r5[12]),
    .Y(_1038_)
  );
  \$_AND_  _1429_ (
    .A(_0948_),
    .B(r6[12]),
    .Y(_1039_)
  );
  \$_OR_  _1430_ (
    .A(_1039_),
    .B(_1038_),
    .Y(_1040_)
  );
  \$_AND_  _1431_ (
    .A(_0951_),
    .B(r7[12]),
    .Y(_1041_)
  );
  \$_AND_  _1432_ (
    .A(_0953_),
    .B(r8[12]),
    .Y(_1042_)
  );
  \$_OR_  _1433_ (
    .A(_1042_),
    .B(_1041_),
    .Y(_1043_)
  );
  \$_OR_  _1434_ (
    .A(_1043_),
    .B(_1040_),
    .Y(_1044_)
  );
  \$_OR_  _1435_ (
    .A(_1044_),
    .B(_1037_),
    .Y(_1045_)
  );
  \$_OR_  _1436_ (
    .A(_1045_),
    .B(_1030_),
    .Y(_1046_)
  );
  \$_OR_  _1437_ (
    .A(_1046_),
    .B(_1025_),
    .Y(reg_src[12])
  );
  \$_AND_  _1438_ (
    .A(_0915_),
    .B(pc[13]),
    .Y(_1047_)
  );
  \$_AND_  _1439_ (
    .A(_0917_),
    .B(r1[13]),
    .Y(_1048_)
  );
  \$_OR_  _1440_ (
    .A(_1048_),
    .B(_1047_),
    .Y(_1049_)
  );
  \$_AND_  _1441_ (
    .A(_0920_),
    .B(r3[13]),
    .Y(_1050_)
  );
  \$_AND_  _1442_ (
    .A(_0922_),
    .B(r4[13]),
    .Y(_1051_)
  );
  \$_OR_  _1443_ (
    .A(_1051_),
    .B(_1050_),
    .Y(_1052_)
  );
  \$_OR_  _1444_ (
    .A(_1052_),
    .B(_1049_),
    .Y(_1053_)
  );
  \$_OR_  _1445_ (
    .A(_1053_),
    .B(_0959_),
    .Y(_1054_)
  );
  \$_AND_  _1446_ (
    .A(_0927_),
    .B(r15[13]),
    .Y(_1055_)
  );
  \$_AND_  _1447_ (
    .A(_0929_),
    .B(r13[13]),
    .Y(_1056_)
  );
  \$_AND_  _1448_ (
    .A(_0931_),
    .B(r14[13]),
    .Y(_1057_)
  );
  \$_OR_  _1449_ (
    .A(_1057_),
    .B(_1056_),
    .Y(_1058_)
  );
  \$_OR_  _1450_ (
    .A(_1058_),
    .B(_1055_),
    .Y(_1059_)
  );
  \$_AND_  _1451_ (
    .A(_0935_),
    .B(r9[13]),
    .Y(_1060_)
  );
  \$_AND_  _1452_ (
    .A(_0937_),
    .B(r10[13]),
    .Y(_1061_)
  );
  \$_OR_  _1453_ (
    .A(_1061_),
    .B(_1060_),
    .Y(_1062_)
  );
  \$_AND_  _1454_ (
    .A(_0940_),
    .B(r11[13]),
    .Y(_1063_)
  );
  \$_AND_  _1455_ (
    .A(_0942_),
    .B(r12[13]),
    .Y(_1064_)
  );
  \$_OR_  _1456_ (
    .A(_1064_),
    .B(_1063_),
    .Y(_1065_)
  );
  \$_OR_  _1457_ (
    .A(_1065_),
    .B(_1062_),
    .Y(_1066_)
  );
  \$_AND_  _1458_ (
    .A(_0946_),
    .B(r5[13]),
    .Y(_1067_)
  );
  \$_AND_  _1459_ (
    .A(_0948_),
    .B(r6[13]),
    .Y(_1068_)
  );
  \$_OR_  _1460_ (
    .A(_1068_),
    .B(_1067_),
    .Y(_1069_)
  );
  \$_AND_  _1461_ (
    .A(_0951_),
    .B(r7[13]),
    .Y(_1070_)
  );
  \$_AND_  _1462_ (
    .A(_0953_),
    .B(r8[13]),
    .Y(_1071_)
  );
  \$_OR_  _1463_ (
    .A(_1071_),
    .B(_1070_),
    .Y(_1072_)
  );
  \$_OR_  _1464_ (
    .A(_1072_),
    .B(_1069_),
    .Y(_1073_)
  );
  \$_OR_  _1465_ (
    .A(_1073_),
    .B(_1066_),
    .Y(_1074_)
  );
  \$_OR_  _1466_ (
    .A(_1074_),
    .B(_1059_),
    .Y(_1075_)
  );
  \$_OR_  _1467_ (
    .A(_1075_),
    .B(_1054_),
    .Y(reg_src[13])
  );
  \$_AND_  _1468_ (
    .A(_0915_),
    .B(pc[14]),
    .Y(_1076_)
  );
  \$_AND_  _1469_ (
    .A(_0917_),
    .B(r1[14]),
    .Y(_1077_)
  );
  \$_OR_  _1470_ (
    .A(_1077_),
    .B(_1076_),
    .Y(_1078_)
  );
  \$_AND_  _1471_ (
    .A(_0920_),
    .B(r3[14]),
    .Y(_1079_)
  );
  \$_AND_  _1472_ (
    .A(_0922_),
    .B(r4[14]),
    .Y(_1080_)
  );
  \$_OR_  _1473_ (
    .A(_1080_),
    .B(_1079_),
    .Y(_1081_)
  );
  \$_OR_  _1474_ (
    .A(_1081_),
    .B(_1078_),
    .Y(_1082_)
  );
  \$_OR_  _1475_ (
    .A(_1082_),
    .B(_0959_),
    .Y(_1083_)
  );
  \$_AND_  _1476_ (
    .A(_0927_),
    .B(r15[14]),
    .Y(_1084_)
  );
  \$_AND_  _1477_ (
    .A(_0929_),
    .B(r13[14]),
    .Y(_1085_)
  );
  \$_AND_  _1478_ (
    .A(_0931_),
    .B(r14[14]),
    .Y(_1086_)
  );
  \$_OR_  _1479_ (
    .A(_1086_),
    .B(_1085_),
    .Y(_1087_)
  );
  \$_OR_  _1480_ (
    .A(_1087_),
    .B(_1084_),
    .Y(_1088_)
  );
  \$_AND_  _1481_ (
    .A(_0935_),
    .B(r9[14]),
    .Y(_1089_)
  );
  \$_AND_  _1482_ (
    .A(_0937_),
    .B(r10[14]),
    .Y(_1090_)
  );
  \$_OR_  _1483_ (
    .A(_1090_),
    .B(_1089_),
    .Y(_1091_)
  );
  \$_AND_  _1484_ (
    .A(_0940_),
    .B(r11[14]),
    .Y(_1092_)
  );
  \$_AND_  _1485_ (
    .A(_0942_),
    .B(r12[14]),
    .Y(_1093_)
  );
  \$_OR_  _1486_ (
    .A(_1093_),
    .B(_1092_),
    .Y(_1094_)
  );
  \$_OR_  _1487_ (
    .A(_1094_),
    .B(_1091_),
    .Y(_1095_)
  );
  \$_AND_  _1488_ (
    .A(_0946_),
    .B(r5[14]),
    .Y(_1096_)
  );
  \$_AND_  _1489_ (
    .A(_0948_),
    .B(r6[14]),
    .Y(_1097_)
  );
  \$_OR_  _1490_ (
    .A(_1097_),
    .B(_1096_),
    .Y(_1098_)
  );
  \$_AND_  _1491_ (
    .A(_0951_),
    .B(r7[14]),
    .Y(_1099_)
  );
  \$_AND_  _1492_ (
    .A(_0953_),
    .B(r8[14]),
    .Y(_1100_)
  );
  \$_OR_  _1493_ (
    .A(_1100_),
    .B(_1099_),
    .Y(_1101_)
  );
  \$_OR_  _1494_ (
    .A(_1101_),
    .B(_1098_),
    .Y(_1102_)
  );
  \$_OR_  _1495_ (
    .A(_1102_),
    .B(_1095_),
    .Y(_1103_)
  );
  \$_OR_  _1496_ (
    .A(_1103_),
    .B(_1088_),
    .Y(_1104_)
  );
  \$_OR_  _1497_ (
    .A(_1104_),
    .B(_1083_),
    .Y(reg_src[14])
  );
  \$_AND_  _1498_ (
    .A(_0915_),
    .B(pc[15]),
    .Y(_1105_)
  );
  \$_AND_  _1499_ (
    .A(_0917_),
    .B(r1[15]),
    .Y(_1106_)
  );
  \$_OR_  _1500_ (
    .A(_1106_),
    .B(_1105_),
    .Y(_1107_)
  );
  \$_AND_  _1501_ (
    .A(_0920_),
    .B(r3[15]),
    .Y(_1108_)
  );
  \$_AND_  _1502_ (
    .A(_0922_),
    .B(r4[15]),
    .Y(_1109_)
  );
  \$_OR_  _1503_ (
    .A(_1109_),
    .B(_1108_),
    .Y(_1110_)
  );
  \$_OR_  _1504_ (
    .A(_1110_),
    .B(_1107_),
    .Y(_1111_)
  );
  \$_OR_  _1505_ (
    .A(_1111_),
    .B(_0959_),
    .Y(_1112_)
  );
  \$_AND_  _1506_ (
    .A(_0927_),
    .B(r15[15]),
    .Y(_1113_)
  );
  \$_AND_  _1507_ (
    .A(_0929_),
    .B(r13[15]),
    .Y(_1114_)
  );
  \$_AND_  _1508_ (
    .A(_0931_),
    .B(r14[15]),
    .Y(_1115_)
  );
  \$_OR_  _1509_ (
    .A(_1115_),
    .B(_1114_),
    .Y(_1116_)
  );
  \$_OR_  _1510_ (
    .A(_1116_),
    .B(_1113_),
    .Y(_1117_)
  );
  \$_AND_  _1511_ (
    .A(_0935_),
    .B(r9[15]),
    .Y(_1118_)
  );
  \$_AND_  _1512_ (
    .A(_0937_),
    .B(r10[15]),
    .Y(_1119_)
  );
  \$_OR_  _1513_ (
    .A(_1119_),
    .B(_1118_),
    .Y(_1120_)
  );
  \$_AND_  _1514_ (
    .A(_0940_),
    .B(r11[15]),
    .Y(_1121_)
  );
  \$_AND_  _1515_ (
    .A(_0942_),
    .B(r12[15]),
    .Y(_1122_)
  );
  \$_OR_  _1516_ (
    .A(_1122_),
    .B(_1121_),
    .Y(_1123_)
  );
  \$_OR_  _1517_ (
    .A(_1123_),
    .B(_1120_),
    .Y(_1124_)
  );
  \$_AND_  _1518_ (
    .A(_0946_),
    .B(r5[15]),
    .Y(_1125_)
  );
  \$_AND_  _1519_ (
    .A(_0948_),
    .B(r6[15]),
    .Y(_1126_)
  );
  \$_OR_  _1520_ (
    .A(_1126_),
    .B(_1125_),
    .Y(_1127_)
  );
  \$_AND_  _1521_ (
    .A(_0951_),
    .B(r7[15]),
    .Y(_1128_)
  );
  \$_AND_  _1522_ (
    .A(_0953_),
    .B(r8[15]),
    .Y(_1129_)
  );
  \$_OR_  _1523_ (
    .A(_1129_),
    .B(_1128_),
    .Y(_1130_)
  );
  \$_OR_  _1524_ (
    .A(_1130_),
    .B(_1127_),
    .Y(_1131_)
  );
  \$_OR_  _1525_ (
    .A(_1131_),
    .B(_1124_),
    .Y(_1132_)
  );
  \$_OR_  _1526_ (
    .A(_1132_),
    .B(_1117_),
    .Y(_1133_)
  );
  \$_OR_  _1527_ (
    .A(_1133_),
    .B(_1112_),
    .Y(reg_src[15])
  );
  \$_AND_  _1528_ (
    .A(_0912_),
    .B(r2[1]),
    .Y(_1134_)
  );
  \$_AND_  _1529_ (
    .A(_0915_),
    .B(pc[1]),
    .Y(_1135_)
  );
  \$_AND_  _1530_ (
    .A(_0917_),
    .B(r1[1]),
    .Y(_1136_)
  );
  \$_OR_  _1531_ (
    .A(_1136_),
    .B(_1135_),
    .Y(_1137_)
  );
  \$_AND_  _1532_ (
    .A(_0920_),
    .B(r3[1]),
    .Y(_1138_)
  );
  \$_AND_  _1533_ (
    .A(_0922_),
    .B(r4[1]),
    .Y(_1139_)
  );
  \$_OR_  _1534_ (
    .A(_1139_),
    .B(_1138_),
    .Y(_1140_)
  );
  \$_OR_  _1535_ (
    .A(_1140_),
    .B(_1137_),
    .Y(_1141_)
  );
  \$_OR_  _1536_ (
    .A(_1141_),
    .B(_1134_),
    .Y(_1142_)
  );
  \$_AND_  _1537_ (
    .A(_0927_),
    .B(r15[1]),
    .Y(_1143_)
  );
  \$_AND_  _1538_ (
    .A(_0929_),
    .B(r13[1]),
    .Y(_1144_)
  );
  \$_AND_  _1539_ (
    .A(_0931_),
    .B(r14[1]),
    .Y(_1145_)
  );
  \$_OR_  _1540_ (
    .A(_1145_),
    .B(_1144_),
    .Y(_1146_)
  );
  \$_OR_  _1541_ (
    .A(_1146_),
    .B(_1143_),
    .Y(_1147_)
  );
  \$_AND_  _1542_ (
    .A(_0935_),
    .B(r9[1]),
    .Y(_1148_)
  );
  \$_AND_  _1543_ (
    .A(_0937_),
    .B(r10[1]),
    .Y(_1149_)
  );
  \$_OR_  _1544_ (
    .A(_1149_),
    .B(_1148_),
    .Y(_1150_)
  );
  \$_AND_  _1545_ (
    .A(_0940_),
    .B(r11[1]),
    .Y(_1151_)
  );
  \$_AND_  _1546_ (
    .A(_0942_),
    .B(r12[1]),
    .Y(_1152_)
  );
  \$_OR_  _1547_ (
    .A(_1152_),
    .B(_1151_),
    .Y(_1153_)
  );
  \$_OR_  _1548_ (
    .A(_1153_),
    .B(_1150_),
    .Y(_1154_)
  );
  \$_AND_  _1549_ (
    .A(_0946_),
    .B(r5[1]),
    .Y(_1155_)
  );
  \$_AND_  _1550_ (
    .A(_0948_),
    .B(r6[1]),
    .Y(_1156_)
  );
  \$_OR_  _1551_ (
    .A(_1156_),
    .B(_1155_),
    .Y(_1157_)
  );
  \$_AND_  _1552_ (
    .A(_0951_),
    .B(r7[1]),
    .Y(_1158_)
  );
  \$_AND_  _1553_ (
    .A(_0953_),
    .B(r8[1]),
    .Y(_1159_)
  );
  \$_OR_  _1554_ (
    .A(_1159_),
    .B(_1158_),
    .Y(_1160_)
  );
  \$_OR_  _1555_ (
    .A(_1160_),
    .B(_1157_),
    .Y(_1161_)
  );
  \$_OR_  _1556_ (
    .A(_1161_),
    .B(_1154_),
    .Y(_1162_)
  );
  \$_OR_  _1557_ (
    .A(_1162_),
    .B(_1147_),
    .Y(_1163_)
  );
  \$_OR_  _1558_ (
    .A(_1163_),
    .B(_1142_),
    .Y(reg_src[1])
  );
  \$_AND_  _1559_ (
    .A(_0912_),
    .B(r2[2]),
    .Y(_1164_)
  );
  \$_AND_  _1560_ (
    .A(_0915_),
    .B(pc[2]),
    .Y(_1165_)
  );
  \$_AND_  _1561_ (
    .A(_0917_),
    .B(r1[2]),
    .Y(_1166_)
  );
  \$_OR_  _1562_ (
    .A(_1166_),
    .B(_1165_),
    .Y(_1167_)
  );
  \$_AND_  _1563_ (
    .A(_0920_),
    .B(r3[2]),
    .Y(_1168_)
  );
  \$_AND_  _1564_ (
    .A(_0922_),
    .B(r4[2]),
    .Y(_1169_)
  );
  \$_OR_  _1565_ (
    .A(_1169_),
    .B(_1168_),
    .Y(_1170_)
  );
  \$_OR_  _1566_ (
    .A(_1170_),
    .B(_1167_),
    .Y(_1171_)
  );
  \$_OR_  _1567_ (
    .A(_1171_),
    .B(_1164_),
    .Y(_1172_)
  );
  \$_AND_  _1568_ (
    .A(_0927_),
    .B(r15[2]),
    .Y(_1173_)
  );
  \$_AND_  _1569_ (
    .A(_0929_),
    .B(r13[2]),
    .Y(_1174_)
  );
  \$_AND_  _1570_ (
    .A(_0931_),
    .B(r14[2]),
    .Y(_1175_)
  );
  \$_OR_  _1571_ (
    .A(_1175_),
    .B(_1174_),
    .Y(_1176_)
  );
  \$_OR_  _1572_ (
    .A(_1176_),
    .B(_1173_),
    .Y(_1177_)
  );
  \$_AND_  _1573_ (
    .A(_0935_),
    .B(r9[2]),
    .Y(_1178_)
  );
  \$_AND_  _1574_ (
    .A(_0937_),
    .B(r10[2]),
    .Y(_1179_)
  );
  \$_OR_  _1575_ (
    .A(_1179_),
    .B(_1178_),
    .Y(_1180_)
  );
  \$_AND_  _1576_ (
    .A(_0940_),
    .B(r11[2]),
    .Y(_1181_)
  );
  \$_AND_  _1577_ (
    .A(_0942_),
    .B(r12[2]),
    .Y(_1182_)
  );
  \$_OR_  _1578_ (
    .A(_1182_),
    .B(_1181_),
    .Y(_1183_)
  );
  \$_OR_  _1579_ (
    .A(_1183_),
    .B(_1180_),
    .Y(_1184_)
  );
  \$_AND_  _1580_ (
    .A(_0946_),
    .B(r5[2]),
    .Y(_1185_)
  );
  \$_AND_  _1581_ (
    .A(_0948_),
    .B(r6[2]),
    .Y(_1186_)
  );
  \$_OR_  _1582_ (
    .A(_1186_),
    .B(_1185_),
    .Y(_1187_)
  );
  \$_AND_  _1583_ (
    .A(_0951_),
    .B(r7[2]),
    .Y(_1188_)
  );
  \$_AND_  _1584_ (
    .A(_0953_),
    .B(r8[2]),
    .Y(_1189_)
  );
  \$_OR_  _1585_ (
    .A(_1189_),
    .B(_1188_),
    .Y(_1190_)
  );
  \$_OR_  _1586_ (
    .A(_1190_),
    .B(_1187_),
    .Y(_1191_)
  );
  \$_OR_  _1587_ (
    .A(_1191_),
    .B(_1184_),
    .Y(_1192_)
  );
  \$_OR_  _1588_ (
    .A(_1192_),
    .B(_1177_),
    .Y(_1193_)
  );
  \$_OR_  _1589_ (
    .A(_1193_),
    .B(_1172_),
    .Y(reg_src[2])
  );
  \$_AND_  _1590_ (
    .A(_0912_),
    .B(gie),
    .Y(_1194_)
  );
  \$_AND_  _1591_ (
    .A(_0915_),
    .B(pc[3]),
    .Y(_1195_)
  );
  \$_AND_  _1592_ (
    .A(_0917_),
    .B(r1[3]),
    .Y(_1196_)
  );
  \$_OR_  _1593_ (
    .A(_1196_),
    .B(_1195_),
    .Y(_1197_)
  );
  \$_AND_  _1594_ (
    .A(_0920_),
    .B(r3[3]),
    .Y(_1198_)
  );
  \$_AND_  _1595_ (
    .A(_0922_),
    .B(r4[3]),
    .Y(_1199_)
  );
  \$_OR_  _1596_ (
    .A(_1199_),
    .B(_1198_),
    .Y(_1200_)
  );
  \$_OR_  _1597_ (
    .A(_1200_),
    .B(_1197_),
    .Y(_1201_)
  );
  \$_OR_  _1598_ (
    .A(_1201_),
    .B(_1194_),
    .Y(_1202_)
  );
  \$_AND_  _1599_ (
    .A(_0927_),
    .B(r15[3]),
    .Y(_1203_)
  );
  \$_AND_  _1600_ (
    .A(_0929_),
    .B(r13[3]),
    .Y(_1204_)
  );
  \$_AND_  _1601_ (
    .A(_0931_),
    .B(r14[3]),
    .Y(_1205_)
  );
  \$_OR_  _1602_ (
    .A(_1205_),
    .B(_1204_),
    .Y(_1206_)
  );
  \$_OR_  _1603_ (
    .A(_1206_),
    .B(_1203_),
    .Y(_1207_)
  );
  \$_AND_  _1604_ (
    .A(_0935_),
    .B(r9[3]),
    .Y(_1208_)
  );
  \$_AND_  _1605_ (
    .A(_0937_),
    .B(r10[3]),
    .Y(_1209_)
  );
  \$_OR_  _1606_ (
    .A(_1209_),
    .B(_1208_),
    .Y(_1210_)
  );
  \$_AND_  _1607_ (
    .A(_0940_),
    .B(r11[3]),
    .Y(_1211_)
  );
  \$_AND_  _1608_ (
    .A(_0942_),
    .B(r12[3]),
    .Y(_1212_)
  );
  \$_OR_  _1609_ (
    .A(_1212_),
    .B(_1211_),
    .Y(_1213_)
  );
  \$_OR_  _1610_ (
    .A(_1213_),
    .B(_1210_),
    .Y(_1214_)
  );
  \$_AND_  _1611_ (
    .A(_0946_),
    .B(r5[3]),
    .Y(_1215_)
  );
  \$_AND_  _1612_ (
    .A(_0948_),
    .B(r6[3]),
    .Y(_1216_)
  );
  \$_OR_  _1613_ (
    .A(_1216_),
    .B(_1215_),
    .Y(_1217_)
  );
  \$_AND_  _1614_ (
    .A(_0951_),
    .B(r7[3]),
    .Y(_1218_)
  );
  \$_AND_  _1615_ (
    .A(_0953_),
    .B(r8[3]),
    .Y(_1219_)
  );
  \$_OR_  _1616_ (
    .A(_1219_),
    .B(_1218_),
    .Y(_1220_)
  );
  \$_OR_  _1617_ (
    .A(_1220_),
    .B(_1217_),
    .Y(_1221_)
  );
  \$_OR_  _1618_ (
    .A(_1221_),
    .B(_1214_),
    .Y(_1222_)
  );
  \$_OR_  _1619_ (
    .A(_1222_),
    .B(_1207_),
    .Y(_1223_)
  );
  \$_OR_  _1620_ (
    .A(_1223_),
    .B(_1202_),
    .Y(reg_src[3])
  );
  \$_AND_  _1621_ (
    .A(_0912_),
    .B(r2[4]),
    .Y(_1224_)
  );
  \$_AND_  _1622_ (
    .A(_0915_),
    .B(pc[4]),
    .Y(_1225_)
  );
  \$_AND_  _1623_ (
    .A(_0917_),
    .B(r1[4]),
    .Y(_1226_)
  );
  \$_OR_  _1624_ (
    .A(_1226_),
    .B(_1225_),
    .Y(_1227_)
  );
  \$_AND_  _1625_ (
    .A(_0920_),
    .B(r3[4]),
    .Y(_1228_)
  );
  \$_AND_  _1626_ (
    .A(_0922_),
    .B(r4[4]),
    .Y(_1229_)
  );
  \$_OR_  _1627_ (
    .A(_1229_),
    .B(_1228_),
    .Y(_1230_)
  );
  \$_OR_  _1628_ (
    .A(_1230_),
    .B(_1227_),
    .Y(_1231_)
  );
  \$_OR_  _1629_ (
    .A(_1231_),
    .B(_1224_),
    .Y(_1232_)
  );
  \$_AND_  _1630_ (
    .A(_0927_),
    .B(r15[4]),
    .Y(_1233_)
  );
  \$_AND_  _1631_ (
    .A(_0929_),
    .B(r13[4]),
    .Y(_1234_)
  );
  \$_AND_  _1632_ (
    .A(_0931_),
    .B(r14[4]),
    .Y(_1235_)
  );
  \$_OR_  _1633_ (
    .A(_1235_),
    .B(_1234_),
    .Y(_1236_)
  );
  \$_OR_  _1634_ (
    .A(_1236_),
    .B(_1233_),
    .Y(_1237_)
  );
  \$_AND_  _1635_ (
    .A(_0935_),
    .B(r9[4]),
    .Y(_1238_)
  );
  \$_AND_  _1636_ (
    .A(_0937_),
    .B(r10[4]),
    .Y(_1239_)
  );
  \$_OR_  _1637_ (
    .A(_1239_),
    .B(_1238_),
    .Y(_1240_)
  );
  \$_AND_  _1638_ (
    .A(_0940_),
    .B(r11[4]),
    .Y(_1241_)
  );
  \$_AND_  _1639_ (
    .A(_0942_),
    .B(r12[4]),
    .Y(_1242_)
  );
  \$_OR_  _1640_ (
    .A(_1242_),
    .B(_1241_),
    .Y(_1243_)
  );
  \$_OR_  _1641_ (
    .A(_1243_),
    .B(_1240_),
    .Y(_1244_)
  );
  \$_AND_  _1642_ (
    .A(_0946_),
    .B(r5[4]),
    .Y(_1245_)
  );
  \$_AND_  _1643_ (
    .A(_0948_),
    .B(r6[4]),
    .Y(_1246_)
  );
  \$_OR_  _1644_ (
    .A(_1246_),
    .B(_1245_),
    .Y(_1247_)
  );
  \$_AND_  _1645_ (
    .A(_0951_),
    .B(r7[4]),
    .Y(_1248_)
  );
  \$_AND_  _1646_ (
    .A(_0953_),
    .B(r8[4]),
    .Y(_1249_)
  );
  \$_OR_  _1647_ (
    .A(_1249_),
    .B(_1248_),
    .Y(_1250_)
  );
  \$_OR_  _1648_ (
    .A(_1250_),
    .B(_1247_),
    .Y(_1251_)
  );
  \$_OR_  _1649_ (
    .A(_1251_),
    .B(_1244_),
    .Y(_1252_)
  );
  \$_OR_  _1650_ (
    .A(_1252_),
    .B(_1237_),
    .Y(_1253_)
  );
  \$_OR_  _1651_ (
    .A(_1253_),
    .B(_1232_),
    .Y(reg_src[4])
  );
  \$_AND_  _1652_ (
    .A(_0912_),
    .B(oscoff),
    .Y(_1254_)
  );
  \$_AND_  _1653_ (
    .A(_0915_),
    .B(pc[5]),
    .Y(_1255_)
  );
  \$_AND_  _1654_ (
    .A(_0917_),
    .B(r1[5]),
    .Y(_1256_)
  );
  \$_OR_  _1655_ (
    .A(_1256_),
    .B(_1255_),
    .Y(_1257_)
  );
  \$_AND_  _1656_ (
    .A(_0920_),
    .B(r3[5]),
    .Y(_1258_)
  );
  \$_AND_  _1657_ (
    .A(_0922_),
    .B(r4[5]),
    .Y(_1259_)
  );
  \$_OR_  _1658_ (
    .A(_1259_),
    .B(_1258_),
    .Y(_1260_)
  );
  \$_OR_  _1659_ (
    .A(_1260_),
    .B(_1257_),
    .Y(_1261_)
  );
  \$_OR_  _1660_ (
    .A(_1261_),
    .B(_1254_),
    .Y(_1262_)
  );
  \$_AND_  _1661_ (
    .A(_0927_),
    .B(r15[5]),
    .Y(_1263_)
  );
  \$_AND_  _1662_ (
    .A(_0929_),
    .B(r13[5]),
    .Y(_1264_)
  );
  \$_AND_  _1663_ (
    .A(_0931_),
    .B(r14[5]),
    .Y(_1265_)
  );
  \$_OR_  _1664_ (
    .A(_1265_),
    .B(_1264_),
    .Y(_1266_)
  );
  \$_OR_  _1665_ (
    .A(_1266_),
    .B(_1263_),
    .Y(_1267_)
  );
  \$_AND_  _1666_ (
    .A(_0935_),
    .B(r9[5]),
    .Y(_1268_)
  );
  \$_AND_  _1667_ (
    .A(_0937_),
    .B(r10[5]),
    .Y(_1269_)
  );
  \$_OR_  _1668_ (
    .A(_1269_),
    .B(_1268_),
    .Y(_1270_)
  );
  \$_AND_  _1669_ (
    .A(_0940_),
    .B(r11[5]),
    .Y(_1271_)
  );
  \$_AND_  _1670_ (
    .A(_0942_),
    .B(r12[5]),
    .Y(_1272_)
  );
  \$_OR_  _1671_ (
    .A(_1272_),
    .B(_1271_),
    .Y(_1273_)
  );
  \$_OR_  _1672_ (
    .A(_1273_),
    .B(_1270_),
    .Y(_1274_)
  );
  \$_AND_  _1673_ (
    .A(_0946_),
    .B(r5[5]),
    .Y(_1275_)
  );
  \$_AND_  _1674_ (
    .A(_0948_),
    .B(r6[5]),
    .Y(_1276_)
  );
  \$_OR_  _1675_ (
    .A(_1276_),
    .B(_1275_),
    .Y(_1277_)
  );
  \$_AND_  _1676_ (
    .A(_0951_),
    .B(r7[5]),
    .Y(_1278_)
  );
  \$_AND_  _1677_ (
    .A(_0953_),
    .B(r8[5]),
    .Y(_1279_)
  );
  \$_OR_  _1678_ (
    .A(_1279_),
    .B(_1278_),
    .Y(_1280_)
  );
  \$_OR_  _1679_ (
    .A(_1280_),
    .B(_1277_),
    .Y(_1281_)
  );
  \$_OR_  _1680_ (
    .A(_1281_),
    .B(_1274_),
    .Y(_1282_)
  );
  \$_OR_  _1681_ (
    .A(_1282_),
    .B(_1267_),
    .Y(_1283_)
  );
  \$_OR_  _1682_ (
    .A(_1283_),
    .B(_1262_),
    .Y(reg_src[5])
  );
  \$_AND_  _1683_ (
    .A(_0915_),
    .B(pc[6]),
    .Y(_1284_)
  );
  \$_AND_  _1684_ (
    .A(_0917_),
    .B(r1[6]),
    .Y(_1285_)
  );
  \$_OR_  _1685_ (
    .A(_1285_),
    .B(_1284_),
    .Y(_1286_)
  );
  \$_AND_  _1686_ (
    .A(_0920_),
    .B(r3[6]),
    .Y(_1287_)
  );
  \$_AND_  _1687_ (
    .A(_0922_),
    .B(r4[6]),
    .Y(_1288_)
  );
  \$_OR_  _1688_ (
    .A(_1288_),
    .B(_1287_),
    .Y(_1289_)
  );
  \$_OR_  _1689_ (
    .A(_1289_),
    .B(_1286_),
    .Y(_1290_)
  );
  \$_OR_  _1690_ (
    .A(_1290_),
    .B(_0959_),
    .Y(_1291_)
  );
  \$_AND_  _1691_ (
    .A(_0927_),
    .B(r15[6]),
    .Y(_1292_)
  );
  \$_AND_  _1692_ (
    .A(_0929_),
    .B(r13[6]),
    .Y(_1293_)
  );
  \$_AND_  _1693_ (
    .A(_0931_),
    .B(r14[6]),
    .Y(_1294_)
  );
  \$_OR_  _1694_ (
    .A(_1294_),
    .B(_1293_),
    .Y(_1295_)
  );
  \$_OR_  _1695_ (
    .A(_1295_),
    .B(_1292_),
    .Y(_1296_)
  );
  \$_AND_  _1696_ (
    .A(_0935_),
    .B(r9[6]),
    .Y(_1297_)
  );
  \$_AND_  _1697_ (
    .A(_0937_),
    .B(r10[6]),
    .Y(_1298_)
  );
  \$_OR_  _1698_ (
    .A(_1298_),
    .B(_1297_),
    .Y(_0015_)
  );
  \$_AND_  _1699_ (
    .A(_0940_),
    .B(r11[6]),
    .Y(_0016_)
  );
  \$_AND_  _1700_ (
    .A(_0942_),
    .B(r12[6]),
    .Y(_0017_)
  );
  \$_OR_  _1701_ (
    .A(_0017_),
    .B(_0016_),
    .Y(_0018_)
  );
  \$_OR_  _1702_ (
    .A(_0018_),
    .B(_0015_),
    .Y(_0019_)
  );
  \$_AND_  _1703_ (
    .A(_0946_),
    .B(r5[6]),
    .Y(_0020_)
  );
  \$_AND_  _1704_ (
    .A(_0948_),
    .B(r6[6]),
    .Y(_0021_)
  );
  \$_OR_  _1705_ (
    .A(_0021_),
    .B(_0020_),
    .Y(_0022_)
  );
  \$_AND_  _1706_ (
    .A(_0951_),
    .B(r7[6]),
    .Y(_0023_)
  );
  \$_AND_  _1707_ (
    .A(_0953_),
    .B(r8[6]),
    .Y(_0024_)
  );
  \$_OR_  _1708_ (
    .A(_0024_),
    .B(_0023_),
    .Y(_0025_)
  );
  \$_OR_  _1709_ (
    .A(_0025_),
    .B(_0022_),
    .Y(_0026_)
  );
  \$_OR_  _1710_ (
    .A(_0026_),
    .B(_0019_),
    .Y(_0027_)
  );
  \$_OR_  _1711_ (
    .A(_0027_),
    .B(_1296_),
    .Y(_0028_)
  );
  \$_OR_  _1712_ (
    .A(_0028_),
    .B(_1291_),
    .Y(reg_src[6])
  );
  \$_AND_  _1713_ (
    .A(_0912_),
    .B(r2[7]),
    .Y(_0029_)
  );
  \$_AND_  _1714_ (
    .A(_0915_),
    .B(pc[7]),
    .Y(_0030_)
  );
  \$_AND_  _1715_ (
    .A(_0917_),
    .B(r1[7]),
    .Y(_0031_)
  );
  \$_OR_  _1716_ (
    .A(_0031_),
    .B(_0030_),
    .Y(_0032_)
  );
  \$_AND_  _1717_ (
    .A(_0920_),
    .B(r3[7]),
    .Y(_0033_)
  );
  \$_AND_  _1718_ (
    .A(_0922_),
    .B(r4[7]),
    .Y(_0034_)
  );
  \$_OR_  _1719_ (
    .A(_0034_),
    .B(_0033_),
    .Y(_0035_)
  );
  \$_OR_  _1720_ (
    .A(_0035_),
    .B(_0032_),
    .Y(_0036_)
  );
  \$_OR_  _1721_ (
    .A(_0036_),
    .B(_0029_),
    .Y(_0037_)
  );
  \$_AND_  _1722_ (
    .A(_0927_),
    .B(r15[7]),
    .Y(_0038_)
  );
  \$_AND_  _1723_ (
    .A(_0929_),
    .B(r13[7]),
    .Y(_0039_)
  );
  \$_AND_  _1724_ (
    .A(_0931_),
    .B(r14[7]),
    .Y(_0040_)
  );
  \$_OR_  _1725_ (
    .A(_0040_),
    .B(_0039_),
    .Y(_0041_)
  );
  \$_OR_  _1726_ (
    .A(_0041_),
    .B(_0038_),
    .Y(_0042_)
  );
  \$_AND_  _1727_ (
    .A(_0935_),
    .B(r9[7]),
    .Y(_0043_)
  );
  \$_AND_  _1728_ (
    .A(_0937_),
    .B(r10[7]),
    .Y(_0044_)
  );
  \$_OR_  _1729_ (
    .A(_0044_),
    .B(_0043_),
    .Y(_0045_)
  );
  \$_AND_  _1730_ (
    .A(_0940_),
    .B(r11[7]),
    .Y(_0046_)
  );
  \$_AND_  _1731_ (
    .A(_0942_),
    .B(r12[7]),
    .Y(_0047_)
  );
  \$_OR_  _1732_ (
    .A(_0047_),
    .B(_0046_),
    .Y(_0048_)
  );
  \$_OR_  _1733_ (
    .A(_0048_),
    .B(_0045_),
    .Y(_0049_)
  );
  \$_AND_  _1734_ (
    .A(_0946_),
    .B(r5[7]),
    .Y(_0050_)
  );
  \$_AND_  _1735_ (
    .A(_0948_),
    .B(r6[7]),
    .Y(_0051_)
  );
  \$_OR_  _1736_ (
    .A(_0051_),
    .B(_0050_),
    .Y(_0052_)
  );
  \$_AND_  _1737_ (
    .A(_0951_),
    .B(r7[7]),
    .Y(_0053_)
  );
  \$_AND_  _1738_ (
    .A(_0953_),
    .B(r8[7]),
    .Y(_0054_)
  );
  \$_OR_  _1739_ (
    .A(_0054_),
    .B(_0053_),
    .Y(_0055_)
  );
  \$_OR_  _1740_ (
    .A(_0055_),
    .B(_0052_),
    .Y(_0056_)
  );
  \$_OR_  _1741_ (
    .A(_0056_),
    .B(_0049_),
    .Y(_0057_)
  );
  \$_OR_  _1742_ (
    .A(_0057_),
    .B(_0042_),
    .Y(_0058_)
  );
  \$_OR_  _1743_ (
    .A(_0058_),
    .B(_0037_),
    .Y(reg_src[7])
  );
  \$_AND_  _1744_ (
    .A(_0912_),
    .B(r2[8]),
    .Y(_0059_)
  );
  \$_AND_  _1745_ (
    .A(_0915_),
    .B(pc[8]),
    .Y(_0060_)
  );
  \$_AND_  _1746_ (
    .A(_0917_),
    .B(r1[8]),
    .Y(_0061_)
  );
  \$_OR_  _1747_ (
    .A(_0061_),
    .B(_0060_),
    .Y(_0062_)
  );
  \$_AND_  _1748_ (
    .A(_0920_),
    .B(r3[8]),
    .Y(_0063_)
  );
  \$_AND_  _1749_ (
    .A(_0922_),
    .B(r4[8]),
    .Y(_0064_)
  );
  \$_OR_  _1750_ (
    .A(_0064_),
    .B(_0063_),
    .Y(_0065_)
  );
  \$_OR_  _1751_ (
    .A(_0065_),
    .B(_0062_),
    .Y(_0066_)
  );
  \$_OR_  _1752_ (
    .A(_0066_),
    .B(_0059_),
    .Y(_0067_)
  );
  \$_AND_  _1753_ (
    .A(_0927_),
    .B(r15[8]),
    .Y(_0068_)
  );
  \$_AND_  _1754_ (
    .A(_0929_),
    .B(r13[8]),
    .Y(_0069_)
  );
  \$_AND_  _1755_ (
    .A(_0931_),
    .B(r14[8]),
    .Y(_0070_)
  );
  \$_OR_  _1756_ (
    .A(_0070_),
    .B(_0069_),
    .Y(_0071_)
  );
  \$_OR_  _1757_ (
    .A(_0071_),
    .B(_0068_),
    .Y(_0072_)
  );
  \$_AND_  _1758_ (
    .A(_0935_),
    .B(r9[8]),
    .Y(_0073_)
  );
  \$_AND_  _1759_ (
    .A(_0937_),
    .B(r10[8]),
    .Y(_0074_)
  );
  \$_OR_  _1760_ (
    .A(_0074_),
    .B(_0073_),
    .Y(_0075_)
  );
  \$_AND_  _1761_ (
    .A(_0940_),
    .B(r11[8]),
    .Y(_0076_)
  );
  \$_AND_  _1762_ (
    .A(_0942_),
    .B(r12[8]),
    .Y(_0077_)
  );
  \$_OR_  _1763_ (
    .A(_0077_),
    .B(_0076_),
    .Y(_0078_)
  );
  \$_OR_  _1764_ (
    .A(_0078_),
    .B(_0075_),
    .Y(_0079_)
  );
  \$_AND_  _1765_ (
    .A(_0946_),
    .B(r5[8]),
    .Y(_0080_)
  );
  \$_AND_  _1766_ (
    .A(_0948_),
    .B(r6[8]),
    .Y(_0081_)
  );
  \$_OR_  _1767_ (
    .A(_0081_),
    .B(_0080_),
    .Y(_0082_)
  );
  \$_AND_  _1768_ (
    .A(_0951_),
    .B(r7[8]),
    .Y(_0083_)
  );
  \$_AND_  _1769_ (
    .A(_0953_),
    .B(r8[8]),
    .Y(_0084_)
  );
  \$_OR_  _1770_ (
    .A(_0084_),
    .B(_0083_),
    .Y(_0085_)
  );
  \$_OR_  _1771_ (
    .A(_0085_),
    .B(_0082_),
    .Y(_0086_)
  );
  \$_OR_  _1772_ (
    .A(_0086_),
    .B(_0079_),
    .Y(_0087_)
  );
  \$_OR_  _1773_ (
    .A(_0087_),
    .B(_0072_),
    .Y(_0088_)
  );
  \$_OR_  _1774_ (
    .A(_0088_),
    .B(_0067_),
    .Y(reg_src[8])
  );
  \$_AND_  _1775_ (
    .A(_0915_),
    .B(pc[9]),
    .Y(_0089_)
  );
  \$_AND_  _1776_ (
    .A(_0917_),
    .B(r1[9]),
    .Y(_0090_)
  );
  \$_OR_  _1777_ (
    .A(_0090_),
    .B(_0089_),
    .Y(_0091_)
  );
  \$_AND_  _1778_ (
    .A(_0920_),
    .B(r3[9]),
    .Y(_0092_)
  );
  \$_AND_  _1779_ (
    .A(_0922_),
    .B(r4[9]),
    .Y(_0093_)
  );
  \$_OR_  _1780_ (
    .A(_0093_),
    .B(_0092_),
    .Y(_0094_)
  );
  \$_OR_  _1781_ (
    .A(_0094_),
    .B(_0091_),
    .Y(_0095_)
  );
  \$_OR_  _1782_ (
    .A(_0095_),
    .B(_0959_),
    .Y(_0096_)
  );
  \$_AND_  _1783_ (
    .A(_0927_),
    .B(r15[9]),
    .Y(_0097_)
  );
  \$_AND_  _1784_ (
    .A(_0929_),
    .B(r13[9]),
    .Y(_0098_)
  );
  \$_AND_  _1785_ (
    .A(_0931_),
    .B(r14[9]),
    .Y(_0099_)
  );
  \$_OR_  _1786_ (
    .A(_0099_),
    .B(_0098_),
    .Y(_0100_)
  );
  \$_OR_  _1787_ (
    .A(_0100_),
    .B(_0097_),
    .Y(_0101_)
  );
  \$_AND_  _1788_ (
    .A(_0935_),
    .B(r9[9]),
    .Y(_0102_)
  );
  \$_AND_  _1789_ (
    .A(_0937_),
    .B(r10[9]),
    .Y(_0103_)
  );
  \$_OR_  _1790_ (
    .A(_0103_),
    .B(_0102_),
    .Y(_0104_)
  );
  \$_AND_  _1791_ (
    .A(_0940_),
    .B(r11[9]),
    .Y(_0105_)
  );
  \$_AND_  _1792_ (
    .A(_0942_),
    .B(r12[9]),
    .Y(_0106_)
  );
  \$_OR_  _1793_ (
    .A(_0106_),
    .B(_0105_),
    .Y(_0107_)
  );
  \$_OR_  _1794_ (
    .A(_0107_),
    .B(_0104_),
    .Y(_0108_)
  );
  \$_AND_  _1795_ (
    .A(_0946_),
    .B(r5[9]),
    .Y(_0109_)
  );
  \$_AND_  _1796_ (
    .A(_0948_),
    .B(r6[9]),
    .Y(_0110_)
  );
  \$_OR_  _1797_ (
    .A(_0110_),
    .B(_0109_),
    .Y(_0111_)
  );
  \$_AND_  _1798_ (
    .A(_0951_),
    .B(r7[9]),
    .Y(_0112_)
  );
  \$_AND_  _1799_ (
    .A(_0953_),
    .B(r8[9]),
    .Y(_0113_)
  );
  \$_OR_  _1800_ (
    .A(_0113_),
    .B(_0112_),
    .Y(_0114_)
  );
  \$_OR_  _1801_ (
    .A(_0114_),
    .B(_0111_),
    .Y(_0115_)
  );
  \$_OR_  _1802_ (
    .A(_0115_),
    .B(_0108_),
    .Y(_0116_)
  );
  \$_OR_  _1803_ (
    .A(_0116_),
    .B(_0101_),
    .Y(_0117_)
  );
  \$_OR_  _1804_ (
    .A(_0117_),
    .B(_0096_),
    .Y(reg_src[9])
  );
  \$_AND_  _1805_ (
    .A(inst_dest[0]),
    .B(reg_dest_wr),
    .Y(_0118_)
  );
  \$_OR_  _1806_ (
    .A(_0118_),
    .B(reg_pc_call),
    .Y(pc_sw_wr)
  );
  \$_AND_  _1807_ (
    .A(inst_dest[2]),
    .B(reg_dest_wr),
    .Y(_0119_)
  );
  \$_OR_  _1808_ (
    .A(_0119_),
    .B(reg_sr_wr),
    .Y(_0120_)
  );
  \$_MUX_  _1809_ (
    .A(r2[4]),
    .B(reg_dest_val[4]),
    .S(_0120_),
    .Y(_0121_)
  );
  \$_AND_  _1810_ (
    .A(_0121_),
    .B(_0120_),
    .Y(_0122_)
  );
  \$_OR_  _1811_ (
    .A(_0122_),
    .B(r2[4]),
    .Y(cpuoff)
  );
  \$_AND_  _1812_ (
    .A(r4[0]),
    .B(inst_dest[4]),
    .Y(_0123_)
  );
  \$_AND_  _1813_ (
    .A(r5[0]),
    .B(inst_dest[5]),
    .Y(_0124_)
  );
  \$_OR_  _1814_ (
    .A(_0124_),
    .B(_0123_),
    .Y(_0125_)
  );
  \$_AND_  _1815_ (
    .A(r6[0]),
    .B(inst_dest[6]),
    .Y(_0126_)
  );
  \$_AND_  _1816_ (
    .A(r7[0]),
    .B(inst_dest[7]),
    .Y(_0127_)
  );
  \$_OR_  _1817_ (
    .A(_0127_),
    .B(_0126_),
    .Y(_0128_)
  );
  \$_OR_  _1818_ (
    .A(_0128_),
    .B(_0125_),
    .Y(_0129_)
  );
  \$_AND_  _1819_ (
    .A(pc[0]),
    .B(inst_dest[0]),
    .Y(_0130_)
  );
  \$_AND_  _1820_ (
    .A(r1[0]),
    .B(inst_dest[1]),
    .Y(_0131_)
  );
  \$_OR_  _1821_ (
    .A(_0131_),
    .B(_0130_),
    .Y(_0132_)
  );
  \$_AND_  _1822_ (
    .A(r2[0]),
    .B(inst_dest[2]),
    .Y(_0133_)
  );
  \$_AND_  _1823_ (
    .A(r3[0]),
    .B(inst_dest[3]),
    .Y(_0134_)
  );
  \$_OR_  _1824_ (
    .A(_0134_),
    .B(_0133_),
    .Y(_0135_)
  );
  \$_OR_  _1825_ (
    .A(_0135_),
    .B(_0132_),
    .Y(_0136_)
  );
  \$_OR_  _1826_ (
    .A(_0136_),
    .B(_0129_),
    .Y(_0137_)
  );
  \$_AND_  _1827_ (
    .A(r12[0]),
    .B(inst_dest[12]),
    .Y(_0138_)
  );
  \$_AND_  _1828_ (
    .A(r13[0]),
    .B(inst_dest[13]),
    .Y(_0139_)
  );
  \$_OR_  _1829_ (
    .A(_0139_),
    .B(_0138_),
    .Y(_0140_)
  );
  \$_AND_  _1830_ (
    .A(r14[0]),
    .B(inst_dest[14]),
    .Y(_0141_)
  );
  \$_AND_  _1831_ (
    .A(r15[0]),
    .B(inst_dest[15]),
    .Y(_0142_)
  );
  \$_OR_  _1832_ (
    .A(_0142_),
    .B(_0141_),
    .Y(_0143_)
  );
  \$_OR_  _1833_ (
    .A(_0143_),
    .B(_0140_),
    .Y(_0144_)
  );
  \$_AND_  _1834_ (
    .A(r8[0]),
    .B(inst_dest[8]),
    .Y(_0145_)
  );
  \$_AND_  _1835_ (
    .A(r9[0]),
    .B(inst_dest[9]),
    .Y(_0146_)
  );
  \$_OR_  _1836_ (
    .A(_0146_),
    .B(_0145_),
    .Y(_0147_)
  );
  \$_AND_  _1837_ (
    .A(r10[0]),
    .B(inst_dest[10]),
    .Y(_0148_)
  );
  \$_AND_  _1838_ (
    .A(r11[0]),
    .B(inst_dest[11]),
    .Y(_0149_)
  );
  \$_OR_  _1839_ (
    .A(_0149_),
    .B(_0148_),
    .Y(_0150_)
  );
  \$_OR_  _1840_ (
    .A(_0150_),
    .B(_0147_),
    .Y(_0151_)
  );
  \$_OR_  _1841_ (
    .A(_0151_),
    .B(_0144_),
    .Y(_0152_)
  );
  \$_OR_  _1842_ (
    .A(_0152_),
    .B(_0137_),
    .Y(reg_dest[0])
  );
  \$_AND_  _1843_ (
    .A(r4[10]),
    .B(inst_dest[4]),
    .Y(_0153_)
  );
  \$_AND_  _1844_ (
    .A(r5[10]),
    .B(inst_dest[5]),
    .Y(_0154_)
  );
  \$_OR_  _1845_ (
    .A(_0154_),
    .B(_0153_),
    .Y(_0155_)
  );
  \$_AND_  _1846_ (
    .A(r6[10]),
    .B(inst_dest[6]),
    .Y(_0156_)
  );
  \$_AND_  _1847_ (
    .A(r7[10]),
    .B(inst_dest[7]),
    .Y(_0157_)
  );
  \$_OR_  _1848_ (
    .A(_0157_),
    .B(_0156_),
    .Y(_0158_)
  );
  \$_OR_  _1849_ (
    .A(_0158_),
    .B(_0155_),
    .Y(_0159_)
  );
  \$_AND_  _1850_ (
    .A(pc[10]),
    .B(inst_dest[0]),
    .Y(_0160_)
  );
  \$_AND_  _1851_ (
    .A(r1[10]),
    .B(inst_dest[1]),
    .Y(_0161_)
  );
  \$_OR_  _1852_ (
    .A(_0161_),
    .B(_0160_),
    .Y(_0162_)
  );
  \$_AND_  _1853_ (
    .A(r2[15]),
    .B(inst_dest[2]),
    .Y(_0163_)
  );
  \$_AND_  _1854_ (
    .A(r3[10]),
    .B(inst_dest[3]),
    .Y(_0164_)
  );
  \$_OR_  _1855_ (
    .A(_0164_),
    .B(_0163_),
    .Y(_0165_)
  );
  \$_OR_  _1856_ (
    .A(_0165_),
    .B(_0162_),
    .Y(_0166_)
  );
  \$_OR_  _1857_ (
    .A(_0166_),
    .B(_0159_),
    .Y(_0167_)
  );
  \$_AND_  _1858_ (
    .A(r12[10]),
    .B(inst_dest[12]),
    .Y(_0168_)
  );
  \$_AND_  _1859_ (
    .A(r13[10]),
    .B(inst_dest[13]),
    .Y(_0169_)
  );
  \$_OR_  _1860_ (
    .A(_0169_),
    .B(_0168_),
    .Y(_0170_)
  );
  \$_AND_  _1861_ (
    .A(r14[10]),
    .B(inst_dest[14]),
    .Y(_0171_)
  );
  \$_AND_  _1862_ (
    .A(r15[10]),
    .B(inst_dest[15]),
    .Y(_0172_)
  );
  \$_OR_  _1863_ (
    .A(_0172_),
    .B(_0171_),
    .Y(_0173_)
  );
  \$_OR_  _1864_ (
    .A(_0173_),
    .B(_0170_),
    .Y(_0174_)
  );
  \$_AND_  _1865_ (
    .A(r8[10]),
    .B(inst_dest[8]),
    .Y(_0175_)
  );
  \$_AND_  _1866_ (
    .A(r9[10]),
    .B(inst_dest[9]),
    .Y(_0176_)
  );
  \$_OR_  _1867_ (
    .A(_0176_),
    .B(_0175_),
    .Y(_0177_)
  );
  \$_AND_  _1868_ (
    .A(r10[10]),
    .B(inst_dest[10]),
    .Y(_0178_)
  );
  \$_AND_  _1869_ (
    .A(r11[10]),
    .B(inst_dest[11]),
    .Y(_0179_)
  );
  \$_OR_  _1870_ (
    .A(_0179_),
    .B(_0178_),
    .Y(_0180_)
  );
  \$_OR_  _1871_ (
    .A(_0180_),
    .B(_0177_),
    .Y(_0181_)
  );
  \$_OR_  _1872_ (
    .A(_0181_),
    .B(_0174_),
    .Y(_0182_)
  );
  \$_OR_  _1873_ (
    .A(_0182_),
    .B(_0167_),
    .Y(reg_dest[10])
  );
  \$_AND_  _1874_ (
    .A(r4[11]),
    .B(inst_dest[4]),
    .Y(_0183_)
  );
  \$_AND_  _1875_ (
    .A(r5[11]),
    .B(inst_dest[5]),
    .Y(_0184_)
  );
  \$_OR_  _1876_ (
    .A(_0184_),
    .B(_0183_),
    .Y(_0185_)
  );
  \$_AND_  _1877_ (
    .A(r6[11]),
    .B(inst_dest[6]),
    .Y(_0186_)
  );
  \$_AND_  _1878_ (
    .A(r7[11]),
    .B(inst_dest[7]),
    .Y(_0187_)
  );
  \$_OR_  _1879_ (
    .A(_0187_),
    .B(_0186_),
    .Y(_0188_)
  );
  \$_OR_  _1880_ (
    .A(_0188_),
    .B(_0185_),
    .Y(_0189_)
  );
  \$_AND_  _1881_ (
    .A(pc[11]),
    .B(inst_dest[0]),
    .Y(_0190_)
  );
  \$_OR_  _1882_ (
    .A(_0190_),
    .B(_0163_),
    .Y(_0191_)
  );
  \$_AND_  _1883_ (
    .A(r1[11]),
    .B(inst_dest[1]),
    .Y(_0192_)
  );
  \$_AND_  _1884_ (
    .A(r3[11]),
    .B(inst_dest[3]),
    .Y(_0193_)
  );
  \$_OR_  _1885_ (
    .A(_0193_),
    .B(_0192_),
    .Y(_0194_)
  );
  \$_OR_  _1886_ (
    .A(_0194_),
    .B(_0191_),
    .Y(_0195_)
  );
  \$_OR_  _1887_ (
    .A(_0195_),
    .B(_0189_),
    .Y(_0196_)
  );
  \$_AND_  _1888_ (
    .A(r12[11]),
    .B(inst_dest[12]),
    .Y(_0197_)
  );
  \$_AND_  _1889_ (
    .A(r13[11]),
    .B(inst_dest[13]),
    .Y(_0198_)
  );
  \$_OR_  _1890_ (
    .A(_0198_),
    .B(_0197_),
    .Y(_0199_)
  );
  \$_AND_  _1891_ (
    .A(r14[11]),
    .B(inst_dest[14]),
    .Y(_0200_)
  );
  \$_AND_  _1892_ (
    .A(r15[11]),
    .B(inst_dest[15]),
    .Y(_0201_)
  );
  \$_OR_  _1893_ (
    .A(_0201_),
    .B(_0200_),
    .Y(_0202_)
  );
  \$_OR_  _1894_ (
    .A(_0202_),
    .B(_0199_),
    .Y(_0203_)
  );
  \$_AND_  _1895_ (
    .A(r8[11]),
    .B(inst_dest[8]),
    .Y(_0204_)
  );
  \$_AND_  _1896_ (
    .A(r9[11]),
    .B(inst_dest[9]),
    .Y(_0205_)
  );
  \$_OR_  _1897_ (
    .A(_0205_),
    .B(_0204_),
    .Y(_0206_)
  );
  \$_AND_  _1898_ (
    .A(r10[11]),
    .B(inst_dest[10]),
    .Y(_0207_)
  );
  \$_AND_  _1899_ (
    .A(r11[11]),
    .B(inst_dest[11]),
    .Y(_0208_)
  );
  \$_OR_  _1900_ (
    .A(_0208_),
    .B(_0207_),
    .Y(_0209_)
  );
  \$_OR_  _1901_ (
    .A(_0209_),
    .B(_0206_),
    .Y(_0210_)
  );
  \$_OR_  _1902_ (
    .A(_0210_),
    .B(_0203_),
    .Y(_0211_)
  );
  \$_OR_  _1903_ (
    .A(_0211_),
    .B(_0196_),
    .Y(reg_dest[11])
  );
  \$_AND_  _1904_ (
    .A(r4[12]),
    .B(inst_dest[4]),
    .Y(_0212_)
  );
  \$_AND_  _1905_ (
    .A(r5[12]),
    .B(inst_dest[5]),
    .Y(_0213_)
  );
  \$_OR_  _1906_ (
    .A(_0213_),
    .B(_0212_),
    .Y(_0214_)
  );
  \$_AND_  _1907_ (
    .A(r6[12]),
    .B(inst_dest[6]),
    .Y(_0215_)
  );
  \$_AND_  _1908_ (
    .A(r7[12]),
    .B(inst_dest[7]),
    .Y(_0216_)
  );
  \$_OR_  _1909_ (
    .A(_0216_),
    .B(_0215_),
    .Y(_0217_)
  );
  \$_OR_  _1910_ (
    .A(_0217_),
    .B(_0214_),
    .Y(_0218_)
  );
  \$_AND_  _1911_ (
    .A(pc[12]),
    .B(inst_dest[0]),
    .Y(_0219_)
  );
  \$_OR_  _1912_ (
    .A(_0219_),
    .B(_0163_),
    .Y(_0220_)
  );
  \$_AND_  _1913_ (
    .A(r1[12]),
    .B(inst_dest[1]),
    .Y(_0221_)
  );
  \$_AND_  _1914_ (
    .A(r3[12]),
    .B(inst_dest[3]),
    .Y(_0222_)
  );
  \$_OR_  _1915_ (
    .A(_0222_),
    .B(_0221_),
    .Y(_0223_)
  );
  \$_OR_  _1916_ (
    .A(_0223_),
    .B(_0220_),
    .Y(_0224_)
  );
  \$_OR_  _1917_ (
    .A(_0224_),
    .B(_0218_),
    .Y(_0225_)
  );
  \$_AND_  _1918_ (
    .A(r12[12]),
    .B(inst_dest[12]),
    .Y(_0226_)
  );
  \$_AND_  _1919_ (
    .A(r13[12]),
    .B(inst_dest[13]),
    .Y(_0227_)
  );
  \$_OR_  _1920_ (
    .A(_0227_),
    .B(_0226_),
    .Y(_0228_)
  );
  \$_AND_  _1921_ (
    .A(r14[12]),
    .B(inst_dest[14]),
    .Y(_0229_)
  );
  \$_AND_  _1922_ (
    .A(r15[12]),
    .B(inst_dest[15]),
    .Y(_0230_)
  );
  \$_OR_  _1923_ (
    .A(_0230_),
    .B(_0229_),
    .Y(_0231_)
  );
  \$_OR_  _1924_ (
    .A(_0231_),
    .B(_0228_),
    .Y(_0232_)
  );
  \$_AND_  _1925_ (
    .A(r8[12]),
    .B(inst_dest[8]),
    .Y(_0233_)
  );
  \$_AND_  _1926_ (
    .A(r9[12]),
    .B(inst_dest[9]),
    .Y(_0234_)
  );
  \$_OR_  _1927_ (
    .A(_0234_),
    .B(_0233_),
    .Y(_0235_)
  );
  \$_AND_  _1928_ (
    .A(r10[12]),
    .B(inst_dest[10]),
    .Y(_0236_)
  );
  \$_AND_  _1929_ (
    .A(r11[12]),
    .B(inst_dest[11]),
    .Y(_0237_)
  );
  \$_OR_  _1930_ (
    .A(_0237_),
    .B(_0236_),
    .Y(_0238_)
  );
  \$_OR_  _1931_ (
    .A(_0238_),
    .B(_0235_),
    .Y(_0239_)
  );
  \$_OR_  _1932_ (
    .A(_0239_),
    .B(_0232_),
    .Y(_0240_)
  );
  \$_OR_  _1933_ (
    .A(_0240_),
    .B(_0225_),
    .Y(reg_dest[12])
  );
  \$_AND_  _1934_ (
    .A(r4[13]),
    .B(inst_dest[4]),
    .Y(_0241_)
  );
  \$_AND_  _1935_ (
    .A(r5[13]),
    .B(inst_dest[5]),
    .Y(_0242_)
  );
  \$_OR_  _1936_ (
    .A(_0242_),
    .B(_0241_),
    .Y(_0243_)
  );
  \$_AND_  _1937_ (
    .A(r6[13]),
    .B(inst_dest[6]),
    .Y(_0244_)
  );
  \$_AND_  _1938_ (
    .A(r7[13]),
    .B(inst_dest[7]),
    .Y(_0245_)
  );
  \$_OR_  _1939_ (
    .A(_0245_),
    .B(_0244_),
    .Y(_0246_)
  );
  \$_OR_  _1940_ (
    .A(_0246_),
    .B(_0243_),
    .Y(_0247_)
  );
  \$_AND_  _1941_ (
    .A(pc[13]),
    .B(inst_dest[0]),
    .Y(_0248_)
  );
  \$_OR_  _1942_ (
    .A(_0248_),
    .B(_0163_),
    .Y(_0249_)
  );
  \$_AND_  _1943_ (
    .A(r1[13]),
    .B(inst_dest[1]),
    .Y(_0250_)
  );
  \$_AND_  _1944_ (
    .A(r3[13]),
    .B(inst_dest[3]),
    .Y(_0251_)
  );
  \$_OR_  _1945_ (
    .A(_0251_),
    .B(_0250_),
    .Y(_0252_)
  );
  \$_OR_  _1946_ (
    .A(_0252_),
    .B(_0249_),
    .Y(_0253_)
  );
  \$_OR_  _1947_ (
    .A(_0253_),
    .B(_0247_),
    .Y(_0254_)
  );
  \$_AND_  _1948_ (
    .A(r12[13]),
    .B(inst_dest[12]),
    .Y(_0255_)
  );
  \$_AND_  _1949_ (
    .A(r13[13]),
    .B(inst_dest[13]),
    .Y(_0256_)
  );
  \$_OR_  _1950_ (
    .A(_0256_),
    .B(_0255_),
    .Y(_0257_)
  );
  \$_AND_  _1951_ (
    .A(r14[13]),
    .B(inst_dest[14]),
    .Y(_0258_)
  );
  \$_AND_  _1952_ (
    .A(r15[13]),
    .B(inst_dest[15]),
    .Y(_0259_)
  );
  \$_OR_  _1953_ (
    .A(_0259_),
    .B(_0258_),
    .Y(_0260_)
  );
  \$_OR_  _1954_ (
    .A(_0260_),
    .B(_0257_),
    .Y(_0261_)
  );
  \$_AND_  _1955_ (
    .A(r8[13]),
    .B(inst_dest[8]),
    .Y(_0262_)
  );
  \$_AND_  _1956_ (
    .A(r9[13]),
    .B(inst_dest[9]),
    .Y(_0263_)
  );
  \$_OR_  _1957_ (
    .A(_0263_),
    .B(_0262_),
    .Y(_0264_)
  );
  \$_AND_  _1958_ (
    .A(r10[13]),
    .B(inst_dest[10]),
    .Y(_0265_)
  );
  \$_AND_  _1959_ (
    .A(r11[13]),
    .B(inst_dest[11]),
    .Y(_0266_)
  );
  \$_OR_  _1960_ (
    .A(_0266_),
    .B(_0265_),
    .Y(_0267_)
  );
  \$_OR_  _1961_ (
    .A(_0267_),
    .B(_0264_),
    .Y(_0268_)
  );
  \$_OR_  _1962_ (
    .A(_0268_),
    .B(_0261_),
    .Y(_0269_)
  );
  \$_OR_  _1963_ (
    .A(_0269_),
    .B(_0254_),
    .Y(reg_dest[13])
  );
  \$_AND_  _1964_ (
    .A(r4[14]),
    .B(inst_dest[4]),
    .Y(_0270_)
  );
  \$_AND_  _1965_ (
    .A(r5[14]),
    .B(inst_dest[5]),
    .Y(_0271_)
  );
  \$_OR_  _1966_ (
    .A(_0271_),
    .B(_0270_),
    .Y(_0272_)
  );
  \$_AND_  _1967_ (
    .A(r6[14]),
    .B(inst_dest[6]),
    .Y(_0273_)
  );
  \$_AND_  _1968_ (
    .A(r7[14]),
    .B(inst_dest[7]),
    .Y(_0274_)
  );
  \$_OR_  _1969_ (
    .A(_0274_),
    .B(_0273_),
    .Y(_0275_)
  );
  \$_OR_  _1970_ (
    .A(_0275_),
    .B(_0272_),
    .Y(_0276_)
  );
  \$_AND_  _1971_ (
    .A(pc[14]),
    .B(inst_dest[0]),
    .Y(_0277_)
  );
  \$_OR_  _1972_ (
    .A(_0277_),
    .B(_0163_),
    .Y(_0278_)
  );
  \$_AND_  _1973_ (
    .A(r1[14]),
    .B(inst_dest[1]),
    .Y(_0279_)
  );
  \$_AND_  _1974_ (
    .A(r3[14]),
    .B(inst_dest[3]),
    .Y(_0280_)
  );
  \$_OR_  _1975_ (
    .A(_0280_),
    .B(_0279_),
    .Y(_0281_)
  );
  \$_OR_  _1976_ (
    .A(_0281_),
    .B(_0278_),
    .Y(_0282_)
  );
  \$_OR_  _1977_ (
    .A(_0282_),
    .B(_0276_),
    .Y(_0283_)
  );
  \$_AND_  _1978_ (
    .A(r12[14]),
    .B(inst_dest[12]),
    .Y(_0284_)
  );
  \$_AND_  _1979_ (
    .A(r13[14]),
    .B(inst_dest[13]),
    .Y(_0285_)
  );
  \$_OR_  _1980_ (
    .A(_0285_),
    .B(_0284_),
    .Y(_0286_)
  );
  \$_AND_  _1981_ (
    .A(r14[14]),
    .B(inst_dest[14]),
    .Y(_0287_)
  );
  \$_AND_  _1982_ (
    .A(r15[14]),
    .B(inst_dest[15]),
    .Y(_0288_)
  );
  \$_OR_  _1983_ (
    .A(_0288_),
    .B(_0287_),
    .Y(_0289_)
  );
  \$_OR_  _1984_ (
    .A(_0289_),
    .B(_0286_),
    .Y(_0290_)
  );
  \$_AND_  _1985_ (
    .A(r8[14]),
    .B(inst_dest[8]),
    .Y(_0291_)
  );
  \$_AND_  _1986_ (
    .A(r9[14]),
    .B(inst_dest[9]),
    .Y(_0292_)
  );
  \$_OR_  _1987_ (
    .A(_0292_),
    .B(_0291_),
    .Y(_0293_)
  );
  \$_AND_  _1988_ (
    .A(r10[14]),
    .B(inst_dest[10]),
    .Y(_0294_)
  );
  \$_AND_  _1989_ (
    .A(r11[14]),
    .B(inst_dest[11]),
    .Y(_0295_)
  );
  \$_OR_  _1990_ (
    .A(_0295_),
    .B(_0294_),
    .Y(_0296_)
  );
  \$_OR_  _1991_ (
    .A(_0296_),
    .B(_0293_),
    .Y(_0297_)
  );
  \$_OR_  _1992_ (
    .A(_0297_),
    .B(_0290_),
    .Y(_0298_)
  );
  \$_OR_  _1993_ (
    .A(_0298_),
    .B(_0283_),
    .Y(reg_dest[14])
  );
  \$_AND_  _1994_ (
    .A(r4[15]),
    .B(inst_dest[4]),
    .Y(_0299_)
  );
  \$_AND_  _1995_ (
    .A(r5[15]),
    .B(inst_dest[5]),
    .Y(_0300_)
  );
  \$_OR_  _1996_ (
    .A(_0300_),
    .B(_0299_),
    .Y(_0301_)
  );
  \$_AND_  _1997_ (
    .A(r6[15]),
    .B(inst_dest[6]),
    .Y(_0302_)
  );
  \$_AND_  _1998_ (
    .A(r7[15]),
    .B(inst_dest[7]),
    .Y(_0303_)
  );
  \$_OR_  _1999_ (
    .A(_0303_),
    .B(_0302_),
    .Y(_0304_)
  );
  \$_OR_  _2000_ (
    .A(_0304_),
    .B(_0301_),
    .Y(_0305_)
  );
  \$_AND_  _2001_ (
    .A(pc[15]),
    .B(inst_dest[0]),
    .Y(_0306_)
  );
  \$_OR_  _2002_ (
    .A(_0306_),
    .B(_0163_),
    .Y(_0307_)
  );
  \$_AND_  _2003_ (
    .A(r1[15]),
    .B(inst_dest[1]),
    .Y(_0308_)
  );
  \$_AND_  _2004_ (
    .A(r3[15]),
    .B(inst_dest[3]),
    .Y(_0309_)
  );
  \$_OR_  _2005_ (
    .A(_0309_),
    .B(_0308_),
    .Y(_0310_)
  );
  \$_OR_  _2006_ (
    .A(_0310_),
    .B(_0307_),
    .Y(_0311_)
  );
  \$_OR_  _2007_ (
    .A(_0311_),
    .B(_0305_),
    .Y(_0312_)
  );
  \$_AND_  _2008_ (
    .A(r12[15]),
    .B(inst_dest[12]),
    .Y(_0313_)
  );
  \$_AND_  _2009_ (
    .A(r13[15]),
    .B(inst_dest[13]),
    .Y(_0314_)
  );
  \$_OR_  _2010_ (
    .A(_0314_),
    .B(_0313_),
    .Y(_0315_)
  );
  \$_AND_  _2011_ (
    .A(r14[15]),
    .B(inst_dest[14]),
    .Y(_0316_)
  );
  \$_AND_  _2012_ (
    .A(r15[15]),
    .B(inst_dest[15]),
    .Y(_0317_)
  );
  \$_OR_  _2013_ (
    .A(_0317_),
    .B(_0316_),
    .Y(_0318_)
  );
  \$_OR_  _2014_ (
    .A(_0318_),
    .B(_0315_),
    .Y(_0319_)
  );
  \$_AND_  _2015_ (
    .A(r8[15]),
    .B(inst_dest[8]),
    .Y(_0320_)
  );
  \$_AND_  _2016_ (
    .A(r9[15]),
    .B(inst_dest[9]),
    .Y(_0321_)
  );
  \$_OR_  _2017_ (
    .A(_0321_),
    .B(_0320_),
    .Y(_0322_)
  );
  \$_AND_  _2018_ (
    .A(r10[15]),
    .B(inst_dest[10]),
    .Y(_0323_)
  );
  \$_AND_  _2019_ (
    .A(r11[15]),
    .B(inst_dest[11]),
    .Y(_0324_)
  );
  \$_OR_  _2020_ (
    .A(_0324_),
    .B(_0323_),
    .Y(_0325_)
  );
  \$_OR_  _2021_ (
    .A(_0325_),
    .B(_0322_),
    .Y(_0326_)
  );
  \$_OR_  _2022_ (
    .A(_0326_),
    .B(_0319_),
    .Y(_0327_)
  );
  \$_OR_  _2023_ (
    .A(_0327_),
    .B(_0312_),
    .Y(reg_dest[15])
  );
  \$_AND_  _2024_ (
    .A(r4[1]),
    .B(inst_dest[4]),
    .Y(_0328_)
  );
  \$_AND_  _2025_ (
    .A(r5[1]),
    .B(inst_dest[5]),
    .Y(_0329_)
  );
  \$_OR_  _2026_ (
    .A(_0329_),
    .B(_0328_),
    .Y(_0330_)
  );
  \$_AND_  _2027_ (
    .A(r6[1]),
    .B(inst_dest[6]),
    .Y(_0331_)
  );
  \$_AND_  _2028_ (
    .A(r7[1]),
    .B(inst_dest[7]),
    .Y(_0332_)
  );
  \$_OR_  _2029_ (
    .A(_0332_),
    .B(_0331_),
    .Y(_0333_)
  );
  \$_OR_  _2030_ (
    .A(_0333_),
    .B(_0330_),
    .Y(_0334_)
  );
  \$_AND_  _2031_ (
    .A(pc[1]),
    .B(inst_dest[0]),
    .Y(_0335_)
  );
  \$_AND_  _2032_ (
    .A(r1[1]),
    .B(inst_dest[1]),
    .Y(_0336_)
  );
  \$_OR_  _2033_ (
    .A(_0336_),
    .B(_0335_),
    .Y(_0337_)
  );
  \$_AND_  _2034_ (
    .A(r2[1]),
    .B(inst_dest[2]),
    .Y(_0338_)
  );
  \$_AND_  _2035_ (
    .A(r3[1]),
    .B(inst_dest[3]),
    .Y(_0339_)
  );
  \$_OR_  _2036_ (
    .A(_0339_),
    .B(_0338_),
    .Y(_0340_)
  );
  \$_OR_  _2037_ (
    .A(_0340_),
    .B(_0337_),
    .Y(_0341_)
  );
  \$_OR_  _2038_ (
    .A(_0341_),
    .B(_0334_),
    .Y(_0342_)
  );
  \$_AND_  _2039_ (
    .A(r12[1]),
    .B(inst_dest[12]),
    .Y(_0343_)
  );
  \$_AND_  _2040_ (
    .A(r13[1]),
    .B(inst_dest[13]),
    .Y(_0344_)
  );
  \$_OR_  _2041_ (
    .A(_0344_),
    .B(_0343_),
    .Y(_0345_)
  );
  \$_AND_  _2042_ (
    .A(r14[1]),
    .B(inst_dest[14]),
    .Y(_0346_)
  );
  \$_AND_  _2043_ (
    .A(r15[1]),
    .B(inst_dest[15]),
    .Y(_0347_)
  );
  \$_OR_  _2044_ (
    .A(_0347_),
    .B(_0346_),
    .Y(_0348_)
  );
  \$_OR_  _2045_ (
    .A(_0348_),
    .B(_0345_),
    .Y(_0349_)
  );
  \$_AND_  _2046_ (
    .A(r8[1]),
    .B(inst_dest[8]),
    .Y(_0350_)
  );
  \$_AND_  _2047_ (
    .A(r9[1]),
    .B(inst_dest[9]),
    .Y(_0351_)
  );
  \$_OR_  _2048_ (
    .A(_0351_),
    .B(_0350_),
    .Y(_0352_)
  );
  \$_AND_  _2049_ (
    .A(r10[1]),
    .B(inst_dest[10]),
    .Y(_0353_)
  );
  \$_AND_  _2050_ (
    .A(r11[1]),
    .B(inst_dest[11]),
    .Y(_0354_)
  );
  \$_OR_  _2051_ (
    .A(_0354_),
    .B(_0353_),
    .Y(_0355_)
  );
  \$_OR_  _2052_ (
    .A(_0355_),
    .B(_0352_),
    .Y(_0356_)
  );
  \$_OR_  _2053_ (
    .A(_0356_),
    .B(_0349_),
    .Y(_0357_)
  );
  \$_OR_  _2054_ (
    .A(_0357_),
    .B(_0342_),
    .Y(reg_dest[1])
  );
  \$_AND_  _2055_ (
    .A(r4[2]),
    .B(inst_dest[4]),
    .Y(_0358_)
  );
  \$_AND_  _2056_ (
    .A(r5[2]),
    .B(inst_dest[5]),
    .Y(_0359_)
  );
  \$_OR_  _2057_ (
    .A(_0359_),
    .B(_0358_),
    .Y(_0360_)
  );
  \$_AND_  _2058_ (
    .A(r6[2]),
    .B(inst_dest[6]),
    .Y(_0361_)
  );
  \$_AND_  _2059_ (
    .A(r7[2]),
    .B(inst_dest[7]),
    .Y(_0362_)
  );
  \$_OR_  _2060_ (
    .A(_0362_),
    .B(_0361_),
    .Y(_0363_)
  );
  \$_OR_  _2061_ (
    .A(_0363_),
    .B(_0360_),
    .Y(_0364_)
  );
  \$_AND_  _2062_ (
    .A(pc[2]),
    .B(inst_dest[0]),
    .Y(_0365_)
  );
  \$_AND_  _2063_ (
    .A(r1[2]),
    .B(inst_dest[1]),
    .Y(_0366_)
  );
  \$_OR_  _2064_ (
    .A(_0366_),
    .B(_0365_),
    .Y(_0367_)
  );
  \$_AND_  _2065_ (
    .A(r2[2]),
    .B(inst_dest[2]),
    .Y(_0368_)
  );
  \$_AND_  _2066_ (
    .A(r3[2]),
    .B(inst_dest[3]),
    .Y(_0369_)
  );
  \$_OR_  _2067_ (
    .A(_0369_),
    .B(_0368_),
    .Y(_0370_)
  );
  \$_OR_  _2068_ (
    .A(_0370_),
    .B(_0367_),
    .Y(_0371_)
  );
  \$_OR_  _2069_ (
    .A(_0371_),
    .B(_0364_),
    .Y(_0372_)
  );
  \$_AND_  _2070_ (
    .A(r12[2]),
    .B(inst_dest[12]),
    .Y(_0373_)
  );
  \$_AND_  _2071_ (
    .A(r13[2]),
    .B(inst_dest[13]),
    .Y(_0374_)
  );
  \$_OR_  _2072_ (
    .A(_0374_),
    .B(_0373_),
    .Y(_0375_)
  );
  \$_AND_  _2073_ (
    .A(r14[2]),
    .B(inst_dest[14]),
    .Y(_0376_)
  );
  \$_AND_  _2074_ (
    .A(r15[2]),
    .B(inst_dest[15]),
    .Y(_0377_)
  );
  \$_OR_  _2075_ (
    .A(_0377_),
    .B(_0376_),
    .Y(_0378_)
  );
  \$_OR_  _2076_ (
    .A(_0378_),
    .B(_0375_),
    .Y(_0379_)
  );
  \$_AND_  _2077_ (
    .A(r8[2]),
    .B(inst_dest[8]),
    .Y(_0380_)
  );
  \$_AND_  _2078_ (
    .A(r9[2]),
    .B(inst_dest[9]),
    .Y(_0381_)
  );
  \$_OR_  _2079_ (
    .A(_0381_),
    .B(_0380_),
    .Y(_0382_)
  );
  \$_AND_  _2080_ (
    .A(r10[2]),
    .B(inst_dest[10]),
    .Y(_0383_)
  );
  \$_AND_  _2081_ (
    .A(r11[2]),
    .B(inst_dest[11]),
    .Y(_0384_)
  );
  \$_OR_  _2082_ (
    .A(_0384_),
    .B(_0383_),
    .Y(_0385_)
  );
  \$_OR_  _2083_ (
    .A(_0385_),
    .B(_0382_),
    .Y(_0386_)
  );
  \$_OR_  _2084_ (
    .A(_0386_),
    .B(_0379_),
    .Y(_0387_)
  );
  \$_OR_  _2085_ (
    .A(_0387_),
    .B(_0372_),
    .Y(reg_dest[2])
  );
  \$_AND_  _2086_ (
    .A(r4[3]),
    .B(inst_dest[4]),
    .Y(_0388_)
  );
  \$_AND_  _2087_ (
    .A(r5[3]),
    .B(inst_dest[5]),
    .Y(_0389_)
  );
  \$_OR_  _2088_ (
    .A(_0389_),
    .B(_0388_),
    .Y(_0390_)
  );
  \$_AND_  _2089_ (
    .A(r6[3]),
    .B(inst_dest[6]),
    .Y(_0391_)
  );
  \$_AND_  _2090_ (
    .A(r7[3]),
    .B(inst_dest[7]),
    .Y(_0392_)
  );
  \$_OR_  _2091_ (
    .A(_0392_),
    .B(_0391_),
    .Y(_0393_)
  );
  \$_OR_  _2092_ (
    .A(_0393_),
    .B(_0390_),
    .Y(_0394_)
  );
  \$_AND_  _2093_ (
    .A(pc[3]),
    .B(inst_dest[0]),
    .Y(_0395_)
  );
  \$_AND_  _2094_ (
    .A(r1[3]),
    .B(inst_dest[1]),
    .Y(_0396_)
  );
  \$_OR_  _2095_ (
    .A(_0396_),
    .B(_0395_),
    .Y(_0397_)
  );
  \$_AND_  _2096_ (
    .A(gie),
    .B(inst_dest[2]),
    .Y(_0398_)
  );
  \$_AND_  _2097_ (
    .A(r3[3]),
    .B(inst_dest[3]),
    .Y(_0399_)
  );
  \$_OR_  _2098_ (
    .A(_0399_),
    .B(_0398_),
    .Y(_0400_)
  );
  \$_OR_  _2099_ (
    .A(_0400_),
    .B(_0397_),
    .Y(_0401_)
  );
  \$_OR_  _2100_ (
    .A(_0401_),
    .B(_0394_),
    .Y(_0402_)
  );
  \$_AND_  _2101_ (
    .A(r12[3]),
    .B(inst_dest[12]),
    .Y(_0403_)
  );
  \$_AND_  _2102_ (
    .A(r13[3]),
    .B(inst_dest[13]),
    .Y(_0404_)
  );
  \$_OR_  _2103_ (
    .A(_0404_),
    .B(_0403_),
    .Y(_0405_)
  );
  \$_AND_  _2104_ (
    .A(r14[3]),
    .B(inst_dest[14]),
    .Y(_0406_)
  );
  \$_AND_  _2105_ (
    .A(r15[3]),
    .B(inst_dest[15]),
    .Y(_0407_)
  );
  \$_OR_  _2106_ (
    .A(_0407_),
    .B(_0406_),
    .Y(_0408_)
  );
  \$_OR_  _2107_ (
    .A(_0408_),
    .B(_0405_),
    .Y(_0409_)
  );
  \$_AND_  _2108_ (
    .A(r8[3]),
    .B(inst_dest[8]),
    .Y(_0410_)
  );
  \$_AND_  _2109_ (
    .A(r9[3]),
    .B(inst_dest[9]),
    .Y(_0411_)
  );
  \$_OR_  _2110_ (
    .A(_0411_),
    .B(_0410_),
    .Y(_0412_)
  );
  \$_AND_  _2111_ (
    .A(r10[3]),
    .B(inst_dest[10]),
    .Y(_0413_)
  );
  \$_AND_  _2112_ (
    .A(r11[3]),
    .B(inst_dest[11]),
    .Y(_0414_)
  );
  \$_OR_  _2113_ (
    .A(_0414_),
    .B(_0413_),
    .Y(_0415_)
  );
  \$_OR_  _2114_ (
    .A(_0415_),
    .B(_0412_),
    .Y(_0416_)
  );
  \$_OR_  _2115_ (
    .A(_0416_),
    .B(_0409_),
    .Y(_0417_)
  );
  \$_OR_  _2116_ (
    .A(_0417_),
    .B(_0402_),
    .Y(reg_dest[3])
  );
  \$_AND_  _2117_ (
    .A(r4[4]),
    .B(inst_dest[4]),
    .Y(_0418_)
  );
  \$_AND_  _2118_ (
    .A(r5[4]),
    .B(inst_dest[5]),
    .Y(_0419_)
  );
  \$_OR_  _2119_ (
    .A(_0419_),
    .B(_0418_),
    .Y(_0420_)
  );
  \$_AND_  _2120_ (
    .A(r6[4]),
    .B(inst_dest[6]),
    .Y(_0421_)
  );
  \$_AND_  _2121_ (
    .A(r7[4]),
    .B(inst_dest[7]),
    .Y(_0422_)
  );
  \$_OR_  _2122_ (
    .A(_0422_),
    .B(_0421_),
    .Y(_0423_)
  );
  \$_OR_  _2123_ (
    .A(_0423_),
    .B(_0420_),
    .Y(_0424_)
  );
  \$_AND_  _2124_ (
    .A(pc[4]),
    .B(inst_dest[0]),
    .Y(_0425_)
  );
  \$_AND_  _2125_ (
    .A(r1[4]),
    .B(inst_dest[1]),
    .Y(_0426_)
  );
  \$_OR_  _2126_ (
    .A(_0426_),
    .B(_0425_),
    .Y(_0427_)
  );
  \$_AND_  _2127_ (
    .A(r2[4]),
    .B(inst_dest[2]),
    .Y(_0428_)
  );
  \$_AND_  _2128_ (
    .A(r3[4]),
    .B(inst_dest[3]),
    .Y(_0429_)
  );
  \$_OR_  _2129_ (
    .A(_0429_),
    .B(_0428_),
    .Y(_0430_)
  );
  \$_OR_  _2130_ (
    .A(_0430_),
    .B(_0427_),
    .Y(_0431_)
  );
  \$_OR_  _2131_ (
    .A(_0431_),
    .B(_0424_),
    .Y(_0432_)
  );
  \$_AND_  _2132_ (
    .A(r12[4]),
    .B(inst_dest[12]),
    .Y(_0433_)
  );
  \$_AND_  _2133_ (
    .A(r13[4]),
    .B(inst_dest[13]),
    .Y(_0434_)
  );
  \$_OR_  _2134_ (
    .A(_0434_),
    .B(_0433_),
    .Y(_0435_)
  );
  \$_AND_  _2135_ (
    .A(r14[4]),
    .B(inst_dest[14]),
    .Y(_0436_)
  );
  \$_AND_  _2136_ (
    .A(r15[4]),
    .B(inst_dest[15]),
    .Y(_0437_)
  );
  \$_OR_  _2137_ (
    .A(_0437_),
    .B(_0436_),
    .Y(_0438_)
  );
  \$_OR_  _2138_ (
    .A(_0438_),
    .B(_0435_),
    .Y(_0439_)
  );
  \$_AND_  _2139_ (
    .A(r8[4]),
    .B(inst_dest[8]),
    .Y(_0440_)
  );
  \$_AND_  _2140_ (
    .A(r9[4]),
    .B(inst_dest[9]),
    .Y(_0441_)
  );
  \$_OR_  _2141_ (
    .A(_0441_),
    .B(_0440_),
    .Y(_0442_)
  );
  \$_AND_  _2142_ (
    .A(r10[4]),
    .B(inst_dest[10]),
    .Y(_0443_)
  );
  \$_AND_  _2143_ (
    .A(r11[4]),
    .B(inst_dest[11]),
    .Y(_0444_)
  );
  \$_OR_  _2144_ (
    .A(_0444_),
    .B(_0443_),
    .Y(_0445_)
  );
  \$_OR_  _2145_ (
    .A(_0445_),
    .B(_0442_),
    .Y(_0446_)
  );
  \$_OR_  _2146_ (
    .A(_0446_),
    .B(_0439_),
    .Y(_0447_)
  );
  \$_OR_  _2147_ (
    .A(_0447_),
    .B(_0432_),
    .Y(reg_dest[4])
  );
  \$_AND_  _2148_ (
    .A(r4[5]),
    .B(inst_dest[4]),
    .Y(_0448_)
  );
  \$_AND_  _2149_ (
    .A(r5[5]),
    .B(inst_dest[5]),
    .Y(_0449_)
  );
  \$_OR_  _2150_ (
    .A(_0449_),
    .B(_0448_),
    .Y(_0450_)
  );
  \$_AND_  _2151_ (
    .A(r6[5]),
    .B(inst_dest[6]),
    .Y(_0451_)
  );
  \$_AND_  _2152_ (
    .A(r7[5]),
    .B(inst_dest[7]),
    .Y(_0452_)
  );
  \$_OR_  _2153_ (
    .A(_0452_),
    .B(_0451_),
    .Y(_0453_)
  );
  \$_OR_  _2154_ (
    .A(_0453_),
    .B(_0450_),
    .Y(_0454_)
  );
  \$_AND_  _2155_ (
    .A(pc[5]),
    .B(inst_dest[0]),
    .Y(_0455_)
  );
  \$_AND_  _2156_ (
    .A(r1[5]),
    .B(inst_dest[1]),
    .Y(_0456_)
  );
  \$_OR_  _2157_ (
    .A(_0456_),
    .B(_0455_),
    .Y(_0457_)
  );
  \$_AND_  _2158_ (
    .A(oscoff),
    .B(inst_dest[2]),
    .Y(_0458_)
  );
  \$_AND_  _2159_ (
    .A(r3[5]),
    .B(inst_dest[3]),
    .Y(_0459_)
  );
  \$_OR_  _2160_ (
    .A(_0459_),
    .B(_0458_),
    .Y(_0460_)
  );
  \$_OR_  _2161_ (
    .A(_0460_),
    .B(_0457_),
    .Y(_0461_)
  );
  \$_OR_  _2162_ (
    .A(_0461_),
    .B(_0454_),
    .Y(_0462_)
  );
  \$_AND_  _2163_ (
    .A(r12[5]),
    .B(inst_dest[12]),
    .Y(_0463_)
  );
  \$_AND_  _2164_ (
    .A(r13[5]),
    .B(inst_dest[13]),
    .Y(_0464_)
  );
  \$_OR_  _2165_ (
    .A(_0464_),
    .B(_0463_),
    .Y(_0465_)
  );
  \$_AND_  _2166_ (
    .A(r14[5]),
    .B(inst_dest[14]),
    .Y(_0466_)
  );
  \$_AND_  _2167_ (
    .A(r15[5]),
    .B(inst_dest[15]),
    .Y(_0467_)
  );
  \$_OR_  _2168_ (
    .A(_0467_),
    .B(_0466_),
    .Y(_0468_)
  );
  \$_OR_  _2169_ (
    .A(_0468_),
    .B(_0465_),
    .Y(_0469_)
  );
  \$_AND_  _2170_ (
    .A(r8[5]),
    .B(inst_dest[8]),
    .Y(_0470_)
  );
  \$_AND_  _2171_ (
    .A(r9[5]),
    .B(inst_dest[9]),
    .Y(_0471_)
  );
  \$_OR_  _2172_ (
    .A(_0471_),
    .B(_0470_),
    .Y(_0472_)
  );
  \$_AND_  _2173_ (
    .A(r10[5]),
    .B(inst_dest[10]),
    .Y(_0473_)
  );
  \$_AND_  _2174_ (
    .A(r11[5]),
    .B(inst_dest[11]),
    .Y(_0474_)
  );
  \$_OR_  _2175_ (
    .A(_0474_),
    .B(_0473_),
    .Y(_0475_)
  );
  \$_OR_  _2176_ (
    .A(_0475_),
    .B(_0472_),
    .Y(_0476_)
  );
  \$_OR_  _2177_ (
    .A(_0476_),
    .B(_0469_),
    .Y(_0477_)
  );
  \$_OR_  _2178_ (
    .A(_0477_),
    .B(_0462_),
    .Y(reg_dest[5])
  );
  \$_AND_  _2179_ (
    .A(r4[6]),
    .B(inst_dest[4]),
    .Y(_0478_)
  );
  \$_AND_  _2180_ (
    .A(r5[6]),
    .B(inst_dest[5]),
    .Y(_0479_)
  );
  \$_OR_  _2181_ (
    .A(_0479_),
    .B(_0478_),
    .Y(_0480_)
  );
  \$_AND_  _2182_ (
    .A(r6[6]),
    .B(inst_dest[6]),
    .Y(_0481_)
  );
  \$_AND_  _2183_ (
    .A(r7[6]),
    .B(inst_dest[7]),
    .Y(_0482_)
  );
  \$_OR_  _2184_ (
    .A(_0482_),
    .B(_0481_),
    .Y(_0483_)
  );
  \$_OR_  _2185_ (
    .A(_0483_),
    .B(_0480_),
    .Y(_0484_)
  );
  \$_AND_  _2186_ (
    .A(pc[6]),
    .B(inst_dest[0]),
    .Y(_0485_)
  );
  \$_OR_  _2187_ (
    .A(_0485_),
    .B(_0163_),
    .Y(_0486_)
  );
  \$_AND_  _2188_ (
    .A(r1[6]),
    .B(inst_dest[1]),
    .Y(_0487_)
  );
  \$_AND_  _2189_ (
    .A(r3[6]),
    .B(inst_dest[3]),
    .Y(_0488_)
  );
  \$_OR_  _2190_ (
    .A(_0488_),
    .B(_0487_),
    .Y(_0489_)
  );
  \$_OR_  _2191_ (
    .A(_0489_),
    .B(_0486_),
    .Y(_0490_)
  );
  \$_OR_  _2192_ (
    .A(_0490_),
    .B(_0484_),
    .Y(_0491_)
  );
  \$_AND_  _2193_ (
    .A(r12[6]),
    .B(inst_dest[12]),
    .Y(_0492_)
  );
  \$_AND_  _2194_ (
    .A(r13[6]),
    .B(inst_dest[13]),
    .Y(_0493_)
  );
  \$_OR_  _2195_ (
    .A(_0493_),
    .B(_0492_),
    .Y(_0494_)
  );
  \$_AND_  _2196_ (
    .A(r14[6]),
    .B(inst_dest[14]),
    .Y(_0495_)
  );
  \$_AND_  _2197_ (
    .A(r15[6]),
    .B(inst_dest[15]),
    .Y(_0496_)
  );
  \$_OR_  _2198_ (
    .A(_0496_),
    .B(_0495_),
    .Y(_0497_)
  );
  \$_OR_  _2199_ (
    .A(_0497_),
    .B(_0494_),
    .Y(_0498_)
  );
  \$_AND_  _2200_ (
    .A(r8[6]),
    .B(inst_dest[8]),
    .Y(_0499_)
  );
  \$_AND_  _2201_ (
    .A(r9[6]),
    .B(inst_dest[9]),
    .Y(_0500_)
  );
  \$_OR_  _2202_ (
    .A(_0500_),
    .B(_0499_),
    .Y(_0501_)
  );
  \$_AND_  _2203_ (
    .A(r10[6]),
    .B(inst_dest[10]),
    .Y(_0502_)
  );
  \$_AND_  _2204_ (
    .A(r11[6]),
    .B(inst_dest[11]),
    .Y(_0503_)
  );
  \$_OR_  _2205_ (
    .A(_0503_),
    .B(_0502_),
    .Y(_0504_)
  );
  \$_OR_  _2206_ (
    .A(_0504_),
    .B(_0501_),
    .Y(_0505_)
  );
  \$_OR_  _2207_ (
    .A(_0505_),
    .B(_0498_),
    .Y(_0506_)
  );
  \$_OR_  _2208_ (
    .A(_0506_),
    .B(_0491_),
    .Y(reg_dest[6])
  );
  \$_AND_  _2209_ (
    .A(r4[7]),
    .B(inst_dest[4]),
    .Y(_0507_)
  );
  \$_AND_  _2210_ (
    .A(r5[7]),
    .B(inst_dest[5]),
    .Y(_0508_)
  );
  \$_OR_  _2211_ (
    .A(_0508_),
    .B(_0507_),
    .Y(_0509_)
  );
  \$_AND_  _2212_ (
    .A(r6[7]),
    .B(inst_dest[6]),
    .Y(_0510_)
  );
  \$_AND_  _2213_ (
    .A(r7[7]),
    .B(inst_dest[7]),
    .Y(_0511_)
  );
  \$_OR_  _2214_ (
    .A(_0511_),
    .B(_0510_),
    .Y(_0512_)
  );
  \$_OR_  _2215_ (
    .A(_0512_),
    .B(_0509_),
    .Y(_0513_)
  );
  \$_AND_  _2216_ (
    .A(pc[7]),
    .B(inst_dest[0]),
    .Y(_0514_)
  );
  \$_AND_  _2217_ (
    .A(r1[7]),
    .B(inst_dest[1]),
    .Y(_0515_)
  );
  \$_OR_  _2218_ (
    .A(_0515_),
    .B(_0514_),
    .Y(_0516_)
  );
  \$_AND_  _2219_ (
    .A(r2[7]),
    .B(inst_dest[2]),
    .Y(_0517_)
  );
  \$_AND_  _2220_ (
    .A(r3[7]),
    .B(inst_dest[3]),
    .Y(_0518_)
  );
  \$_OR_  _2221_ (
    .A(_0518_),
    .B(_0517_),
    .Y(_0519_)
  );
  \$_OR_  _2222_ (
    .A(_0519_),
    .B(_0516_),
    .Y(_0520_)
  );
  \$_OR_  _2223_ (
    .A(_0520_),
    .B(_0513_),
    .Y(_0521_)
  );
  \$_AND_  _2224_ (
    .A(r12[7]),
    .B(inst_dest[12]),
    .Y(_0522_)
  );
  \$_AND_  _2225_ (
    .A(r13[7]),
    .B(inst_dest[13]),
    .Y(_0523_)
  );
  \$_OR_  _2226_ (
    .A(_0523_),
    .B(_0522_),
    .Y(_0524_)
  );
  \$_AND_  _2227_ (
    .A(r14[7]),
    .B(inst_dest[14]),
    .Y(_0525_)
  );
  \$_AND_  _2228_ (
    .A(r15[7]),
    .B(inst_dest[15]),
    .Y(_0526_)
  );
  \$_OR_  _2229_ (
    .A(_0526_),
    .B(_0525_),
    .Y(_0527_)
  );
  \$_OR_  _2230_ (
    .A(_0527_),
    .B(_0524_),
    .Y(_0528_)
  );
  \$_AND_  _2231_ (
    .A(r8[7]),
    .B(inst_dest[8]),
    .Y(_0529_)
  );
  \$_AND_  _2232_ (
    .A(r9[7]),
    .B(inst_dest[9]),
    .Y(_0530_)
  );
  \$_OR_  _2233_ (
    .A(_0530_),
    .B(_0529_),
    .Y(_0531_)
  );
  \$_AND_  _2234_ (
    .A(r10[7]),
    .B(inst_dest[10]),
    .Y(_0532_)
  );
  \$_AND_  _2235_ (
    .A(r11[7]),
    .B(inst_dest[11]),
    .Y(_0533_)
  );
  \$_OR_  _2236_ (
    .A(_0533_),
    .B(_0532_),
    .Y(_0534_)
  );
  \$_OR_  _2237_ (
    .A(_0534_),
    .B(_0531_),
    .Y(_0535_)
  );
  \$_OR_  _2238_ (
    .A(_0535_),
    .B(_0528_),
    .Y(_0536_)
  );
  \$_OR_  _2239_ (
    .A(_0536_),
    .B(_0521_),
    .Y(reg_dest[7])
  );
  \$_AND_  _2240_ (
    .A(r4[8]),
    .B(inst_dest[4]),
    .Y(_0537_)
  );
  \$_AND_  _2241_ (
    .A(r5[8]),
    .B(inst_dest[5]),
    .Y(_0538_)
  );
  \$_OR_  _2242_ (
    .A(_0538_),
    .B(_0537_),
    .Y(_0539_)
  );
  \$_AND_  _2243_ (
    .A(r6[8]),
    .B(inst_dest[6]),
    .Y(_0540_)
  );
  \$_AND_  _2244_ (
    .A(r7[8]),
    .B(inst_dest[7]),
    .Y(_0541_)
  );
  \$_OR_  _2245_ (
    .A(_0541_),
    .B(_0540_),
    .Y(_0542_)
  );
  \$_OR_  _2246_ (
    .A(_0542_),
    .B(_0539_),
    .Y(_0543_)
  );
  \$_AND_  _2247_ (
    .A(pc[8]),
    .B(inst_dest[0]),
    .Y(_0544_)
  );
  \$_AND_  _2248_ (
    .A(r1[8]),
    .B(inst_dest[1]),
    .Y(_0545_)
  );
  \$_OR_  _2249_ (
    .A(_0545_),
    .B(_0544_),
    .Y(_0546_)
  );
  \$_AND_  _2250_ (
    .A(r2[8]),
    .B(inst_dest[2]),
    .Y(_0547_)
  );
  \$_AND_  _2251_ (
    .A(r3[8]),
    .B(inst_dest[3]),
    .Y(_0548_)
  );
  \$_OR_  _2252_ (
    .A(_0548_),
    .B(_0547_),
    .Y(_0549_)
  );
  \$_OR_  _2253_ (
    .A(_0549_),
    .B(_0546_),
    .Y(_0550_)
  );
  \$_OR_  _2254_ (
    .A(_0550_),
    .B(_0543_),
    .Y(_0551_)
  );
  \$_AND_  _2255_ (
    .A(r12[8]),
    .B(inst_dest[12]),
    .Y(_0552_)
  );
  \$_AND_  _2256_ (
    .A(r13[8]),
    .B(inst_dest[13]),
    .Y(_0553_)
  );
  \$_OR_  _2257_ (
    .A(_0553_),
    .B(_0552_),
    .Y(_0554_)
  );
  \$_AND_  _2258_ (
    .A(r14[8]),
    .B(inst_dest[14]),
    .Y(_0555_)
  );
  \$_AND_  _2259_ (
    .A(r15[8]),
    .B(inst_dest[15]),
    .Y(_0556_)
  );
  \$_OR_  _2260_ (
    .A(_0556_),
    .B(_0555_),
    .Y(_0557_)
  );
  \$_OR_  _2261_ (
    .A(_0557_),
    .B(_0554_),
    .Y(_0558_)
  );
  \$_AND_  _2262_ (
    .A(r8[8]),
    .B(inst_dest[8]),
    .Y(_0559_)
  );
  \$_AND_  _2263_ (
    .A(r9[8]),
    .B(inst_dest[9]),
    .Y(_0560_)
  );
  \$_OR_  _2264_ (
    .A(_0560_),
    .B(_0559_),
    .Y(_0561_)
  );
  \$_AND_  _2265_ (
    .A(r10[8]),
    .B(inst_dest[10]),
    .Y(_0562_)
  );
  \$_AND_  _2266_ (
    .A(r11[8]),
    .B(inst_dest[11]),
    .Y(_0563_)
  );
  \$_OR_  _2267_ (
    .A(_0563_),
    .B(_0562_),
    .Y(_0564_)
  );
  \$_OR_  _2268_ (
    .A(_0564_),
    .B(_0561_),
    .Y(_0565_)
  );
  \$_OR_  _2269_ (
    .A(_0565_),
    .B(_0558_),
    .Y(_0566_)
  );
  \$_OR_  _2270_ (
    .A(_0566_),
    .B(_0551_),
    .Y(reg_dest[8])
  );
  \$_AND_  _2271_ (
    .A(r4[9]),
    .B(inst_dest[4]),
    .Y(_0567_)
  );
  \$_AND_  _2272_ (
    .A(r5[9]),
    .B(inst_dest[5]),
    .Y(_0568_)
  );
  \$_OR_  _2273_ (
    .A(_0568_),
    .B(_0567_),
    .Y(_0569_)
  );
  \$_AND_  _2274_ (
    .A(r6[9]),
    .B(inst_dest[6]),
    .Y(_0570_)
  );
  \$_AND_  _2275_ (
    .A(r7[9]),
    .B(inst_dest[7]),
    .Y(_0571_)
  );
  \$_OR_  _2276_ (
    .A(_0571_),
    .B(_0570_),
    .Y(_0572_)
  );
  \$_OR_  _2277_ (
    .A(_0572_),
    .B(_0569_),
    .Y(_0573_)
  );
  \$_AND_  _2278_ (
    .A(pc[9]),
    .B(inst_dest[0]),
    .Y(_0574_)
  );
  \$_OR_  _2279_ (
    .A(_0574_),
    .B(_0163_),
    .Y(_0575_)
  );
  \$_AND_  _2280_ (
    .A(r1[9]),
    .B(inst_dest[1]),
    .Y(_0576_)
  );
  \$_AND_  _2281_ (
    .A(r3[9]),
    .B(inst_dest[3]),
    .Y(_0577_)
  );
  \$_OR_  _2282_ (
    .A(_0577_),
    .B(_0576_),
    .Y(_0578_)
  );
  \$_OR_  _2283_ (
    .A(_0578_),
    .B(_0575_),
    .Y(_0579_)
  );
  \$_OR_  _2284_ (
    .A(_0579_),
    .B(_0573_),
    .Y(_0580_)
  );
  \$_AND_  _2285_ (
    .A(r12[9]),
    .B(inst_dest[12]),
    .Y(_0581_)
  );
  \$_AND_  _2286_ (
    .A(r13[9]),
    .B(inst_dest[13]),
    .Y(_0582_)
  );
  \$_OR_  _2287_ (
    .A(_0582_),
    .B(_0581_),
    .Y(_0583_)
  );
  \$_AND_  _2288_ (
    .A(r14[9]),
    .B(inst_dest[14]),
    .Y(_0584_)
  );
  \$_AND_  _2289_ (
    .A(r15[9]),
    .B(inst_dest[15]),
    .Y(_0585_)
  );
  \$_OR_  _2290_ (
    .A(_0585_),
    .B(_0584_),
    .Y(_0586_)
  );
  \$_OR_  _2291_ (
    .A(_0586_),
    .B(_0583_),
    .Y(_0587_)
  );
  \$_AND_  _2292_ (
    .A(r8[9]),
    .B(inst_dest[8]),
    .Y(_0588_)
  );
  \$_AND_  _2293_ (
    .A(r9[9]),
    .B(inst_dest[9]),
    .Y(_0589_)
  );
  \$_OR_  _2294_ (
    .A(_0589_),
    .B(_0588_),
    .Y(_0590_)
  );
  \$_AND_  _2295_ (
    .A(r10[9]),
    .B(inst_dest[10]),
    .Y(_0591_)
  );
  \$_AND_  _2296_ (
    .A(r11[9]),
    .B(inst_dest[11]),
    .Y(_0592_)
  );
  \$_OR_  _2297_ (
    .A(_0592_),
    .B(_0591_),
    .Y(_0593_)
  );
  \$_OR_  _2298_ (
    .A(_0593_),
    .B(_0590_),
    .Y(_0594_)
  );
  \$_OR_  _2299_ (
    .A(_0594_),
    .B(_0587_),
    .Y(_0595_)
  );
  \$_OR_  _2300_ (
    .A(_0595_),
    .B(_0580_),
    .Y(reg_dest[9])
  );
  \$_INV_  _2301_ (
    .A(reg_incr),
    .Y(_0596_)
  );
  \$_INV_  _2302_ (
    .A(_0917_),
    .Y(_0597_)
  );
  \$_OR_  _2303_ (
    .A(_0597_),
    .B(_0596_),
    .Y(_0598_)
  );
  \$_AND_  _2304_ (
    .A(inst_dest[1]),
    .B(reg_dest_wr),
    .Y(_0599_)
  );
  \$_INV_  _2305_ (
    .A(_0599_),
    .Y(_0600_)
  );
  \$_INV_  _2306_ (
    .A(reg_sp_wr),
    .Y(_0601_)
  );
  \$_AND_  _2307_ (
    .A(_0601_),
    .B(r1[0]),
    .Y(_0602_)
  );
  \$_AND_  _2308_ (
    .A(_0602_),
    .B(_0600_),
    .Y(_0603_)
  );
  \$_AND_  _2309_ (
    .A(_0603_),
    .B(_0598_),
    .Y(_0006_[0])
  );
  \$_INV_  _2310_ (
    .A(inst_bw),
    .Y(_0604_)
  );
  \$_AND_  _2311_ (
    .A(reg_dest_val[10]),
    .B(_0604_),
    .Y(pc_sw[10])
  );
  \$_AND_  _2312_ (
    .A(_0597_),
    .B(inst_bw),
    .Y(_0605_)
  );
  \$_INV_  _2313_ (
    .A(_0605_),
    .Y(_0606_)
  );
  \$_AND_  _2314_ (
    .A(_0606_),
    .B(reg_src[1]),
    .Y(_0607_)
  );
  \$_XOR_  _2315_ (
    .A(_0606_),
    .B(reg_src[1]),
    .Y(_0608_)
  );
  \$_AND_  _2316_ (
    .A(_0605_),
    .B(reg_src[0]),
    .Y(_0609_)
  );
  \$_AND_  _2317_ (
    .A(_0609_),
    .B(_0608_),
    .Y(_0610_)
  );
  \$_OR_  _2318_ (
    .A(_0610_),
    .B(_0607_),
    .Y(_0611_)
  );
  \$_AND_  _2319_ (
    .A(_0611_),
    .B(reg_src[2]),
    .Y(_0612_)
  );
  \$_AND_  _2320_ (
    .A(_0612_),
    .B(reg_src[3]),
    .Y(_0613_)
  );
  \$_AND_  _2321_ (
    .A(_0613_),
    .B(reg_src[4]),
    .Y(_0614_)
  );
  \$_AND_  _2322_ (
    .A(_0614_),
    .B(reg_src[5]),
    .Y(_0615_)
  );
  \$_AND_  _2323_ (
    .A(_0615_),
    .B(reg_src[6]),
    .Y(_0616_)
  );
  \$_AND_  _2324_ (
    .A(_0616_),
    .B(reg_src[7]),
    .Y(_0617_)
  );
  \$_AND_  _2325_ (
    .A(_0617_),
    .B(reg_src[8]),
    .Y(_0618_)
  );
  \$_AND_  _2326_ (
    .A(_0618_),
    .B(reg_src[9]),
    .Y(_0619_)
  );
  \$_XOR_  _2327_ (
    .A(_0619_),
    .B(reg_src[10]),
    .Y(_0620_)
  );
  \$_MUX_  _2328_ (
    .A(_0620_),
    .B(r1[10]),
    .S(_0598_),
    .Y(_0621_)
  );
  \$_MUX_  _2329_ (
    .A(_0621_),
    .B(reg_sp_val[10]),
    .S(reg_sp_wr),
    .Y(_0622_)
  );
  \$_MUX_  _2330_ (
    .A(_0622_),
    .B(pc_sw[10]),
    .S(_0599_),
    .Y(_0006_[10])
  );
  \$_AND_  _2331_ (
    .A(reg_dest_val[11]),
    .B(_0604_),
    .Y(pc_sw[11])
  );
  \$_AND_  _2332_ (
    .A(_0619_),
    .B(reg_src[10]),
    .Y(_0623_)
  );
  \$_XOR_  _2333_ (
    .A(_0623_),
    .B(reg_src[11]),
    .Y(_0624_)
  );
  \$_MUX_  _2334_ (
    .A(_0624_),
    .B(r1[11]),
    .S(_0598_),
    .Y(_0625_)
  );
  \$_MUX_  _2335_ (
    .A(_0625_),
    .B(reg_sp_val[11]),
    .S(reg_sp_wr),
    .Y(_0626_)
  );
  \$_MUX_  _2336_ (
    .A(_0626_),
    .B(pc_sw[11]),
    .S(_0599_),
    .Y(_0006_[11])
  );
  \$_AND_  _2337_ (
    .A(reg_dest_val[12]),
    .B(_0604_),
    .Y(pc_sw[12])
  );
  \$_AND_  _2338_ (
    .A(_0623_),
    .B(reg_src[11]),
    .Y(_0627_)
  );
  \$_XOR_  _2339_ (
    .A(_0627_),
    .B(reg_src[12]),
    .Y(_0628_)
  );
  \$_MUX_  _2340_ (
    .A(_0628_),
    .B(r1[12]),
    .S(_0598_),
    .Y(_0629_)
  );
  \$_MUX_  _2341_ (
    .A(_0629_),
    .B(reg_sp_val[12]),
    .S(reg_sp_wr),
    .Y(_0630_)
  );
  \$_MUX_  _2342_ (
    .A(_0630_),
    .B(pc_sw[12]),
    .S(_0599_),
    .Y(_0006_[12])
  );
  \$_AND_  _2343_ (
    .A(reg_dest_val[13]),
    .B(_0604_),
    .Y(pc_sw[13])
  );
  \$_AND_  _2344_ (
    .A(_0627_),
    .B(reg_src[12]),
    .Y(_0631_)
  );
  \$_XOR_  _2345_ (
    .A(_0631_),
    .B(reg_src[13]),
    .Y(_0632_)
  );
  \$_MUX_  _2346_ (
    .A(_0632_),
    .B(r1[13]),
    .S(_0598_),
    .Y(_0633_)
  );
  \$_MUX_  _2347_ (
    .A(_0633_),
    .B(reg_sp_val[13]),
    .S(reg_sp_wr),
    .Y(_0634_)
  );
  \$_MUX_  _2348_ (
    .A(_0634_),
    .B(pc_sw[13]),
    .S(_0599_),
    .Y(_0006_[13])
  );
  \$_AND_  _2349_ (
    .A(reg_dest_val[14]),
    .B(_0604_),
    .Y(pc_sw[14])
  );
  \$_AND_  _2350_ (
    .A(_0631_),
    .B(reg_src[13]),
    .Y(_0635_)
  );
  \$_XOR_  _2351_ (
    .A(_0635_),
    .B(reg_src[14]),
    .Y(_0636_)
  );
  \$_MUX_  _2352_ (
    .A(_0636_),
    .B(r1[14]),
    .S(_0598_),
    .Y(_0637_)
  );
  \$_MUX_  _2353_ (
    .A(_0637_),
    .B(reg_sp_val[14]),
    .S(reg_sp_wr),
    .Y(_0638_)
  );
  \$_MUX_  _2354_ (
    .A(_0638_),
    .B(pc_sw[14]),
    .S(_0599_),
    .Y(_0006_[14])
  );
  \$_AND_  _2355_ (
    .A(reg_dest_val[15]),
    .B(_0604_),
    .Y(pc_sw[15])
  );
  \$_AND_  _2356_ (
    .A(_0635_),
    .B(reg_src[14]),
    .Y(_0639_)
  );
  \$_XOR_  _2357_ (
    .A(_0639_),
    .B(reg_src[15]),
    .Y(_0640_)
  );
  \$_MUX_  _2358_ (
    .A(_0640_),
    .B(r1[15]),
    .S(_0598_),
    .Y(_0641_)
  );
  \$_MUX_  _2359_ (
    .A(_0641_),
    .B(reg_sp_val[15]),
    .S(reg_sp_wr),
    .Y(_0642_)
  );
  \$_MUX_  _2360_ (
    .A(_0642_),
    .B(pc_sw[15]),
    .S(_0599_),
    .Y(_0006_[15])
  );
  \$_XOR_  _2361_ (
    .A(_0609_),
    .B(_0608_),
    .Y(_0643_)
  );
  \$_MUX_  _2362_ (
    .A(_0643_),
    .B(r1[1]),
    .S(_0598_),
    .Y(_0644_)
  );
  \$_MUX_  _2363_ (
    .A(_0644_),
    .B(reg_sp_val[1]),
    .S(reg_sp_wr),
    .Y(_0645_)
  );
  \$_MUX_  _2364_ (
    .A(_0645_),
    .B(reg_dest_val[1]),
    .S(_0599_),
    .Y(_0006_[1])
  );
  \$_XOR_  _2365_ (
    .A(_0611_),
    .B(reg_src[2]),
    .Y(_0646_)
  );
  \$_MUX_  _2366_ (
    .A(_0646_),
    .B(r1[2]),
    .S(_0598_),
    .Y(_0647_)
  );
  \$_MUX_  _2367_ (
    .A(_0647_),
    .B(reg_sp_val[2]),
    .S(reg_sp_wr),
    .Y(_0648_)
  );
  \$_MUX_  _2368_ (
    .A(_0648_),
    .B(reg_dest_val[2]),
    .S(_0599_),
    .Y(_0006_[2])
  );
  \$_XOR_  _2369_ (
    .A(_0612_),
    .B(reg_src[3]),
    .Y(_0649_)
  );
  \$_MUX_  _2370_ (
    .A(_0649_),
    .B(r1[3]),
    .S(_0598_),
    .Y(_0650_)
  );
  \$_MUX_  _2371_ (
    .A(_0650_),
    .B(reg_sp_val[3]),
    .S(reg_sp_wr),
    .Y(_0651_)
  );
  \$_MUX_  _2372_ (
    .A(_0651_),
    .B(reg_dest_val[3]),
    .S(_0599_),
    .Y(_0006_[3])
  );
  \$_XOR_  _2373_ (
    .A(_0613_),
    .B(reg_src[4]),
    .Y(_0652_)
  );
  \$_MUX_  _2374_ (
    .A(_0652_),
    .B(r1[4]),
    .S(_0598_),
    .Y(_0653_)
  );
  \$_MUX_  _2375_ (
    .A(_0653_),
    .B(reg_sp_val[4]),
    .S(reg_sp_wr),
    .Y(_0654_)
  );
  \$_MUX_  _2376_ (
    .A(_0654_),
    .B(reg_dest_val[4]),
    .S(_0599_),
    .Y(_0006_[4])
  );
  \$_XOR_  _2377_ (
    .A(_0614_),
    .B(reg_src[5]),
    .Y(_0655_)
  );
  \$_MUX_  _2378_ (
    .A(_0655_),
    .B(r1[5]),
    .S(_0598_),
    .Y(_0656_)
  );
  \$_MUX_  _2379_ (
    .A(_0656_),
    .B(reg_sp_val[5]),
    .S(reg_sp_wr),
    .Y(_0657_)
  );
  \$_MUX_  _2380_ (
    .A(_0657_),
    .B(reg_dest_val[5]),
    .S(_0599_),
    .Y(_0006_[5])
  );
  \$_XOR_  _2381_ (
    .A(_0615_),
    .B(reg_src[6]),
    .Y(_0658_)
  );
  \$_MUX_  _2382_ (
    .A(_0658_),
    .B(r1[6]),
    .S(_0598_),
    .Y(_0659_)
  );
  \$_MUX_  _2383_ (
    .A(_0659_),
    .B(reg_sp_val[6]),
    .S(reg_sp_wr),
    .Y(_0660_)
  );
  \$_MUX_  _2384_ (
    .A(_0660_),
    .B(reg_dest_val[6]),
    .S(_0599_),
    .Y(_0006_[6])
  );
  \$_XOR_  _2385_ (
    .A(_0616_),
    .B(reg_src[7]),
    .Y(_0661_)
  );
  \$_MUX_  _2386_ (
    .A(_0661_),
    .B(r1[7]),
    .S(_0598_),
    .Y(_0662_)
  );
  \$_MUX_  _2387_ (
    .A(_0662_),
    .B(reg_sp_val[7]),
    .S(reg_sp_wr),
    .Y(_0663_)
  );
  \$_MUX_  _2388_ (
    .A(_0663_),
    .B(reg_dest_val[7]),
    .S(_0599_),
    .Y(_0006_[7])
  );
  \$_AND_  _2389_ (
    .A(reg_dest_val[8]),
    .B(_0604_),
    .Y(pc_sw[8])
  );
  \$_XOR_  _2390_ (
    .A(_0617_),
    .B(reg_src[8]),
    .Y(_0664_)
  );
  \$_MUX_  _2391_ (
    .A(_0664_),
    .B(r1[8]),
    .S(_0598_),
    .Y(_0665_)
  );
  \$_MUX_  _2392_ (
    .A(_0665_),
    .B(reg_sp_val[8]),
    .S(reg_sp_wr),
    .Y(_0666_)
  );
  \$_MUX_  _2393_ (
    .A(_0666_),
    .B(pc_sw[8]),
    .S(_0599_),
    .Y(_0006_[8])
  );
  \$_AND_  _2394_ (
    .A(reg_dest_val[9]),
    .B(_0604_),
    .Y(pc_sw[9])
  );
  \$_XOR_  _2395_ (
    .A(_0618_),
    .B(reg_src[9]),
    .Y(_0667_)
  );
  \$_MUX_  _2396_ (
    .A(_0667_),
    .B(r1[9]),
    .S(_0598_),
    .Y(_0668_)
  );
  \$_MUX_  _2397_ (
    .A(_0668_),
    .B(reg_sp_val[9]),
    .S(reg_sp_wr),
    .Y(_0669_)
  );
  \$_MUX_  _2398_ (
    .A(_0669_),
    .B(pc_sw[9]),
    .S(_0599_),
    .Y(_0006_[9])
  );
  \$_MUX_  _2399_ (
    .A(r2[0]),
    .B(reg_dest_val[0]),
    .S(_0120_),
    .Y(_0670_)
  );
  \$_MUX_  _2400_ (
    .A(_0670_),
    .B(alu_stat[0]),
    .S(alu_stat_wr[0]),
    .Y(_0671_)
  );
  \$_AND_  _2401_ (
    .A(_0671_),
    .B(_0914_),
    .Y(_0007_[0])
  );
  \$_MUX_  _2402_ (
    .A(r2[1]),
    .B(reg_dest_val[1]),
    .S(_0120_),
    .Y(_0672_)
  );
  \$_MUX_  _2403_ (
    .A(_0672_),
    .B(alu_stat[1]),
    .S(alu_stat_wr[1]),
    .Y(_0673_)
  );
  \$_AND_  _2404_ (
    .A(_0673_),
    .B(_0914_),
    .Y(_0007_[1])
  );
  \$_MUX_  _2405_ (
    .A(r2[2]),
    .B(reg_dest_val[2]),
    .S(_0120_),
    .Y(_0674_)
  );
  \$_MUX_  _2406_ (
    .A(_0674_),
    .B(alu_stat[2]),
    .S(alu_stat_wr[2]),
    .Y(_0675_)
  );
  \$_AND_  _2407_ (
    .A(_0675_),
    .B(_0914_),
    .Y(_0007_[2])
  );
  \$_MUX_  _2408_ (
    .A(gie),
    .B(reg_dest_val[3]),
    .S(_0120_),
    .Y(_0676_)
  );
  \$_AND_  _2409_ (
    .A(_0676_),
    .B(_0914_),
    .Y(_0007_[3])
  );
  \$_AND_  _2410_ (
    .A(_0121_),
    .B(_0914_),
    .Y(_0007_[4])
  );
  \$_MUX_  _2411_ (
    .A(oscoff),
    .B(reg_dest_val[5]),
    .S(_0120_),
    .Y(_0677_)
  );
  \$_AND_  _2412_ (
    .A(_0677_),
    .B(_0914_),
    .Y(_0007_[5])
  );
  \$_MUX_  _2413_ (
    .A(r2[7]),
    .B(reg_dest_val[7]),
    .S(_0120_),
    .Y(_0678_)
  );
  \$_AND_  _2414_ (
    .A(_0678_),
    .B(_0914_),
    .Y(_0007_[7])
  );
  \$_MUX_  _2415_ (
    .A(r2[8]),
    .B(pc_sw[8]),
    .S(_0120_),
    .Y(_0679_)
  );
  \$_MUX_  _2416_ (
    .A(_0679_),
    .B(alu_stat[3]),
    .S(alu_stat_wr[3]),
    .Y(_0680_)
  );
  \$_AND_  _2417_ (
    .A(_0680_),
    .B(_0914_),
    .Y(_0007_[8])
  );
  \$_AND_  _2418_ (
    .A(inst_dest[3]),
    .B(reg_dest_wr),
    .Y(_0681_)
  );
  \$_MUX_  _2419_ (
    .A(r3[0]),
    .B(reg_dest_val[0]),
    .S(_0681_),
    .Y(_0008_[0])
  );
  \$_INV_  _2420_ (
    .A(_0681_),
    .Y(_0682_)
  );
  \$_MUX_  _2421_ (
    .A(pc_sw[10]),
    .B(r3[10]),
    .S(_0682_),
    .Y(_0008_[10])
  );
  \$_MUX_  _2422_ (
    .A(pc_sw[11]),
    .B(r3[11]),
    .S(_0682_),
    .Y(_0008_[11])
  );
  \$_MUX_  _2423_ (
    .A(pc_sw[12]),
    .B(r3[12]),
    .S(_0682_),
    .Y(_0008_[12])
  );
  \$_MUX_  _2424_ (
    .A(pc_sw[13]),
    .B(r3[13]),
    .S(_0682_),
    .Y(_0008_[13])
  );
  \$_MUX_  _2425_ (
    .A(pc_sw[14]),
    .B(r3[14]),
    .S(_0682_),
    .Y(_0008_[14])
  );
  \$_MUX_  _2426_ (
    .A(pc_sw[15]),
    .B(r3[15]),
    .S(_0682_),
    .Y(_0008_[15])
  );
  \$_MUX_  _2427_ (
    .A(r3[1]),
    .B(reg_dest_val[1]),
    .S(_0681_),
    .Y(_0008_[1])
  );
  \$_MUX_  _2428_ (
    .A(r3[2]),
    .B(reg_dest_val[2]),
    .S(_0681_),
    .Y(_0008_[2])
  );
  \$_MUX_  _2429_ (
    .A(r3[3]),
    .B(reg_dest_val[3]),
    .S(_0681_),
    .Y(_0008_[3])
  );
  \$_MUX_  _2430_ (
    .A(r3[4]),
    .B(reg_dest_val[4]),
    .S(_0681_),
    .Y(_0008_[4])
  );
  \$_MUX_  _2431_ (
    .A(r3[5]),
    .B(reg_dest_val[5]),
    .S(_0681_),
    .Y(_0008_[5])
  );
  \$_MUX_  _2432_ (
    .A(r3[6]),
    .B(reg_dest_val[6]),
    .S(_0681_),
    .Y(_0008_[6])
  );
  \$_MUX_  _2433_ (
    .A(r3[7]),
    .B(reg_dest_val[7]),
    .S(_0681_),
    .Y(_0008_[7])
  );
  \$_MUX_  _2434_ (
    .A(pc_sw[8]),
    .B(r3[8]),
    .S(_0682_),
    .Y(_0008_[8])
  );
  \$_MUX_  _2435_ (
    .A(pc_sw[9]),
    .B(r3[9]),
    .S(_0682_),
    .Y(_0008_[9])
  );
  \$_AND_  _2436_ (
    .A(inst_dest[4]),
    .B(reg_dest_wr),
    .Y(_0683_)
  );
  \$_INV_  _2437_ (
    .A(_0922_),
    .Y(_0684_)
  );
  \$_OR_  _2438_ (
    .A(_0684_),
    .B(_0596_),
    .Y(_0685_)
  );
  \$_XOR_  _2439_ (
    .A(_0605_),
    .B(reg_src[0]),
    .Y(_0686_)
  );
  \$_MUX_  _2440_ (
    .A(_0686_),
    .B(r4[0]),
    .S(_0685_),
    .Y(_0687_)
  );
  \$_MUX_  _2441_ (
    .A(_0687_),
    .B(reg_dest_val[0]),
    .S(_0683_),
    .Y(_0009_[0])
  );
  \$_MUX_  _2442_ (
    .A(_0620_),
    .B(r4[10]),
    .S(_0685_),
    .Y(_0688_)
  );
  \$_MUX_  _2443_ (
    .A(_0688_),
    .B(pc_sw[10]),
    .S(_0683_),
    .Y(_0009_[10])
  );
  \$_MUX_  _2444_ (
    .A(_0624_),
    .B(r4[11]),
    .S(_0685_),
    .Y(_0689_)
  );
  \$_MUX_  _2445_ (
    .A(_0689_),
    .B(pc_sw[11]),
    .S(_0683_),
    .Y(_0009_[11])
  );
  \$_MUX_  _2446_ (
    .A(_0628_),
    .B(r4[12]),
    .S(_0685_),
    .Y(_0690_)
  );
  \$_MUX_  _2447_ (
    .A(_0690_),
    .B(pc_sw[12]),
    .S(_0683_),
    .Y(_0009_[12])
  );
  \$_MUX_  _2448_ (
    .A(_0632_),
    .B(r4[13]),
    .S(_0685_),
    .Y(_0691_)
  );
  \$_MUX_  _2449_ (
    .A(_0691_),
    .B(pc_sw[13]),
    .S(_0683_),
    .Y(_0009_[13])
  );
  \$_MUX_  _2450_ (
    .A(_0636_),
    .B(r4[14]),
    .S(_0685_),
    .Y(_0692_)
  );
  \$_MUX_  _2451_ (
    .A(_0692_),
    .B(pc_sw[14]),
    .S(_0683_),
    .Y(_0009_[14])
  );
  \$_MUX_  _2452_ (
    .A(_0640_),
    .B(r4[15]),
    .S(_0685_),
    .Y(_0693_)
  );
  \$_MUX_  _2453_ (
    .A(_0693_),
    .B(pc_sw[15]),
    .S(_0683_),
    .Y(_0009_[15])
  );
  \$_MUX_  _2454_ (
    .A(_0643_),
    .B(r4[1]),
    .S(_0685_),
    .Y(_0694_)
  );
  \$_MUX_  _2455_ (
    .A(_0694_),
    .B(reg_dest_val[1]),
    .S(_0683_),
    .Y(_0009_[1])
  );
  \$_MUX_  _2456_ (
    .A(_0646_),
    .B(r4[2]),
    .S(_0685_),
    .Y(_0695_)
  );
  \$_MUX_  _2457_ (
    .A(_0695_),
    .B(reg_dest_val[2]),
    .S(_0683_),
    .Y(_0009_[2])
  );
  \$_MUX_  _2458_ (
    .A(_0649_),
    .B(r4[3]),
    .S(_0685_),
    .Y(_0696_)
  );
  \$_MUX_  _2459_ (
    .A(_0696_),
    .B(reg_dest_val[3]),
    .S(_0683_),
    .Y(_0009_[3])
  );
  \$_MUX_  _2460_ (
    .A(_0652_),
    .B(r4[4]),
    .S(_0685_),
    .Y(_0697_)
  );
  \$_MUX_  _2461_ (
    .A(_0697_),
    .B(reg_dest_val[4]),
    .S(_0683_),
    .Y(_0009_[4])
  );
  \$_MUX_  _2462_ (
    .A(_0655_),
    .B(r4[5]),
    .S(_0685_),
    .Y(_0698_)
  );
  \$_MUX_  _2463_ (
    .A(_0698_),
    .B(reg_dest_val[5]),
    .S(_0683_),
    .Y(_0009_[5])
  );
  \$_MUX_  _2464_ (
    .A(_0658_),
    .B(r4[6]),
    .S(_0685_),
    .Y(_0699_)
  );
  \$_MUX_  _2465_ (
    .A(_0699_),
    .B(reg_dest_val[6]),
    .S(_0683_),
    .Y(_0009_[6])
  );
  \$_MUX_  _2466_ (
    .A(_0661_),
    .B(r4[7]),
    .S(_0685_),
    .Y(_0700_)
  );
  \$_MUX_  _2467_ (
    .A(_0700_),
    .B(reg_dest_val[7]),
    .S(_0683_),
    .Y(_0009_[7])
  );
  \$_MUX_  _2468_ (
    .A(_0664_),
    .B(r4[8]),
    .S(_0685_),
    .Y(_0701_)
  );
  \$_MUX_  _2469_ (
    .A(_0701_),
    .B(pc_sw[8]),
    .S(_0683_),
    .Y(_0009_[8])
  );
  \$_MUX_  _2470_ (
    .A(_0667_),
    .B(r4[9]),
    .S(_0685_),
    .Y(_0702_)
  );
  \$_MUX_  _2471_ (
    .A(_0702_),
    .B(pc_sw[9]),
    .S(_0683_),
    .Y(_0009_[9])
  );
  \$_AND_  _2472_ (
    .A(inst_dest[5]),
    .B(reg_dest_wr),
    .Y(_0703_)
  );
  \$_INV_  _2473_ (
    .A(_0946_),
    .Y(_0704_)
  );
  \$_OR_  _2474_ (
    .A(_0704_),
    .B(_0596_),
    .Y(_0705_)
  );
  \$_MUX_  _2475_ (
    .A(_0686_),
    .B(r5[0]),
    .S(_0705_),
    .Y(_0706_)
  );
  \$_MUX_  _2476_ (
    .A(_0706_),
    .B(reg_dest_val[0]),
    .S(_0703_),
    .Y(_0010_[0])
  );
  \$_MUX_  _2477_ (
    .A(_0620_),
    .B(r5[10]),
    .S(_0705_),
    .Y(_0707_)
  );
  \$_MUX_  _2478_ (
    .A(_0707_),
    .B(pc_sw[10]),
    .S(_0703_),
    .Y(_0010_[10])
  );
  \$_MUX_  _2479_ (
    .A(_0624_),
    .B(r5[11]),
    .S(_0705_),
    .Y(_0708_)
  );
  \$_MUX_  _2480_ (
    .A(_0708_),
    .B(pc_sw[11]),
    .S(_0703_),
    .Y(_0010_[11])
  );
  \$_MUX_  _2481_ (
    .A(_0628_),
    .B(r5[12]),
    .S(_0705_),
    .Y(_0709_)
  );
  \$_MUX_  _2482_ (
    .A(_0709_),
    .B(pc_sw[12]),
    .S(_0703_),
    .Y(_0010_[12])
  );
  \$_MUX_  _2483_ (
    .A(_0632_),
    .B(r5[13]),
    .S(_0705_),
    .Y(_0710_)
  );
  \$_MUX_  _2484_ (
    .A(_0710_),
    .B(pc_sw[13]),
    .S(_0703_),
    .Y(_0010_[13])
  );
  \$_MUX_  _2485_ (
    .A(_0636_),
    .B(r5[14]),
    .S(_0705_),
    .Y(_0711_)
  );
  \$_MUX_  _2486_ (
    .A(_0711_),
    .B(pc_sw[14]),
    .S(_0703_),
    .Y(_0010_[14])
  );
  \$_MUX_  _2487_ (
    .A(_0640_),
    .B(r5[15]),
    .S(_0705_),
    .Y(_0712_)
  );
  \$_MUX_  _2488_ (
    .A(_0712_),
    .B(pc_sw[15]),
    .S(_0703_),
    .Y(_0010_[15])
  );
  \$_MUX_  _2489_ (
    .A(_0643_),
    .B(r5[1]),
    .S(_0705_),
    .Y(_0713_)
  );
  \$_MUX_  _2490_ (
    .A(_0713_),
    .B(reg_dest_val[1]),
    .S(_0703_),
    .Y(_0010_[1])
  );
  \$_MUX_  _2491_ (
    .A(_0646_),
    .B(r5[2]),
    .S(_0705_),
    .Y(_0714_)
  );
  \$_MUX_  _2492_ (
    .A(_0714_),
    .B(reg_dest_val[2]),
    .S(_0703_),
    .Y(_0010_[2])
  );
  \$_MUX_  _2493_ (
    .A(_0649_),
    .B(r5[3]),
    .S(_0705_),
    .Y(_0715_)
  );
  \$_MUX_  _2494_ (
    .A(_0715_),
    .B(reg_dest_val[3]),
    .S(_0703_),
    .Y(_0010_[3])
  );
  \$_MUX_  _2495_ (
    .A(_0652_),
    .B(r5[4]),
    .S(_0705_),
    .Y(_0716_)
  );
  \$_MUX_  _2496_ (
    .A(_0716_),
    .B(reg_dest_val[4]),
    .S(_0703_),
    .Y(_0010_[4])
  );
  \$_MUX_  _2497_ (
    .A(_0655_),
    .B(r5[5]),
    .S(_0705_),
    .Y(_0717_)
  );
  \$_MUX_  _2498_ (
    .A(_0717_),
    .B(reg_dest_val[5]),
    .S(_0703_),
    .Y(_0010_[5])
  );
  \$_MUX_  _2499_ (
    .A(_0658_),
    .B(r5[6]),
    .S(_0705_),
    .Y(_0718_)
  );
  \$_MUX_  _2500_ (
    .A(_0718_),
    .B(reg_dest_val[6]),
    .S(_0703_),
    .Y(_0010_[6])
  );
  \$_MUX_  _2501_ (
    .A(_0661_),
    .B(r5[7]),
    .S(_0705_),
    .Y(_0719_)
  );
  \$_MUX_  _2502_ (
    .A(_0719_),
    .B(reg_dest_val[7]),
    .S(_0703_),
    .Y(_0010_[7])
  );
  \$_MUX_  _2503_ (
    .A(_0664_),
    .B(r5[8]),
    .S(_0705_),
    .Y(_0720_)
  );
  \$_MUX_  _2504_ (
    .A(_0720_),
    .B(pc_sw[8]),
    .S(_0703_),
    .Y(_0010_[8])
  );
  \$_MUX_  _2505_ (
    .A(_0667_),
    .B(r5[9]),
    .S(_0705_),
    .Y(_0721_)
  );
  \$_MUX_  _2506_ (
    .A(_0721_),
    .B(pc_sw[9]),
    .S(_0703_),
    .Y(_0010_[9])
  );
  \$_AND_  _2507_ (
    .A(inst_dest[6]),
    .B(reg_dest_wr),
    .Y(_0722_)
  );
  \$_INV_  _2508_ (
    .A(_0948_),
    .Y(_0723_)
  );
  \$_OR_  _2509_ (
    .A(_0723_),
    .B(_0596_),
    .Y(_0724_)
  );
  \$_MUX_  _2510_ (
    .A(_0686_),
    .B(r6[0]),
    .S(_0724_),
    .Y(_0725_)
  );
  \$_MUX_  _2511_ (
    .A(_0725_),
    .B(reg_dest_val[0]),
    .S(_0722_),
    .Y(_0011_[0])
  );
  \$_MUX_  _2512_ (
    .A(_0620_),
    .B(r6[10]),
    .S(_0724_),
    .Y(_0726_)
  );
  \$_MUX_  _2513_ (
    .A(_0726_),
    .B(pc_sw[10]),
    .S(_0722_),
    .Y(_0011_[10])
  );
  \$_MUX_  _2514_ (
    .A(_0624_),
    .B(r6[11]),
    .S(_0724_),
    .Y(_0727_)
  );
  \$_MUX_  _2515_ (
    .A(_0727_),
    .B(pc_sw[11]),
    .S(_0722_),
    .Y(_0011_[11])
  );
  \$_MUX_  _2516_ (
    .A(_0628_),
    .B(r6[12]),
    .S(_0724_),
    .Y(_0728_)
  );
  \$_MUX_  _2517_ (
    .A(_0728_),
    .B(pc_sw[12]),
    .S(_0722_),
    .Y(_0011_[12])
  );
  \$_MUX_  _2518_ (
    .A(_0632_),
    .B(r6[13]),
    .S(_0724_),
    .Y(_0729_)
  );
  \$_MUX_  _2519_ (
    .A(_0729_),
    .B(pc_sw[13]),
    .S(_0722_),
    .Y(_0011_[13])
  );
  \$_MUX_  _2520_ (
    .A(_0636_),
    .B(r6[14]),
    .S(_0724_),
    .Y(_0730_)
  );
  \$_MUX_  _2521_ (
    .A(_0730_),
    .B(pc_sw[14]),
    .S(_0722_),
    .Y(_0011_[14])
  );
  \$_MUX_  _2522_ (
    .A(_0640_),
    .B(r6[15]),
    .S(_0724_),
    .Y(_0731_)
  );
  \$_MUX_  _2523_ (
    .A(_0731_),
    .B(pc_sw[15]),
    .S(_0722_),
    .Y(_0011_[15])
  );
  \$_MUX_  _2524_ (
    .A(_0643_),
    .B(r6[1]),
    .S(_0724_),
    .Y(_0732_)
  );
  \$_MUX_  _2525_ (
    .A(_0732_),
    .B(reg_dest_val[1]),
    .S(_0722_),
    .Y(_0011_[1])
  );
  \$_MUX_  _2526_ (
    .A(_0646_),
    .B(r6[2]),
    .S(_0724_),
    .Y(_0733_)
  );
  \$_MUX_  _2527_ (
    .A(_0733_),
    .B(reg_dest_val[2]),
    .S(_0722_),
    .Y(_0011_[2])
  );
  \$_MUX_  _2528_ (
    .A(_0649_),
    .B(r6[3]),
    .S(_0724_),
    .Y(_0734_)
  );
  \$_MUX_  _2529_ (
    .A(_0734_),
    .B(reg_dest_val[3]),
    .S(_0722_),
    .Y(_0011_[3])
  );
  \$_MUX_  _2530_ (
    .A(_0652_),
    .B(r6[4]),
    .S(_0724_),
    .Y(_0735_)
  );
  \$_MUX_  _2531_ (
    .A(_0735_),
    .B(reg_dest_val[4]),
    .S(_0722_),
    .Y(_0011_[4])
  );
  \$_MUX_  _2532_ (
    .A(_0655_),
    .B(r6[5]),
    .S(_0724_),
    .Y(_0736_)
  );
  \$_MUX_  _2533_ (
    .A(_0736_),
    .B(reg_dest_val[5]),
    .S(_0722_),
    .Y(_0011_[5])
  );
  \$_MUX_  _2534_ (
    .A(_0658_),
    .B(r6[6]),
    .S(_0724_),
    .Y(_0737_)
  );
  \$_MUX_  _2535_ (
    .A(_0737_),
    .B(reg_dest_val[6]),
    .S(_0722_),
    .Y(_0011_[6])
  );
  \$_MUX_  _2536_ (
    .A(_0661_),
    .B(r6[7]),
    .S(_0724_),
    .Y(_0738_)
  );
  \$_MUX_  _2537_ (
    .A(_0738_),
    .B(reg_dest_val[7]),
    .S(_0722_),
    .Y(_0011_[7])
  );
  \$_MUX_  _2538_ (
    .A(_0664_),
    .B(r6[8]),
    .S(_0724_),
    .Y(_0739_)
  );
  \$_MUX_  _2539_ (
    .A(_0739_),
    .B(pc_sw[8]),
    .S(_0722_),
    .Y(_0011_[8])
  );
  \$_MUX_  _2540_ (
    .A(_0667_),
    .B(r6[9]),
    .S(_0724_),
    .Y(_0740_)
  );
  \$_MUX_  _2541_ (
    .A(_0740_),
    .B(pc_sw[9]),
    .S(_0722_),
    .Y(_0011_[9])
  );
  \$_AND_  _2542_ (
    .A(inst_dest[7]),
    .B(reg_dest_wr),
    .Y(_0741_)
  );
  \$_INV_  _2543_ (
    .A(_0951_),
    .Y(_0742_)
  );
  \$_OR_  _2544_ (
    .A(_0742_),
    .B(_0596_),
    .Y(_0743_)
  );
  \$_MUX_  _2545_ (
    .A(_0686_),
    .B(r7[0]),
    .S(_0743_),
    .Y(_0744_)
  );
  \$_MUX_  _2546_ (
    .A(_0744_),
    .B(reg_dest_val[0]),
    .S(_0741_),
    .Y(_0012_[0])
  );
  \$_MUX_  _2547_ (
    .A(_0620_),
    .B(r7[10]),
    .S(_0743_),
    .Y(_0745_)
  );
  \$_MUX_  _2548_ (
    .A(_0745_),
    .B(pc_sw[10]),
    .S(_0741_),
    .Y(_0012_[10])
  );
  \$_MUX_  _2549_ (
    .A(_0624_),
    .B(r7[11]),
    .S(_0743_),
    .Y(_0746_)
  );
  \$_MUX_  _2550_ (
    .A(_0746_),
    .B(pc_sw[11]),
    .S(_0741_),
    .Y(_0012_[11])
  );
  \$_MUX_  _2551_ (
    .A(_0628_),
    .B(r7[12]),
    .S(_0743_),
    .Y(_0747_)
  );
  \$_MUX_  _2552_ (
    .A(_0747_),
    .B(pc_sw[12]),
    .S(_0741_),
    .Y(_0012_[12])
  );
  \$_MUX_  _2553_ (
    .A(_0632_),
    .B(r7[13]),
    .S(_0743_),
    .Y(_0748_)
  );
  \$_MUX_  _2554_ (
    .A(_0748_),
    .B(pc_sw[13]),
    .S(_0741_),
    .Y(_0012_[13])
  );
  \$_MUX_  _2555_ (
    .A(_0636_),
    .B(r7[14]),
    .S(_0743_),
    .Y(_0749_)
  );
  \$_MUX_  _2556_ (
    .A(_0749_),
    .B(pc_sw[14]),
    .S(_0741_),
    .Y(_0012_[14])
  );
  \$_MUX_  _2557_ (
    .A(_0640_),
    .B(r7[15]),
    .S(_0743_),
    .Y(_0750_)
  );
  \$_MUX_  _2558_ (
    .A(_0750_),
    .B(pc_sw[15]),
    .S(_0741_),
    .Y(_0012_[15])
  );
  \$_MUX_  _2559_ (
    .A(_0643_),
    .B(r7[1]),
    .S(_0743_),
    .Y(_0751_)
  );
  \$_MUX_  _2560_ (
    .A(_0751_),
    .B(reg_dest_val[1]),
    .S(_0741_),
    .Y(_0012_[1])
  );
  \$_MUX_  _2561_ (
    .A(_0646_),
    .B(r7[2]),
    .S(_0743_),
    .Y(_0752_)
  );
  \$_MUX_  _2562_ (
    .A(_0752_),
    .B(reg_dest_val[2]),
    .S(_0741_),
    .Y(_0012_[2])
  );
  \$_MUX_  _2563_ (
    .A(_0649_),
    .B(r7[3]),
    .S(_0743_),
    .Y(_0753_)
  );
  \$_MUX_  _2564_ (
    .A(_0753_),
    .B(reg_dest_val[3]),
    .S(_0741_),
    .Y(_0012_[3])
  );
  \$_MUX_  _2565_ (
    .A(_0652_),
    .B(r7[4]),
    .S(_0743_),
    .Y(_0754_)
  );
  \$_MUX_  _2566_ (
    .A(_0754_),
    .B(reg_dest_val[4]),
    .S(_0741_),
    .Y(_0012_[4])
  );
  \$_MUX_  _2567_ (
    .A(_0655_),
    .B(r7[5]),
    .S(_0743_),
    .Y(_0755_)
  );
  \$_MUX_  _2568_ (
    .A(_0755_),
    .B(reg_dest_val[5]),
    .S(_0741_),
    .Y(_0012_[5])
  );
  \$_MUX_  _2569_ (
    .A(_0658_),
    .B(r7[6]),
    .S(_0743_),
    .Y(_0756_)
  );
  \$_MUX_  _2570_ (
    .A(_0756_),
    .B(reg_dest_val[6]),
    .S(_0741_),
    .Y(_0012_[6])
  );
  \$_MUX_  _2571_ (
    .A(_0661_),
    .B(r7[7]),
    .S(_0743_),
    .Y(_0757_)
  );
  \$_MUX_  _2572_ (
    .A(_0757_),
    .B(reg_dest_val[7]),
    .S(_0741_),
    .Y(_0012_[7])
  );
  \$_MUX_  _2573_ (
    .A(_0664_),
    .B(r7[8]),
    .S(_0743_),
    .Y(_0758_)
  );
  \$_MUX_  _2574_ (
    .A(_0758_),
    .B(pc_sw[8]),
    .S(_0741_),
    .Y(_0012_[8])
  );
  \$_MUX_  _2575_ (
    .A(_0667_),
    .B(r7[9]),
    .S(_0743_),
    .Y(_0759_)
  );
  \$_MUX_  _2576_ (
    .A(_0759_),
    .B(pc_sw[9]),
    .S(_0741_),
    .Y(_0012_[9])
  );
  \$_AND_  _2577_ (
    .A(inst_dest[8]),
    .B(reg_dest_wr),
    .Y(_0760_)
  );
  \$_INV_  _2578_ (
    .A(_0953_),
    .Y(_0761_)
  );
  \$_OR_  _2579_ (
    .A(_0761_),
    .B(_0596_),
    .Y(_0762_)
  );
  \$_MUX_  _2580_ (
    .A(_0686_),
    .B(r8[0]),
    .S(_0762_),
    .Y(_0763_)
  );
  \$_MUX_  _2581_ (
    .A(_0763_),
    .B(reg_dest_val[0]),
    .S(_0760_),
    .Y(_0013_[0])
  );
  \$_MUX_  _2582_ (
    .A(_0620_),
    .B(r8[10]),
    .S(_0762_),
    .Y(_0764_)
  );
  \$_MUX_  _2583_ (
    .A(_0764_),
    .B(pc_sw[10]),
    .S(_0760_),
    .Y(_0013_[10])
  );
  \$_MUX_  _2584_ (
    .A(_0624_),
    .B(r8[11]),
    .S(_0762_),
    .Y(_0765_)
  );
  \$_MUX_  _2585_ (
    .A(_0765_),
    .B(pc_sw[11]),
    .S(_0760_),
    .Y(_0013_[11])
  );
  \$_MUX_  _2586_ (
    .A(_0628_),
    .B(r8[12]),
    .S(_0762_),
    .Y(_0766_)
  );
  \$_MUX_  _2587_ (
    .A(_0766_),
    .B(pc_sw[12]),
    .S(_0760_),
    .Y(_0013_[12])
  );
  \$_MUX_  _2588_ (
    .A(_0632_),
    .B(r8[13]),
    .S(_0762_),
    .Y(_0767_)
  );
  \$_MUX_  _2589_ (
    .A(_0767_),
    .B(pc_sw[13]),
    .S(_0760_),
    .Y(_0013_[13])
  );
  \$_MUX_  _2590_ (
    .A(_0636_),
    .B(r8[14]),
    .S(_0762_),
    .Y(_0768_)
  );
  \$_MUX_  _2591_ (
    .A(_0768_),
    .B(pc_sw[14]),
    .S(_0760_),
    .Y(_0013_[14])
  );
  \$_MUX_  _2592_ (
    .A(_0640_),
    .B(r8[15]),
    .S(_0762_),
    .Y(_0769_)
  );
  \$_MUX_  _2593_ (
    .A(_0769_),
    .B(pc_sw[15]),
    .S(_0760_),
    .Y(_0013_[15])
  );
  \$_MUX_  _2594_ (
    .A(_0643_),
    .B(r8[1]),
    .S(_0762_),
    .Y(_0770_)
  );
  \$_MUX_  _2595_ (
    .A(_0770_),
    .B(reg_dest_val[1]),
    .S(_0760_),
    .Y(_0013_[1])
  );
  \$_MUX_  _2596_ (
    .A(_0646_),
    .B(r8[2]),
    .S(_0762_),
    .Y(_0771_)
  );
  \$_MUX_  _2597_ (
    .A(_0771_),
    .B(reg_dest_val[2]),
    .S(_0760_),
    .Y(_0013_[2])
  );
  \$_MUX_  _2598_ (
    .A(_0649_),
    .B(r8[3]),
    .S(_0762_),
    .Y(_0772_)
  );
  \$_MUX_  _2599_ (
    .A(_0772_),
    .B(reg_dest_val[3]),
    .S(_0760_),
    .Y(_0013_[3])
  );
  \$_MUX_  _2600_ (
    .A(_0652_),
    .B(r8[4]),
    .S(_0762_),
    .Y(_0773_)
  );
  \$_MUX_  _2601_ (
    .A(_0773_),
    .B(reg_dest_val[4]),
    .S(_0760_),
    .Y(_0013_[4])
  );
  \$_MUX_  _2602_ (
    .A(_0655_),
    .B(r8[5]),
    .S(_0762_),
    .Y(_0774_)
  );
  \$_MUX_  _2603_ (
    .A(_0774_),
    .B(reg_dest_val[5]),
    .S(_0760_),
    .Y(_0013_[5])
  );
  \$_MUX_  _2604_ (
    .A(_0658_),
    .B(r8[6]),
    .S(_0762_),
    .Y(_0775_)
  );
  \$_MUX_  _2605_ (
    .A(_0775_),
    .B(reg_dest_val[6]),
    .S(_0760_),
    .Y(_0013_[6])
  );
  \$_MUX_  _2606_ (
    .A(_0661_),
    .B(r8[7]),
    .S(_0762_),
    .Y(_0776_)
  );
  \$_MUX_  _2607_ (
    .A(_0776_),
    .B(reg_dest_val[7]),
    .S(_0760_),
    .Y(_0013_[7])
  );
  \$_MUX_  _2608_ (
    .A(_0664_),
    .B(r8[8]),
    .S(_0762_),
    .Y(_0777_)
  );
  \$_MUX_  _2609_ (
    .A(_0777_),
    .B(pc_sw[8]),
    .S(_0760_),
    .Y(_0013_[8])
  );
  \$_MUX_  _2610_ (
    .A(_0667_),
    .B(r8[9]),
    .S(_0762_),
    .Y(_0778_)
  );
  \$_MUX_  _2611_ (
    .A(_0778_),
    .B(pc_sw[9]),
    .S(_0760_),
    .Y(_0013_[9])
  );
  \$_AND_  _2612_ (
    .A(inst_dest[9]),
    .B(reg_dest_wr),
    .Y(_0779_)
  );
  \$_INV_  _2613_ (
    .A(_0935_),
    .Y(_0780_)
  );
  \$_OR_  _2614_ (
    .A(_0780_),
    .B(_0596_),
    .Y(_0781_)
  );
  \$_MUX_  _2615_ (
    .A(_0686_),
    .B(r9[0]),
    .S(_0781_),
    .Y(_0782_)
  );
  \$_MUX_  _2616_ (
    .A(_0782_),
    .B(reg_dest_val[0]),
    .S(_0779_),
    .Y(_0014_[0])
  );
  \$_MUX_  _2617_ (
    .A(_0620_),
    .B(r9[10]),
    .S(_0781_),
    .Y(_0783_)
  );
  \$_MUX_  _2618_ (
    .A(_0783_),
    .B(pc_sw[10]),
    .S(_0779_),
    .Y(_0014_[10])
  );
  \$_MUX_  _2619_ (
    .A(_0624_),
    .B(r9[11]),
    .S(_0781_),
    .Y(_0784_)
  );
  \$_MUX_  _2620_ (
    .A(_0784_),
    .B(pc_sw[11]),
    .S(_0779_),
    .Y(_0014_[11])
  );
  \$_MUX_  _2621_ (
    .A(_0628_),
    .B(r9[12]),
    .S(_0781_),
    .Y(_0785_)
  );
  \$_MUX_  _2622_ (
    .A(_0785_),
    .B(pc_sw[12]),
    .S(_0779_),
    .Y(_0014_[12])
  );
  \$_MUX_  _2623_ (
    .A(_0632_),
    .B(r9[13]),
    .S(_0781_),
    .Y(_0786_)
  );
  \$_MUX_  _2624_ (
    .A(_0786_),
    .B(pc_sw[13]),
    .S(_0779_),
    .Y(_0014_[13])
  );
  \$_MUX_  _2625_ (
    .A(_0636_),
    .B(r9[14]),
    .S(_0781_),
    .Y(_0787_)
  );
  \$_MUX_  _2626_ (
    .A(_0787_),
    .B(pc_sw[14]),
    .S(_0779_),
    .Y(_0014_[14])
  );
  \$_MUX_  _2627_ (
    .A(_0640_),
    .B(r9[15]),
    .S(_0781_),
    .Y(_0788_)
  );
  \$_MUX_  _2628_ (
    .A(_0788_),
    .B(pc_sw[15]),
    .S(_0779_),
    .Y(_0014_[15])
  );
  \$_MUX_  _2629_ (
    .A(_0643_),
    .B(r9[1]),
    .S(_0781_),
    .Y(_0789_)
  );
  \$_MUX_  _2630_ (
    .A(_0789_),
    .B(reg_dest_val[1]),
    .S(_0779_),
    .Y(_0014_[1])
  );
  \$_MUX_  _2631_ (
    .A(_0646_),
    .B(r9[2]),
    .S(_0781_),
    .Y(_0790_)
  );
  \$_MUX_  _2632_ (
    .A(_0790_),
    .B(reg_dest_val[2]),
    .S(_0779_),
    .Y(_0014_[2])
  );
  \$_MUX_  _2633_ (
    .A(_0649_),
    .B(r9[3]),
    .S(_0781_),
    .Y(_0791_)
  );
  \$_MUX_  _2634_ (
    .A(_0791_),
    .B(reg_dest_val[3]),
    .S(_0779_),
    .Y(_0014_[3])
  );
  \$_MUX_  _2635_ (
    .A(_0652_),
    .B(r9[4]),
    .S(_0781_),
    .Y(_0792_)
  );
  \$_MUX_  _2636_ (
    .A(_0792_),
    .B(reg_dest_val[4]),
    .S(_0779_),
    .Y(_0014_[4])
  );
  \$_MUX_  _2637_ (
    .A(_0655_),
    .B(r9[5]),
    .S(_0781_),
    .Y(_0793_)
  );
  \$_MUX_  _2638_ (
    .A(_0793_),
    .B(reg_dest_val[5]),
    .S(_0779_),
    .Y(_0014_[5])
  );
  \$_MUX_  _2639_ (
    .A(_0658_),
    .B(r9[6]),
    .S(_0781_),
    .Y(_0794_)
  );
  \$_MUX_  _2640_ (
    .A(_0794_),
    .B(reg_dest_val[6]),
    .S(_0779_),
    .Y(_0014_[6])
  );
  \$_MUX_  _2641_ (
    .A(_0661_),
    .B(r9[7]),
    .S(_0781_),
    .Y(_0795_)
  );
  \$_MUX_  _2642_ (
    .A(_0795_),
    .B(reg_dest_val[7]),
    .S(_0779_),
    .Y(_0014_[7])
  );
  \$_MUX_  _2643_ (
    .A(_0664_),
    .B(r9[8]),
    .S(_0781_),
    .Y(_0796_)
  );
  \$_MUX_  _2644_ (
    .A(_0796_),
    .B(pc_sw[8]),
    .S(_0779_),
    .Y(_0014_[8])
  );
  \$_MUX_  _2645_ (
    .A(_0667_),
    .B(r9[9]),
    .S(_0781_),
    .Y(_0797_)
  );
  \$_MUX_  _2646_ (
    .A(_0797_),
    .B(pc_sw[9]),
    .S(_0779_),
    .Y(_0014_[9])
  );
  \$_AND_  _2647_ (
    .A(inst_dest[10]),
    .B(reg_dest_wr),
    .Y(_0798_)
  );
  \$_INV_  _2648_ (
    .A(_0937_),
    .Y(_0799_)
  );
  \$_OR_  _2649_ (
    .A(_0799_),
    .B(_0596_),
    .Y(_0800_)
  );
  \$_MUX_  _2650_ (
    .A(_0686_),
    .B(r10[0]),
    .S(_0800_),
    .Y(_0801_)
  );
  \$_MUX_  _2651_ (
    .A(_0801_),
    .B(reg_dest_val[0]),
    .S(_0798_),
    .Y(_0000_[0])
  );
  \$_MUX_  _2652_ (
    .A(_0620_),
    .B(r10[10]),
    .S(_0800_),
    .Y(_0802_)
  );
  \$_MUX_  _2653_ (
    .A(_0802_),
    .B(pc_sw[10]),
    .S(_0798_),
    .Y(_0000_[10])
  );
  \$_MUX_  _2654_ (
    .A(_0624_),
    .B(r10[11]),
    .S(_0800_),
    .Y(_0803_)
  );
  \$_MUX_  _2655_ (
    .A(_0803_),
    .B(pc_sw[11]),
    .S(_0798_),
    .Y(_0000_[11])
  );
  \$_MUX_  _2656_ (
    .A(_0628_),
    .B(r10[12]),
    .S(_0800_),
    .Y(_0804_)
  );
  \$_MUX_  _2657_ (
    .A(_0804_),
    .B(pc_sw[12]),
    .S(_0798_),
    .Y(_0000_[12])
  );
  \$_MUX_  _2658_ (
    .A(_0632_),
    .B(r10[13]),
    .S(_0800_),
    .Y(_0805_)
  );
  \$_MUX_  _2659_ (
    .A(_0805_),
    .B(pc_sw[13]),
    .S(_0798_),
    .Y(_0000_[13])
  );
  \$_MUX_  _2660_ (
    .A(_0636_),
    .B(r10[14]),
    .S(_0800_),
    .Y(_0806_)
  );
  \$_MUX_  _2661_ (
    .A(_0806_),
    .B(pc_sw[14]),
    .S(_0798_),
    .Y(_0000_[14])
  );
  \$_MUX_  _2662_ (
    .A(_0640_),
    .B(r10[15]),
    .S(_0800_),
    .Y(_0807_)
  );
  \$_MUX_  _2663_ (
    .A(_0807_),
    .B(pc_sw[15]),
    .S(_0798_),
    .Y(_0000_[15])
  );
  \$_MUX_  _2664_ (
    .A(_0643_),
    .B(r10[1]),
    .S(_0800_),
    .Y(_0808_)
  );
  \$_MUX_  _2665_ (
    .A(_0808_),
    .B(reg_dest_val[1]),
    .S(_0798_),
    .Y(_0000_[1])
  );
  \$_MUX_  _2666_ (
    .A(_0646_),
    .B(r10[2]),
    .S(_0800_),
    .Y(_0809_)
  );
  \$_MUX_  _2667_ (
    .A(_0809_),
    .B(reg_dest_val[2]),
    .S(_0798_),
    .Y(_0000_[2])
  );
  \$_MUX_  _2668_ (
    .A(_0649_),
    .B(r10[3]),
    .S(_0800_),
    .Y(_0810_)
  );
  \$_MUX_  _2669_ (
    .A(_0810_),
    .B(reg_dest_val[3]),
    .S(_0798_),
    .Y(_0000_[3])
  );
  \$_MUX_  _2670_ (
    .A(_0652_),
    .B(r10[4]),
    .S(_0800_),
    .Y(_0811_)
  );
  \$_MUX_  _2671_ (
    .A(_0811_),
    .B(reg_dest_val[4]),
    .S(_0798_),
    .Y(_0000_[4])
  );
  \$_MUX_  _2672_ (
    .A(_0655_),
    .B(r10[5]),
    .S(_0800_),
    .Y(_0812_)
  );
  \$_MUX_  _2673_ (
    .A(_0812_),
    .B(reg_dest_val[5]),
    .S(_0798_),
    .Y(_0000_[5])
  );
  \$_MUX_  _2674_ (
    .A(_0658_),
    .B(r10[6]),
    .S(_0800_),
    .Y(_0813_)
  );
  \$_MUX_  _2675_ (
    .A(_0813_),
    .B(reg_dest_val[6]),
    .S(_0798_),
    .Y(_0000_[6])
  );
  \$_MUX_  _2676_ (
    .A(_0661_),
    .B(r10[7]),
    .S(_0800_),
    .Y(_0814_)
  );
  \$_MUX_  _2677_ (
    .A(_0814_),
    .B(reg_dest_val[7]),
    .S(_0798_),
    .Y(_0000_[7])
  );
  \$_MUX_  _2678_ (
    .A(_0664_),
    .B(r10[8]),
    .S(_0800_),
    .Y(_0815_)
  );
  \$_MUX_  _2679_ (
    .A(_0815_),
    .B(pc_sw[8]),
    .S(_0798_),
    .Y(_0000_[8])
  );
  \$_MUX_  _2680_ (
    .A(_0667_),
    .B(r10[9]),
    .S(_0800_),
    .Y(_0816_)
  );
  \$_MUX_  _2681_ (
    .A(_0816_),
    .B(pc_sw[9]),
    .S(_0798_),
    .Y(_0000_[9])
  );
  \$_AND_  _2682_ (
    .A(inst_dest[11]),
    .B(reg_dest_wr),
    .Y(_0817_)
  );
  \$_INV_  _2683_ (
    .A(_0940_),
    .Y(_0818_)
  );
  \$_OR_  _2684_ (
    .A(_0818_),
    .B(_0596_),
    .Y(_0819_)
  );
  \$_MUX_  _2685_ (
    .A(_0686_),
    .B(r11[0]),
    .S(_0819_),
    .Y(_0820_)
  );
  \$_MUX_  _2686_ (
    .A(_0820_),
    .B(reg_dest_val[0]),
    .S(_0817_),
    .Y(_0001_[0])
  );
  \$_MUX_  _2687_ (
    .A(_0620_),
    .B(r11[10]),
    .S(_0819_),
    .Y(_0821_)
  );
  \$_MUX_  _2688_ (
    .A(_0821_),
    .B(pc_sw[10]),
    .S(_0817_),
    .Y(_0001_[10])
  );
  \$_MUX_  _2689_ (
    .A(_0624_),
    .B(r11[11]),
    .S(_0819_),
    .Y(_0822_)
  );
  \$_MUX_  _2690_ (
    .A(_0822_),
    .B(pc_sw[11]),
    .S(_0817_),
    .Y(_0001_[11])
  );
  \$_MUX_  _2691_ (
    .A(_0628_),
    .B(r11[12]),
    .S(_0819_),
    .Y(_0823_)
  );
  \$_MUX_  _2692_ (
    .A(_0823_),
    .B(pc_sw[12]),
    .S(_0817_),
    .Y(_0001_[12])
  );
  \$_MUX_  _2693_ (
    .A(_0632_),
    .B(r11[13]),
    .S(_0819_),
    .Y(_0824_)
  );
  \$_MUX_  _2694_ (
    .A(_0824_),
    .B(pc_sw[13]),
    .S(_0817_),
    .Y(_0001_[13])
  );
  \$_MUX_  _2695_ (
    .A(_0636_),
    .B(r11[14]),
    .S(_0819_),
    .Y(_0825_)
  );
  \$_MUX_  _2696_ (
    .A(_0825_),
    .B(pc_sw[14]),
    .S(_0817_),
    .Y(_0001_[14])
  );
  \$_MUX_  _2697_ (
    .A(_0640_),
    .B(r11[15]),
    .S(_0819_),
    .Y(_0826_)
  );
  \$_MUX_  _2698_ (
    .A(_0826_),
    .B(pc_sw[15]),
    .S(_0817_),
    .Y(_0001_[15])
  );
  \$_MUX_  _2699_ (
    .A(_0643_),
    .B(r11[1]),
    .S(_0819_),
    .Y(_0827_)
  );
  \$_MUX_  _2700_ (
    .A(_0827_),
    .B(reg_dest_val[1]),
    .S(_0817_),
    .Y(_0001_[1])
  );
  \$_MUX_  _2701_ (
    .A(_0646_),
    .B(r11[2]),
    .S(_0819_),
    .Y(_0828_)
  );
  \$_MUX_  _2702_ (
    .A(_0828_),
    .B(reg_dest_val[2]),
    .S(_0817_),
    .Y(_0001_[2])
  );
  \$_MUX_  _2703_ (
    .A(_0649_),
    .B(r11[3]),
    .S(_0819_),
    .Y(_0829_)
  );
  \$_MUX_  _2704_ (
    .A(_0829_),
    .B(reg_dest_val[3]),
    .S(_0817_),
    .Y(_0001_[3])
  );
  \$_MUX_  _2705_ (
    .A(_0652_),
    .B(r11[4]),
    .S(_0819_),
    .Y(_0830_)
  );
  \$_MUX_  _2706_ (
    .A(_0830_),
    .B(reg_dest_val[4]),
    .S(_0817_),
    .Y(_0001_[4])
  );
  \$_MUX_  _2707_ (
    .A(_0655_),
    .B(r11[5]),
    .S(_0819_),
    .Y(_0831_)
  );
  \$_MUX_  _2708_ (
    .A(_0831_),
    .B(reg_dest_val[5]),
    .S(_0817_),
    .Y(_0001_[5])
  );
  \$_MUX_  _2709_ (
    .A(_0658_),
    .B(r11[6]),
    .S(_0819_),
    .Y(_0832_)
  );
  \$_MUX_  _2710_ (
    .A(_0832_),
    .B(reg_dest_val[6]),
    .S(_0817_),
    .Y(_0001_[6])
  );
  \$_MUX_  _2711_ (
    .A(_0661_),
    .B(r11[7]),
    .S(_0819_),
    .Y(_0833_)
  );
  \$_MUX_  _2712_ (
    .A(_0833_),
    .B(reg_dest_val[7]),
    .S(_0817_),
    .Y(_0001_[7])
  );
  \$_MUX_  _2713_ (
    .A(_0664_),
    .B(r11[8]),
    .S(_0819_),
    .Y(_0834_)
  );
  \$_MUX_  _2714_ (
    .A(_0834_),
    .B(pc_sw[8]),
    .S(_0817_),
    .Y(_0001_[8])
  );
  \$_MUX_  _2715_ (
    .A(_0667_),
    .B(r11[9]),
    .S(_0819_),
    .Y(_0835_)
  );
  \$_MUX_  _2716_ (
    .A(_0835_),
    .B(pc_sw[9]),
    .S(_0817_),
    .Y(_0001_[9])
  );
  \$_AND_  _2717_ (
    .A(inst_dest[12]),
    .B(reg_dest_wr),
    .Y(_0836_)
  );
  \$_INV_  _2718_ (
    .A(_0942_),
    .Y(_0837_)
  );
  \$_OR_  _2719_ (
    .A(_0837_),
    .B(_0596_),
    .Y(_0838_)
  );
  \$_MUX_  _2720_ (
    .A(_0686_),
    .B(r12[0]),
    .S(_0838_),
    .Y(_0839_)
  );
  \$_MUX_  _2721_ (
    .A(_0839_),
    .B(reg_dest_val[0]),
    .S(_0836_),
    .Y(_0002_[0])
  );
  \$_MUX_  _2722_ (
    .A(_0620_),
    .B(r12[10]),
    .S(_0838_),
    .Y(_0840_)
  );
  \$_MUX_  _2723_ (
    .A(_0840_),
    .B(pc_sw[10]),
    .S(_0836_),
    .Y(_0002_[10])
  );
  \$_MUX_  _2724_ (
    .A(_0624_),
    .B(r12[11]),
    .S(_0838_),
    .Y(_0841_)
  );
  \$_MUX_  _2725_ (
    .A(_0841_),
    .B(pc_sw[11]),
    .S(_0836_),
    .Y(_0002_[11])
  );
  \$_MUX_  _2726_ (
    .A(_0628_),
    .B(r12[12]),
    .S(_0838_),
    .Y(_0842_)
  );
  \$_MUX_  _2727_ (
    .A(_0842_),
    .B(pc_sw[12]),
    .S(_0836_),
    .Y(_0002_[12])
  );
  \$_MUX_  _2728_ (
    .A(_0632_),
    .B(r12[13]),
    .S(_0838_),
    .Y(_0843_)
  );
  \$_MUX_  _2729_ (
    .A(_0843_),
    .B(pc_sw[13]),
    .S(_0836_),
    .Y(_0002_[13])
  );
  \$_MUX_  _2730_ (
    .A(_0636_),
    .B(r12[14]),
    .S(_0838_),
    .Y(_0844_)
  );
  \$_MUX_  _2731_ (
    .A(_0844_),
    .B(pc_sw[14]),
    .S(_0836_),
    .Y(_0002_[14])
  );
  \$_MUX_  _2732_ (
    .A(_0640_),
    .B(r12[15]),
    .S(_0838_),
    .Y(_0845_)
  );
  \$_MUX_  _2733_ (
    .A(_0845_),
    .B(pc_sw[15]),
    .S(_0836_),
    .Y(_0002_[15])
  );
  \$_MUX_  _2734_ (
    .A(_0643_),
    .B(r12[1]),
    .S(_0838_),
    .Y(_0846_)
  );
  \$_MUX_  _2735_ (
    .A(_0846_),
    .B(reg_dest_val[1]),
    .S(_0836_),
    .Y(_0002_[1])
  );
  \$_MUX_  _2736_ (
    .A(_0646_),
    .B(r12[2]),
    .S(_0838_),
    .Y(_0847_)
  );
  \$_MUX_  _2737_ (
    .A(_0847_),
    .B(reg_dest_val[2]),
    .S(_0836_),
    .Y(_0002_[2])
  );
  \$_MUX_  _2738_ (
    .A(_0649_),
    .B(r12[3]),
    .S(_0838_),
    .Y(_0848_)
  );
  \$_MUX_  _2739_ (
    .A(_0848_),
    .B(reg_dest_val[3]),
    .S(_0836_),
    .Y(_0002_[3])
  );
  \$_MUX_  _2740_ (
    .A(_0652_),
    .B(r12[4]),
    .S(_0838_),
    .Y(_0849_)
  );
  \$_MUX_  _2741_ (
    .A(_0849_),
    .B(reg_dest_val[4]),
    .S(_0836_),
    .Y(_0002_[4])
  );
  \$_MUX_  _2742_ (
    .A(_0655_),
    .B(r12[5]),
    .S(_0838_),
    .Y(_0850_)
  );
  \$_MUX_  _2743_ (
    .A(_0850_),
    .B(reg_dest_val[5]),
    .S(_0836_),
    .Y(_0002_[5])
  );
  \$_MUX_  _2744_ (
    .A(_0658_),
    .B(r12[6]),
    .S(_0838_),
    .Y(_0851_)
  );
  \$_MUX_  _2745_ (
    .A(_0851_),
    .B(reg_dest_val[6]),
    .S(_0836_),
    .Y(_0002_[6])
  );
  \$_MUX_  _2746_ (
    .A(_0661_),
    .B(r12[7]),
    .S(_0838_),
    .Y(_0852_)
  );
  \$_MUX_  _2747_ (
    .A(_0852_),
    .B(reg_dest_val[7]),
    .S(_0836_),
    .Y(_0002_[7])
  );
  \$_MUX_  _2748_ (
    .A(_0664_),
    .B(r12[8]),
    .S(_0838_),
    .Y(_0853_)
  );
  \$_MUX_  _2749_ (
    .A(_0853_),
    .B(pc_sw[8]),
    .S(_0836_),
    .Y(_0002_[8])
  );
  \$_MUX_  _2750_ (
    .A(_0667_),
    .B(r12[9]),
    .S(_0838_),
    .Y(_0854_)
  );
  \$_MUX_  _2751_ (
    .A(_0854_),
    .B(pc_sw[9]),
    .S(_0836_),
    .Y(_0002_[9])
  );
  \$_AND_  _2752_ (
    .A(inst_dest[13]),
    .B(reg_dest_wr),
    .Y(_0855_)
  );
  \$_INV_  _2753_ (
    .A(_0929_),
    .Y(_0856_)
  );
  \$_OR_  _2754_ (
    .A(_0856_),
    .B(_0596_),
    .Y(_0857_)
  );
  \$_MUX_  _2755_ (
    .A(_0686_),
    .B(r13[0]),
    .S(_0857_),
    .Y(_0858_)
  );
  \$_MUX_  _2756_ (
    .A(_0858_),
    .B(reg_dest_val[0]),
    .S(_0855_),
    .Y(_0003_[0])
  );
  \$_MUX_  _2757_ (
    .A(_0620_),
    .B(r13[10]),
    .S(_0857_),
    .Y(_0859_)
  );
  \$_MUX_  _2758_ (
    .A(_0859_),
    .B(pc_sw[10]),
    .S(_0855_),
    .Y(_0003_[10])
  );
  \$_MUX_  _2759_ (
    .A(_0624_),
    .B(r13[11]),
    .S(_0857_),
    .Y(_0860_)
  );
  \$_MUX_  _2760_ (
    .A(_0860_),
    .B(pc_sw[11]),
    .S(_0855_),
    .Y(_0003_[11])
  );
  \$_MUX_  _2761_ (
    .A(_0628_),
    .B(r13[12]),
    .S(_0857_),
    .Y(_0861_)
  );
  \$_MUX_  _2762_ (
    .A(_0861_),
    .B(pc_sw[12]),
    .S(_0855_),
    .Y(_0003_[12])
  );
  \$_MUX_  _2763_ (
    .A(_0632_),
    .B(r13[13]),
    .S(_0857_),
    .Y(_0862_)
  );
  \$_MUX_  _2764_ (
    .A(_0862_),
    .B(pc_sw[13]),
    .S(_0855_),
    .Y(_0003_[13])
  );
  \$_MUX_  _2765_ (
    .A(_0636_),
    .B(r13[14]),
    .S(_0857_),
    .Y(_0863_)
  );
  \$_MUX_  _2766_ (
    .A(_0863_),
    .B(pc_sw[14]),
    .S(_0855_),
    .Y(_0003_[14])
  );
  \$_MUX_  _2767_ (
    .A(_0640_),
    .B(r13[15]),
    .S(_0857_),
    .Y(_0864_)
  );
  \$_MUX_  _2768_ (
    .A(_0864_),
    .B(pc_sw[15]),
    .S(_0855_),
    .Y(_0003_[15])
  );
  \$_MUX_  _2769_ (
    .A(_0643_),
    .B(r13[1]),
    .S(_0857_),
    .Y(_0865_)
  );
  \$_MUX_  _2770_ (
    .A(_0865_),
    .B(reg_dest_val[1]),
    .S(_0855_),
    .Y(_0003_[1])
  );
  \$_MUX_  _2771_ (
    .A(_0646_),
    .B(r13[2]),
    .S(_0857_),
    .Y(_0866_)
  );
  \$_MUX_  _2772_ (
    .A(_0866_),
    .B(reg_dest_val[2]),
    .S(_0855_),
    .Y(_0003_[2])
  );
  \$_MUX_  _2773_ (
    .A(_0649_),
    .B(r13[3]),
    .S(_0857_),
    .Y(_0867_)
  );
  \$_MUX_  _2774_ (
    .A(_0867_),
    .B(reg_dest_val[3]),
    .S(_0855_),
    .Y(_0003_[3])
  );
  \$_MUX_  _2775_ (
    .A(_0652_),
    .B(r13[4]),
    .S(_0857_),
    .Y(_0868_)
  );
  \$_MUX_  _2776_ (
    .A(_0868_),
    .B(reg_dest_val[4]),
    .S(_0855_),
    .Y(_0003_[4])
  );
  \$_MUX_  _2777_ (
    .A(_0655_),
    .B(r13[5]),
    .S(_0857_),
    .Y(_0869_)
  );
  \$_MUX_  _2778_ (
    .A(_0869_),
    .B(reg_dest_val[5]),
    .S(_0855_),
    .Y(_0003_[5])
  );
  \$_MUX_  _2779_ (
    .A(_0658_),
    .B(r13[6]),
    .S(_0857_),
    .Y(_0870_)
  );
  \$_MUX_  _2780_ (
    .A(_0870_),
    .B(reg_dest_val[6]),
    .S(_0855_),
    .Y(_0003_[6])
  );
  \$_MUX_  _2781_ (
    .A(_0661_),
    .B(r13[7]),
    .S(_0857_),
    .Y(_0871_)
  );
  \$_MUX_  _2782_ (
    .A(_0871_),
    .B(reg_dest_val[7]),
    .S(_0855_),
    .Y(_0003_[7])
  );
  \$_MUX_  _2783_ (
    .A(_0664_),
    .B(r13[8]),
    .S(_0857_),
    .Y(_0872_)
  );
  \$_MUX_  _2784_ (
    .A(_0872_),
    .B(pc_sw[8]),
    .S(_0855_),
    .Y(_0003_[8])
  );
  \$_MUX_  _2785_ (
    .A(_0667_),
    .B(r13[9]),
    .S(_0857_),
    .Y(_0873_)
  );
  \$_MUX_  _2786_ (
    .A(_0873_),
    .B(pc_sw[9]),
    .S(_0855_),
    .Y(_0003_[9])
  );
  \$_AND_  _2787_ (
    .A(inst_dest[14]),
    .B(reg_dest_wr),
    .Y(_0874_)
  );
  \$_INV_  _2788_ (
    .A(_0931_),
    .Y(_0875_)
  );
  \$_OR_  _2789_ (
    .A(_0875_),
    .B(_0596_),
    .Y(_0876_)
  );
  \$_MUX_  _2790_ (
    .A(_0686_),
    .B(r14[0]),
    .S(_0876_),
    .Y(_0877_)
  );
  \$_MUX_  _2791_ (
    .A(_0877_),
    .B(reg_dest_val[0]),
    .S(_0874_),
    .Y(_0004_[0])
  );
  \$_MUX_  _2792_ (
    .A(_0620_),
    .B(r14[10]),
    .S(_0876_),
    .Y(_0878_)
  );
  \$_MUX_  _2793_ (
    .A(_0878_),
    .B(pc_sw[10]),
    .S(_0874_),
    .Y(_0004_[10])
  );
  \$_MUX_  _2794_ (
    .A(_0624_),
    .B(r14[11]),
    .S(_0876_),
    .Y(_0879_)
  );
  \$_MUX_  _2795_ (
    .A(_0879_),
    .B(pc_sw[11]),
    .S(_0874_),
    .Y(_0004_[11])
  );
  \$_MUX_  _2796_ (
    .A(_0628_),
    .B(r14[12]),
    .S(_0876_),
    .Y(_0880_)
  );
  \$_MUX_  _2797_ (
    .A(_0880_),
    .B(pc_sw[12]),
    .S(_0874_),
    .Y(_0004_[12])
  );
  \$_MUX_  _2798_ (
    .A(_0632_),
    .B(r14[13]),
    .S(_0876_),
    .Y(_0881_)
  );
  \$_MUX_  _2799_ (
    .A(_0881_),
    .B(pc_sw[13]),
    .S(_0874_),
    .Y(_0004_[13])
  );
  \$_MUX_  _2800_ (
    .A(_0636_),
    .B(r14[14]),
    .S(_0876_),
    .Y(_0882_)
  );
  \$_MUX_  _2801_ (
    .A(_0882_),
    .B(pc_sw[14]),
    .S(_0874_),
    .Y(_0004_[14])
  );
  \$_MUX_  _2802_ (
    .A(_0640_),
    .B(r14[15]),
    .S(_0876_),
    .Y(_0883_)
  );
  \$_MUX_  _2803_ (
    .A(_0883_),
    .B(pc_sw[15]),
    .S(_0874_),
    .Y(_0004_[15])
  );
  \$_MUX_  _2804_ (
    .A(_0643_),
    .B(r14[1]),
    .S(_0876_),
    .Y(_0884_)
  );
  \$_MUX_  _2805_ (
    .A(_0884_),
    .B(reg_dest_val[1]),
    .S(_0874_),
    .Y(_0004_[1])
  );
  \$_MUX_  _2806_ (
    .A(_0646_),
    .B(r14[2]),
    .S(_0876_),
    .Y(_0885_)
  );
  \$_MUX_  _2807_ (
    .A(_0885_),
    .B(reg_dest_val[2]),
    .S(_0874_),
    .Y(_0004_[2])
  );
  \$_MUX_  _2808_ (
    .A(_0649_),
    .B(r14[3]),
    .S(_0876_),
    .Y(_0886_)
  );
  \$_MUX_  _2809_ (
    .A(_0886_),
    .B(reg_dest_val[3]),
    .S(_0874_),
    .Y(_0004_[3])
  );
  \$_MUX_  _2810_ (
    .A(_0652_),
    .B(r14[4]),
    .S(_0876_),
    .Y(_0887_)
  );
  \$_MUX_  _2811_ (
    .A(_0887_),
    .B(reg_dest_val[4]),
    .S(_0874_),
    .Y(_0004_[4])
  );
  \$_MUX_  _2812_ (
    .A(_0655_),
    .B(r14[5]),
    .S(_0876_),
    .Y(_0888_)
  );
  \$_MUX_  _2813_ (
    .A(_0888_),
    .B(reg_dest_val[5]),
    .S(_0874_),
    .Y(_0004_[5])
  );
  \$_MUX_  _2814_ (
    .A(_0658_),
    .B(r14[6]),
    .S(_0876_),
    .Y(_0889_)
  );
  \$_MUX_  _2815_ (
    .A(_0889_),
    .B(reg_dest_val[6]),
    .S(_0874_),
    .Y(_0004_[6])
  );
  \$_MUX_  _2816_ (
    .A(_0661_),
    .B(r14[7]),
    .S(_0876_),
    .Y(_0890_)
  );
  \$_MUX_  _2817_ (
    .A(_0890_),
    .B(reg_dest_val[7]),
    .S(_0874_),
    .Y(_0004_[7])
  );
  \$_MUX_  _2818_ (
    .A(_0664_),
    .B(r14[8]),
    .S(_0876_),
    .Y(_0891_)
  );
  \$_MUX_  _2819_ (
    .A(_0891_),
    .B(pc_sw[8]),
    .S(_0874_),
    .Y(_0004_[8])
  );
  \$_MUX_  _2820_ (
    .A(_0667_),
    .B(r14[9]),
    .S(_0876_),
    .Y(_0892_)
  );
  \$_MUX_  _2821_ (
    .A(_0892_),
    .B(pc_sw[9]),
    .S(_0874_),
    .Y(_0004_[9])
  );
  \$_AND_  _2822_ (
    .A(inst_dest[15]),
    .B(reg_dest_wr),
    .Y(_0893_)
  );
  \$_INV_  _2823_ (
    .A(_0927_),
    .Y(_0894_)
  );
  \$_OR_  _2824_ (
    .A(_0894_),
    .B(_0596_),
    .Y(_0895_)
  );
  \$_MUX_  _2825_ (
    .A(_0686_),
    .B(r15[0]),
    .S(_0895_),
    .Y(_0896_)
  );
  \$_MUX_  _2826_ (
    .A(_0896_),
    .B(reg_dest_val[0]),
    .S(_0893_),
    .Y(_0005_[0])
  );
  \$_MUX_  _2827_ (
    .A(_0620_),
    .B(r15[10]),
    .S(_0895_),
    .Y(_0897_)
  );
  \$_MUX_  _2828_ (
    .A(_0897_),
    .B(pc_sw[10]),
    .S(_0893_),
    .Y(_0005_[10])
  );
  \$_MUX_  _2829_ (
    .A(_0624_),
    .B(r15[11]),
    .S(_0895_),
    .Y(_0898_)
  );
  \$_MUX_  _2830_ (
    .A(_0898_),
    .B(pc_sw[11]),
    .S(_0893_),
    .Y(_0005_[11])
  );
  \$_MUX_  _2831_ (
    .A(_0628_),
    .B(r15[12]),
    .S(_0895_),
    .Y(_0899_)
  );
  \$_MUX_  _2832_ (
    .A(_0899_),
    .B(pc_sw[12]),
    .S(_0893_),
    .Y(_0005_[12])
  );
  \$_MUX_  _2833_ (
    .A(_0632_),
    .B(r15[13]),
    .S(_0895_),
    .Y(_0900_)
  );
  \$_MUX_  _2834_ (
    .A(_0900_),
    .B(pc_sw[13]),
    .S(_0893_),
    .Y(_0005_[13])
  );
  \$_MUX_  _2835_ (
    .A(_0636_),
    .B(r15[14]),
    .S(_0895_),
    .Y(_0901_)
  );
  \$_MUX_  _2836_ (
    .A(_0901_),
    .B(pc_sw[14]),
    .S(_0893_),
    .Y(_0005_[14])
  );
  \$_MUX_  _2837_ (
    .A(_0640_),
    .B(r15[15]),
    .S(_0895_),
    .Y(_0902_)
  );
  \$_MUX_  _2838_ (
    .A(_0902_),
    .B(pc_sw[15]),
    .S(_0893_),
    .Y(_0005_[15])
  );
  \$_MUX_  _2839_ (
    .A(_0643_),
    .B(r15[1]),
    .S(_0895_),
    .Y(_0903_)
  );
  \$_MUX_  _2840_ (
    .A(_0903_),
    .B(reg_dest_val[1]),
    .S(_0893_),
    .Y(_0005_[1])
  );
  \$_MUX_  _2841_ (
    .A(_0646_),
    .B(r15[2]),
    .S(_0895_),
    .Y(_0904_)
  );
  \$_MUX_  _2842_ (
    .A(_0904_),
    .B(reg_dest_val[2]),
    .S(_0893_),
    .Y(_0005_[2])
  );
  \$_MUX_  _2843_ (
    .A(_0649_),
    .B(r15[3]),
    .S(_0895_),
    .Y(_0905_)
  );
  \$_MUX_  _2844_ (
    .A(_0905_),
    .B(reg_dest_val[3]),
    .S(_0893_),
    .Y(_0005_[3])
  );
  \$_MUX_  _2845_ (
    .A(_0652_),
    .B(r15[4]),
    .S(_0895_),
    .Y(_0906_)
  );
  \$_MUX_  _2846_ (
    .A(_0906_),
    .B(reg_dest_val[4]),
    .S(_0893_),
    .Y(_0005_[4])
  );
  \$_MUX_  _2847_ (
    .A(_0655_),
    .B(r15[5]),
    .S(_0895_),
    .Y(_0907_)
  );
  \$_MUX_  _2848_ (
    .A(_0907_),
    .B(reg_dest_val[5]),
    .S(_0893_),
    .Y(_0005_[5])
  );
  \$_MUX_  _2849_ (
    .A(_0658_),
    .B(r15[6]),
    .S(_0895_),
    .Y(_0908_)
  );
  \$_MUX_  _2850_ (
    .A(_0908_),
    .B(reg_dest_val[6]),
    .S(_0893_),
    .Y(_0005_[6])
  );
  \$_MUX_  _2851_ (
    .A(_0661_),
    .B(r15[7]),
    .S(_0895_),
    .Y(_0909_)
  );
  \$_MUX_  _2852_ (
    .A(_0909_),
    .B(reg_dest_val[7]),
    .S(_0893_),
    .Y(_0005_[7])
  );
  \$_MUX_  _2853_ (
    .A(_0664_),
    .B(r15[8]),
    .S(_0895_),
    .Y(_0910_)
  );
  \$_MUX_  _2854_ (
    .A(_0910_),
    .B(pc_sw[8]),
    .S(_0893_),
    .Y(_0005_[8])
  );
  \$_MUX_  _2855_ (
    .A(_0667_),
    .B(r15[9]),
    .S(_0895_),
    .Y(_0911_)
  );
  \$_MUX_  _2856_ (
    .A(_0911_),
    .B(pc_sw[9]),
    .S(_0893_),
    .Y(_0005_[9])
  );
  \$_DFF_PP0_  \r1_reg[0]  /* _2857_ */ (
    .C(mclk),
    .D(_0006_[0]),
    .Q(r1[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[10]  /* _2858_ */ (
    .C(mclk),
    .D(_0006_[10]),
    .Q(r1[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[11]  /* _2859_ */ (
    .C(mclk),
    .D(_0006_[11]),
    .Q(r1[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[12]  /* _2860_ */ (
    .C(mclk),
    .D(_0006_[12]),
    .Q(r1[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[13]  /* _2861_ */ (
    .C(mclk),
    .D(_0006_[13]),
    .Q(r1[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[14]  /* _2862_ */ (
    .C(mclk),
    .D(_0006_[14]),
    .Q(r1[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[15]  /* _2863_ */ (
    .C(mclk),
    .D(_0006_[15]),
    .Q(r1[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[1]  /* _2864_ */ (
    .C(mclk),
    .D(_0006_[1]),
    .Q(r1[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[2]  /* _2865_ */ (
    .C(mclk),
    .D(_0006_[2]),
    .Q(r1[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[3]  /* _2866_ */ (
    .C(mclk),
    .D(_0006_[3]),
    .Q(r1[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[4]  /* _2867_ */ (
    .C(mclk),
    .D(_0006_[4]),
    .Q(r1[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[5]  /* _2868_ */ (
    .C(mclk),
    .D(_0006_[5]),
    .Q(r1[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[6]  /* _2869_ */ (
    .C(mclk),
    .D(_0006_[6]),
    .Q(r1[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[7]  /* _2870_ */ (
    .C(mclk),
    .D(_0006_[7]),
    .Q(r1[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[8]  /* _2871_ */ (
    .C(mclk),
    .D(_0006_[8]),
    .Q(r1[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r1_reg[9]  /* _2872_ */ (
    .C(mclk),
    .D(_0006_[9]),
    .Q(r1[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[0]  /* _2873_ */ (
    .C(mclk),
    .D(_0007_[0]),
    .Q(r2[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[15]  /* _2874_ */ (
    .C(mclk),
    .D(1'b0),
    .Q(r2[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[1]  /* _2875_ */ (
    .C(mclk),
    .D(_0007_[1]),
    .Q(r2[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[2]  /* _2876_ */ (
    .C(mclk),
    .D(_0007_[2]),
    .Q(r2[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  gie_reg /* _2877_ */ (
    .C(mclk),
    .D(_0007_[3]),
    .Q(gie),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[4]  /* _2878_ */ (
    .C(mclk),
    .D(_0007_[4]),
    .Q(r2[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  oscoff_reg /* _2879_ */ (
    .C(mclk),
    .D(_0007_[5]),
    .Q(oscoff),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[7]  /* _2880_ */ (
    .C(mclk),
    .D(_0007_[7]),
    .Q(r2[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r2_reg[8]  /* _2881_ */ (
    .C(mclk),
    .D(_0007_[8]),
    .Q(r2[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[0]  /* _2882_ */ (
    .C(mclk),
    .D(_0008_[0]),
    .Q(r3[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[10]  /* _2883_ */ (
    .C(mclk),
    .D(_0008_[10]),
    .Q(r3[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[11]  /* _2884_ */ (
    .C(mclk),
    .D(_0008_[11]),
    .Q(r3[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[12]  /* _2885_ */ (
    .C(mclk),
    .D(_0008_[12]),
    .Q(r3[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[13]  /* _2886_ */ (
    .C(mclk),
    .D(_0008_[13]),
    .Q(r3[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[14]  /* _2887_ */ (
    .C(mclk),
    .D(_0008_[14]),
    .Q(r3[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[15]  /* _2888_ */ (
    .C(mclk),
    .D(_0008_[15]),
    .Q(r3[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[1]  /* _2889_ */ (
    .C(mclk),
    .D(_0008_[1]),
    .Q(r3[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[2]  /* _2890_ */ (
    .C(mclk),
    .D(_0008_[2]),
    .Q(r3[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[3]  /* _2891_ */ (
    .C(mclk),
    .D(_0008_[3]),
    .Q(r3[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[4]  /* _2892_ */ (
    .C(mclk),
    .D(_0008_[4]),
    .Q(r3[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[5]  /* _2893_ */ (
    .C(mclk),
    .D(_0008_[5]),
    .Q(r3[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[6]  /* _2894_ */ (
    .C(mclk),
    .D(_0008_[6]),
    .Q(r3[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[7]  /* _2895_ */ (
    .C(mclk),
    .D(_0008_[7]),
    .Q(r3[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[8]  /* _2896_ */ (
    .C(mclk),
    .D(_0008_[8]),
    .Q(r3[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r3_reg[9]  /* _2897_ */ (
    .C(mclk),
    .D(_0008_[9]),
    .Q(r3[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[0]  /* _2898_ */ (
    .C(mclk),
    .D(_0009_[0]),
    .Q(r4[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[10]  /* _2899_ */ (
    .C(mclk),
    .D(_0009_[10]),
    .Q(r4[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[11]  /* _2900_ */ (
    .C(mclk),
    .D(_0009_[11]),
    .Q(r4[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[12]  /* _2901_ */ (
    .C(mclk),
    .D(_0009_[12]),
    .Q(r4[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[13]  /* _2902_ */ (
    .C(mclk),
    .D(_0009_[13]),
    .Q(r4[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[14]  /* _2903_ */ (
    .C(mclk),
    .D(_0009_[14]),
    .Q(r4[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[15]  /* _2904_ */ (
    .C(mclk),
    .D(_0009_[15]),
    .Q(r4[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[1]  /* _2905_ */ (
    .C(mclk),
    .D(_0009_[1]),
    .Q(r4[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[2]  /* _2906_ */ (
    .C(mclk),
    .D(_0009_[2]),
    .Q(r4[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[3]  /* _2907_ */ (
    .C(mclk),
    .D(_0009_[3]),
    .Q(r4[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[4]  /* _2908_ */ (
    .C(mclk),
    .D(_0009_[4]),
    .Q(r4[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[5]  /* _2909_ */ (
    .C(mclk),
    .D(_0009_[5]),
    .Q(r4[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[6]  /* _2910_ */ (
    .C(mclk),
    .D(_0009_[6]),
    .Q(r4[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[7]  /* _2911_ */ (
    .C(mclk),
    .D(_0009_[7]),
    .Q(r4[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[8]  /* _2912_ */ (
    .C(mclk),
    .D(_0009_[8]),
    .Q(r4[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r4_reg[9]  /* _2913_ */ (
    .C(mclk),
    .D(_0009_[9]),
    .Q(r4[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[0]  /* _2914_ */ (
    .C(mclk),
    .D(_0010_[0]),
    .Q(r5[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[10]  /* _2915_ */ (
    .C(mclk),
    .D(_0010_[10]),
    .Q(r5[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[11]  /* _2916_ */ (
    .C(mclk),
    .D(_0010_[11]),
    .Q(r5[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[12]  /* _2917_ */ (
    .C(mclk),
    .D(_0010_[12]),
    .Q(r5[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[13]  /* _2918_ */ (
    .C(mclk),
    .D(_0010_[13]),
    .Q(r5[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[14]  /* _2919_ */ (
    .C(mclk),
    .D(_0010_[14]),
    .Q(r5[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[15]  /* _2920_ */ (
    .C(mclk),
    .D(_0010_[15]),
    .Q(r5[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[1]  /* _2921_ */ (
    .C(mclk),
    .D(_0010_[1]),
    .Q(r5[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[2]  /* _2922_ */ (
    .C(mclk),
    .D(_0010_[2]),
    .Q(r5[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[3]  /* _2923_ */ (
    .C(mclk),
    .D(_0010_[3]),
    .Q(r5[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[4]  /* _2924_ */ (
    .C(mclk),
    .D(_0010_[4]),
    .Q(r5[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[5]  /* _2925_ */ (
    .C(mclk),
    .D(_0010_[5]),
    .Q(r5[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[6]  /* _2926_ */ (
    .C(mclk),
    .D(_0010_[6]),
    .Q(r5[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[7]  /* _2927_ */ (
    .C(mclk),
    .D(_0010_[7]),
    .Q(r5[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[8]  /* _2928_ */ (
    .C(mclk),
    .D(_0010_[8]),
    .Q(r5[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r5_reg[9]  /* _2929_ */ (
    .C(mclk),
    .D(_0010_[9]),
    .Q(r5[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[0]  /* _2930_ */ (
    .C(mclk),
    .D(_0011_[0]),
    .Q(r6[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[10]  /* _2931_ */ (
    .C(mclk),
    .D(_0011_[10]),
    .Q(r6[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[11]  /* _2932_ */ (
    .C(mclk),
    .D(_0011_[11]),
    .Q(r6[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[12]  /* _2933_ */ (
    .C(mclk),
    .D(_0011_[12]),
    .Q(r6[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[13]  /* _2934_ */ (
    .C(mclk),
    .D(_0011_[13]),
    .Q(r6[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[14]  /* _2935_ */ (
    .C(mclk),
    .D(_0011_[14]),
    .Q(r6[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[15]  /* _2936_ */ (
    .C(mclk),
    .D(_0011_[15]),
    .Q(r6[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[1]  /* _2937_ */ (
    .C(mclk),
    .D(_0011_[1]),
    .Q(r6[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[2]  /* _2938_ */ (
    .C(mclk),
    .D(_0011_[2]),
    .Q(r6[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[3]  /* _2939_ */ (
    .C(mclk),
    .D(_0011_[3]),
    .Q(r6[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[4]  /* _2940_ */ (
    .C(mclk),
    .D(_0011_[4]),
    .Q(r6[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[5]  /* _2941_ */ (
    .C(mclk),
    .D(_0011_[5]),
    .Q(r6[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[6]  /* _2942_ */ (
    .C(mclk),
    .D(_0011_[6]),
    .Q(r6[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[7]  /* _2943_ */ (
    .C(mclk),
    .D(_0011_[7]),
    .Q(r6[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[8]  /* _2944_ */ (
    .C(mclk),
    .D(_0011_[8]),
    .Q(r6[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r6_reg[9]  /* _2945_ */ (
    .C(mclk),
    .D(_0011_[9]),
    .Q(r6[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[0]  /* _2946_ */ (
    .C(mclk),
    .D(_0012_[0]),
    .Q(r7[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[10]  /* _2947_ */ (
    .C(mclk),
    .D(_0012_[10]),
    .Q(r7[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[11]  /* _2948_ */ (
    .C(mclk),
    .D(_0012_[11]),
    .Q(r7[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[12]  /* _2949_ */ (
    .C(mclk),
    .D(_0012_[12]),
    .Q(r7[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[13]  /* _2950_ */ (
    .C(mclk),
    .D(_0012_[13]),
    .Q(r7[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[14]  /* _2951_ */ (
    .C(mclk),
    .D(_0012_[14]),
    .Q(r7[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[15]  /* _2952_ */ (
    .C(mclk),
    .D(_0012_[15]),
    .Q(r7[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[1]  /* _2953_ */ (
    .C(mclk),
    .D(_0012_[1]),
    .Q(r7[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[2]  /* _2954_ */ (
    .C(mclk),
    .D(_0012_[2]),
    .Q(r7[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[3]  /* _2955_ */ (
    .C(mclk),
    .D(_0012_[3]),
    .Q(r7[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[4]  /* _2956_ */ (
    .C(mclk),
    .D(_0012_[4]),
    .Q(r7[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[5]  /* _2957_ */ (
    .C(mclk),
    .D(_0012_[5]),
    .Q(r7[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[6]  /* _2958_ */ (
    .C(mclk),
    .D(_0012_[6]),
    .Q(r7[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[7]  /* _2959_ */ (
    .C(mclk),
    .D(_0012_[7]),
    .Q(r7[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[8]  /* _2960_ */ (
    .C(mclk),
    .D(_0012_[8]),
    .Q(r7[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r7_reg[9]  /* _2961_ */ (
    .C(mclk),
    .D(_0012_[9]),
    .Q(r7[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[0]  /* _2962_ */ (
    .C(mclk),
    .D(_0013_[0]),
    .Q(r8[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[10]  /* _2963_ */ (
    .C(mclk),
    .D(_0013_[10]),
    .Q(r8[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[11]  /* _2964_ */ (
    .C(mclk),
    .D(_0013_[11]),
    .Q(r8[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[12]  /* _2965_ */ (
    .C(mclk),
    .D(_0013_[12]),
    .Q(r8[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[13]  /* _2966_ */ (
    .C(mclk),
    .D(_0013_[13]),
    .Q(r8[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[14]  /* _2967_ */ (
    .C(mclk),
    .D(_0013_[14]),
    .Q(r8[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[15]  /* _2968_ */ (
    .C(mclk),
    .D(_0013_[15]),
    .Q(r8[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[1]  /* _2969_ */ (
    .C(mclk),
    .D(_0013_[1]),
    .Q(r8[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[2]  /* _2970_ */ (
    .C(mclk),
    .D(_0013_[2]),
    .Q(r8[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[3]  /* _2971_ */ (
    .C(mclk),
    .D(_0013_[3]),
    .Q(r8[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[4]  /* _2972_ */ (
    .C(mclk),
    .D(_0013_[4]),
    .Q(r8[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[5]  /* _2973_ */ (
    .C(mclk),
    .D(_0013_[5]),
    .Q(r8[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[6]  /* _2974_ */ (
    .C(mclk),
    .D(_0013_[6]),
    .Q(r8[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[7]  /* _2975_ */ (
    .C(mclk),
    .D(_0013_[7]),
    .Q(r8[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[8]  /* _2976_ */ (
    .C(mclk),
    .D(_0013_[8]),
    .Q(r8[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r8_reg[9]  /* _2977_ */ (
    .C(mclk),
    .D(_0013_[9]),
    .Q(r8[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[0]  /* _2978_ */ (
    .C(mclk),
    .D(_0014_[0]),
    .Q(r9[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[10]  /* _2979_ */ (
    .C(mclk),
    .D(_0014_[10]),
    .Q(r9[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[11]  /* _2980_ */ (
    .C(mclk),
    .D(_0014_[11]),
    .Q(r9[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[12]  /* _2981_ */ (
    .C(mclk),
    .D(_0014_[12]),
    .Q(r9[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[13]  /* _2982_ */ (
    .C(mclk),
    .D(_0014_[13]),
    .Q(r9[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[14]  /* _2983_ */ (
    .C(mclk),
    .D(_0014_[14]),
    .Q(r9[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[15]  /* _2984_ */ (
    .C(mclk),
    .D(_0014_[15]),
    .Q(r9[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[1]  /* _2985_ */ (
    .C(mclk),
    .D(_0014_[1]),
    .Q(r9[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[2]  /* _2986_ */ (
    .C(mclk),
    .D(_0014_[2]),
    .Q(r9[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[3]  /* _2987_ */ (
    .C(mclk),
    .D(_0014_[3]),
    .Q(r9[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[4]  /* _2988_ */ (
    .C(mclk),
    .D(_0014_[4]),
    .Q(r9[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[5]  /* _2989_ */ (
    .C(mclk),
    .D(_0014_[5]),
    .Q(r9[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[6]  /* _2990_ */ (
    .C(mclk),
    .D(_0014_[6]),
    .Q(r9[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[7]  /* _2991_ */ (
    .C(mclk),
    .D(_0014_[7]),
    .Q(r9[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[8]  /* _2992_ */ (
    .C(mclk),
    .D(_0014_[8]),
    .Q(r9[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r9_reg[9]  /* _2993_ */ (
    .C(mclk),
    .D(_0014_[9]),
    .Q(r9[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[0]  /* _2994_ */ (
    .C(mclk),
    .D(_0000_[0]),
    .Q(r10[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[10]  /* _2995_ */ (
    .C(mclk),
    .D(_0000_[10]),
    .Q(r10[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[11]  /* _2996_ */ (
    .C(mclk),
    .D(_0000_[11]),
    .Q(r10[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[12]  /* _2997_ */ (
    .C(mclk),
    .D(_0000_[12]),
    .Q(r10[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[13]  /* _2998_ */ (
    .C(mclk),
    .D(_0000_[13]),
    .Q(r10[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[14]  /* _2999_ */ (
    .C(mclk),
    .D(_0000_[14]),
    .Q(r10[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[15]  /* _3000_ */ (
    .C(mclk),
    .D(_0000_[15]),
    .Q(r10[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[1]  /* _3001_ */ (
    .C(mclk),
    .D(_0000_[1]),
    .Q(r10[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[2]  /* _3002_ */ (
    .C(mclk),
    .D(_0000_[2]),
    .Q(r10[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[3]  /* _3003_ */ (
    .C(mclk),
    .D(_0000_[3]),
    .Q(r10[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[4]  /* _3004_ */ (
    .C(mclk),
    .D(_0000_[4]),
    .Q(r10[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[5]  /* _3005_ */ (
    .C(mclk),
    .D(_0000_[5]),
    .Q(r10[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[6]  /* _3006_ */ (
    .C(mclk),
    .D(_0000_[6]),
    .Q(r10[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[7]  /* _3007_ */ (
    .C(mclk),
    .D(_0000_[7]),
    .Q(r10[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[8]  /* _3008_ */ (
    .C(mclk),
    .D(_0000_[8]),
    .Q(r10[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r10_reg[9]  /* _3009_ */ (
    .C(mclk),
    .D(_0000_[9]),
    .Q(r10[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[0]  /* _3010_ */ (
    .C(mclk),
    .D(_0001_[0]),
    .Q(r11[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[10]  /* _3011_ */ (
    .C(mclk),
    .D(_0001_[10]),
    .Q(r11[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[11]  /* _3012_ */ (
    .C(mclk),
    .D(_0001_[11]),
    .Q(r11[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[12]  /* _3013_ */ (
    .C(mclk),
    .D(_0001_[12]),
    .Q(r11[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[13]  /* _3014_ */ (
    .C(mclk),
    .D(_0001_[13]),
    .Q(r11[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[14]  /* _3015_ */ (
    .C(mclk),
    .D(_0001_[14]),
    .Q(r11[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[15]  /* _3016_ */ (
    .C(mclk),
    .D(_0001_[15]),
    .Q(r11[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[1]  /* _3017_ */ (
    .C(mclk),
    .D(_0001_[1]),
    .Q(r11[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[2]  /* _3018_ */ (
    .C(mclk),
    .D(_0001_[2]),
    .Q(r11[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[3]  /* _3019_ */ (
    .C(mclk),
    .D(_0001_[3]),
    .Q(r11[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[4]  /* _3020_ */ (
    .C(mclk),
    .D(_0001_[4]),
    .Q(r11[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[5]  /* _3021_ */ (
    .C(mclk),
    .D(_0001_[5]),
    .Q(r11[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[6]  /* _3022_ */ (
    .C(mclk),
    .D(_0001_[6]),
    .Q(r11[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[7]  /* _3023_ */ (
    .C(mclk),
    .D(_0001_[7]),
    .Q(r11[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[8]  /* _3024_ */ (
    .C(mclk),
    .D(_0001_[8]),
    .Q(r11[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r11_reg[9]  /* _3025_ */ (
    .C(mclk),
    .D(_0001_[9]),
    .Q(r11[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[0]  /* _3026_ */ (
    .C(mclk),
    .D(_0002_[0]),
    .Q(r12[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[10]  /* _3027_ */ (
    .C(mclk),
    .D(_0002_[10]),
    .Q(r12[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[11]  /* _3028_ */ (
    .C(mclk),
    .D(_0002_[11]),
    .Q(r12[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[12]  /* _3029_ */ (
    .C(mclk),
    .D(_0002_[12]),
    .Q(r12[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[13]  /* _3030_ */ (
    .C(mclk),
    .D(_0002_[13]),
    .Q(r12[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[14]  /* _3031_ */ (
    .C(mclk),
    .D(_0002_[14]),
    .Q(r12[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[15]  /* _3032_ */ (
    .C(mclk),
    .D(_0002_[15]),
    .Q(r12[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[1]  /* _3033_ */ (
    .C(mclk),
    .D(_0002_[1]),
    .Q(r12[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[2]  /* _3034_ */ (
    .C(mclk),
    .D(_0002_[2]),
    .Q(r12[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[3]  /* _3035_ */ (
    .C(mclk),
    .D(_0002_[3]),
    .Q(r12[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[4]  /* _3036_ */ (
    .C(mclk),
    .D(_0002_[4]),
    .Q(r12[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[5]  /* _3037_ */ (
    .C(mclk),
    .D(_0002_[5]),
    .Q(r12[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[6]  /* _3038_ */ (
    .C(mclk),
    .D(_0002_[6]),
    .Q(r12[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[7]  /* _3039_ */ (
    .C(mclk),
    .D(_0002_[7]),
    .Q(r12[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[8]  /* _3040_ */ (
    .C(mclk),
    .D(_0002_[8]),
    .Q(r12[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r12_reg[9]  /* _3041_ */ (
    .C(mclk),
    .D(_0002_[9]),
    .Q(r12[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[0]  /* _3042_ */ (
    .C(mclk),
    .D(_0003_[0]),
    .Q(r13[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[10]  /* _3043_ */ (
    .C(mclk),
    .D(_0003_[10]),
    .Q(r13[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[11]  /* _3044_ */ (
    .C(mclk),
    .D(_0003_[11]),
    .Q(r13[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[12]  /* _3045_ */ (
    .C(mclk),
    .D(_0003_[12]),
    .Q(r13[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[13]  /* _3046_ */ (
    .C(mclk),
    .D(_0003_[13]),
    .Q(r13[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[14]  /* _3047_ */ (
    .C(mclk),
    .D(_0003_[14]),
    .Q(r13[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[15]  /* _3048_ */ (
    .C(mclk),
    .D(_0003_[15]),
    .Q(r13[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[1]  /* _3049_ */ (
    .C(mclk),
    .D(_0003_[1]),
    .Q(r13[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[2]  /* _3050_ */ (
    .C(mclk),
    .D(_0003_[2]),
    .Q(r13[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[3]  /* _3051_ */ (
    .C(mclk),
    .D(_0003_[3]),
    .Q(r13[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[4]  /* _3052_ */ (
    .C(mclk),
    .D(_0003_[4]),
    .Q(r13[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[5]  /* _3053_ */ (
    .C(mclk),
    .D(_0003_[5]),
    .Q(r13[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[6]  /* _3054_ */ (
    .C(mclk),
    .D(_0003_[6]),
    .Q(r13[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[7]  /* _3055_ */ (
    .C(mclk),
    .D(_0003_[7]),
    .Q(r13[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[8]  /* _3056_ */ (
    .C(mclk),
    .D(_0003_[8]),
    .Q(r13[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r13_reg[9]  /* _3057_ */ (
    .C(mclk),
    .D(_0003_[9]),
    .Q(r13[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[0]  /* _3058_ */ (
    .C(mclk),
    .D(_0004_[0]),
    .Q(r14[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[10]  /* _3059_ */ (
    .C(mclk),
    .D(_0004_[10]),
    .Q(r14[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[11]  /* _3060_ */ (
    .C(mclk),
    .D(_0004_[11]),
    .Q(r14[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[12]  /* _3061_ */ (
    .C(mclk),
    .D(_0004_[12]),
    .Q(r14[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[13]  /* _3062_ */ (
    .C(mclk),
    .D(_0004_[13]),
    .Q(r14[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[14]  /* _3063_ */ (
    .C(mclk),
    .D(_0004_[14]),
    .Q(r14[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[15]  /* _3064_ */ (
    .C(mclk),
    .D(_0004_[15]),
    .Q(r14[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[1]  /* _3065_ */ (
    .C(mclk),
    .D(_0004_[1]),
    .Q(r14[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[2]  /* _3066_ */ (
    .C(mclk),
    .D(_0004_[2]),
    .Q(r14[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[3]  /* _3067_ */ (
    .C(mclk),
    .D(_0004_[3]),
    .Q(r14[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[4]  /* _3068_ */ (
    .C(mclk),
    .D(_0004_[4]),
    .Q(r14[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[5]  /* _3069_ */ (
    .C(mclk),
    .D(_0004_[5]),
    .Q(r14[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[6]  /* _3070_ */ (
    .C(mclk),
    .D(_0004_[6]),
    .Q(r14[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[7]  /* _3071_ */ (
    .C(mclk),
    .D(_0004_[7]),
    .Q(r14[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[8]  /* _3072_ */ (
    .C(mclk),
    .D(_0004_[8]),
    .Q(r14[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r14_reg[9]  /* _3073_ */ (
    .C(mclk),
    .D(_0004_[9]),
    .Q(r14[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[0]  /* _3074_ */ (
    .C(mclk),
    .D(_0005_[0]),
    .Q(r15[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[10]  /* _3075_ */ (
    .C(mclk),
    .D(_0005_[10]),
    .Q(r15[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[11]  /* _3076_ */ (
    .C(mclk),
    .D(_0005_[11]),
    .Q(r15[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[12]  /* _3077_ */ (
    .C(mclk),
    .D(_0005_[12]),
    .Q(r15[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[13]  /* _3078_ */ (
    .C(mclk),
    .D(_0005_[13]),
    .Q(r15[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[14]  /* _3079_ */ (
    .C(mclk),
    .D(_0005_[14]),
    .Q(r15[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[15]  /* _3080_ */ (
    .C(mclk),
    .D(_0005_[15]),
    .Q(r15[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[1]  /* _3081_ */ (
    .C(mclk),
    .D(_0005_[1]),
    .Q(r15[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[2]  /* _3082_ */ (
    .C(mclk),
    .D(_0005_[2]),
    .Q(r15[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[3]  /* _3083_ */ (
    .C(mclk),
    .D(_0005_[3]),
    .Q(r15[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[4]  /* _3084_ */ (
    .C(mclk),
    .D(_0005_[4]),
    .Q(r15[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[5]  /* _3085_ */ (
    .C(mclk),
    .D(_0005_[5]),
    .Q(r15[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[6]  /* _3086_ */ (
    .C(mclk),
    .D(_0005_[6]),
    .Q(r15[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[7]  /* _3087_ */ (
    .C(mclk),
    .D(_0005_[7]),
    .Q(r15[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[8]  /* _3088_ */ (
    .C(mclk),
    .D(_0005_[8]),
    .Q(r15[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \r15_reg[9]  /* _3089_ */ (
    .C(mclk),
    .D(_0005_[9]),
    .Q(r15[9]),
    .R(puc_rst)
  );
  assign mclk_r1 = mclk;
  assign mclk_r10 = mclk;
  assign mclk_r11 = mclk;
  assign mclk_r12 = mclk;
  assign mclk_r13 = mclk;
  assign mclk_r14 = mclk;
  assign mclk_r15 = mclk;
  assign mclk_r2 = mclk;
  assign mclk_r3 = mclk;
  assign mclk_r4 = mclk;
  assign mclk_r5 = mclk;
  assign mclk_r6 = mclk;
  assign mclk_r7 = mclk;
  assign mclk_r8 = mclk;
  assign mclk_r9 = mclk;
  assign pc_sw[7:0] = reg_dest_val[7:0];
  assign r0 = pc;
  assign { r2[14:9], r2[6:5], r2[3] } = { r2[15], r2[15], r2[15], r2[15], r2[15], r2[15], r2[15], oscoff, gie };
  assign reg_dest_val_in = { pc_sw[15:8], reg_dest_val[7:0] };
  assign scg0 = r2[15];
  assign scg1 = r2[7];
  assign status = { r2[8], r2[2:0] };
endmodule

module omsp_sfr(cpu_id, nmi_pnd, nmi_wkup, per_dout, wdtie, wdtifg_sw_clr, wdtifg_sw_set, mclk, nmi, nmi_acc, per_addr, per_din, per_en, per_we, puc_rst, scan_mode, wdtifg, wdtnmies);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  output [31:0] cpu_id;
  wire [15:0] cpu_id_hi_rd;
  wire [15:0] cpu_id_lo_rd;
  wire [7:0] ie1;
  wire [7:0] ie1_nxt;
  wire [7:0] ifg1;
  wire [7:0] ifg1_nxt;
  input mclk;
  input nmi;
  input nmi_acc;
  wire nmi_capture;
  wire nmi_dly;
  output nmi_pnd;
  wire nmi_pol;
  wire nmi_s;
  output nmi_wkup;
  wire nmie;
  wire nmiifg;
  input [13:0] per_addr;
  input [15:0] per_din;
  output [15:0] per_dout;
  input per_en;
  input [1:0] per_we;
  input puc_rst;
  wire [2:0] reg_addr;
  wire [7:0] reg_rd;
  input scan_mode;
  output wdtie;
  input wdtifg;
  output wdtifg_sw_clr;
  output wdtifg_sw_set;
  input wdtnmies;
  \$_INV_  _067_ (
    .A(per_addr[12]),
    .Y(_015_)
  );
  \$_AND_  _068_ (
    .A(_015_),
    .B(per_en),
    .Y(_016_)
  );
  \$_INV_  _069_ (
    .A(per_addr[13]),
    .Y(_017_)
  );
  \$_INV_  _070_ (
    .A(per_addr[2]),
    .Y(_018_)
  );
  \$_AND_  _071_ (
    .A(_018_),
    .B(_017_),
    .Y(_019_)
  );
  \$_INV_  _072_ (
    .A(per_addr[3]),
    .Y(_020_)
  );
  \$_INV_  _073_ (
    .A(per_addr[4]),
    .Y(_021_)
  );
  \$_AND_  _074_ (
    .A(_021_),
    .B(_020_),
    .Y(_022_)
  );
  \$_AND_  _075_ (
    .A(_022_),
    .B(_019_),
    .Y(_023_)
  );
  \$_AND_  _076_ (
    .A(_023_),
    .B(_016_),
    .Y(_024_)
  );
  \$_INV_  _077_ (
    .A(per_addr[11]),
    .Y(_025_)
  );
  \$_INV_  _078_ (
    .A(per_addr[9]),
    .Y(_026_)
  );
  \$_INV_  _079_ (
    .A(per_addr[10]),
    .Y(_027_)
  );
  \$_AND_  _080_ (
    .A(_027_),
    .B(_026_),
    .Y(_028_)
  );
  \$_AND_  _081_ (
    .A(_028_),
    .B(_025_),
    .Y(_029_)
  );
  \$_INV_  _082_ (
    .A(per_addr[5]),
    .Y(_030_)
  );
  \$_INV_  _083_ (
    .A(per_addr[6]),
    .Y(_031_)
  );
  \$_AND_  _084_ (
    .A(_031_),
    .B(_030_),
    .Y(_032_)
  );
  \$_INV_  _085_ (
    .A(per_addr[7]),
    .Y(_033_)
  );
  \$_INV_  _086_ (
    .A(per_addr[8]),
    .Y(_034_)
  );
  \$_AND_  _087_ (
    .A(_034_),
    .B(_033_),
    .Y(_035_)
  );
  \$_AND_  _088_ (
    .A(_035_),
    .B(_032_),
    .Y(_036_)
  );
  \$_AND_  _089_ (
    .A(_036_),
    .B(_029_),
    .Y(_037_)
  );
  \$_AND_  _090_ (
    .A(_037_),
    .B(_024_),
    .Y(_038_)
  );
  \$_INV_  _091_ (
    .A(per_we[0]),
    .Y(_039_)
  );
  \$_INV_  _092_ (
    .A(per_we[1]),
    .Y(_040_)
  );
  \$_AND_  _093_ (
    .A(_040_),
    .B(_039_),
    .Y(_041_)
  );
  \$_AND_  _094_ (
    .A(_041_),
    .B(_038_),
    .Y(_042_)
  );
  \$_INV_  _095_ (
    .A(per_addr[0]),
    .Y(_043_)
  );
  \$_AND_  _096_ (
    .A(per_addr[1]),
    .B(_043_),
    .Y(_044_)
  );
  \$_AND_  _097_ (
    .A(_044_),
    .B(_042_),
    .Y(cpu_id_lo_rd[9])
  );
  \$_AND_  _098_ (
    .A(per_addr[1]),
    .B(per_addr[0]),
    .Y(_045_)
  );
  \$_AND_  _099_ (
    .A(_045_),
    .B(_042_),
    .Y(cpu_id_hi_rd[11])
  );
  \$_INV_  _100_ (
    .A(per_din[0]),
    .Y(_046_)
  );
  \$_INV_  _101_ (
    .A(per_addr[1]),
    .Y(_047_)
  );
  \$_AND_  _102_ (
    .A(_047_),
    .B(per_addr[0]),
    .Y(_048_)
  );
  \$_AND_  _103_ (
    .A(_038_),
    .B(per_we[0]),
    .Y(_049_)
  );
  \$_AND_  _104_ (
    .A(_049_),
    .B(_048_),
    .Y(_050_)
  );
  \$_AND_  _105_ (
    .A(_050_),
    .B(_046_),
    .Y(wdtifg_sw_clr)
  );
  \$_AND_  _106_ (
    .A(_050_),
    .B(per_din[0]),
    .Y(wdtifg_sw_set)
  );
  \$_AND_  _107_ (
    .A(ifg1[4]),
    .B(ie1[4]),
    .Y(nmi_pnd)
  );
  \$_AND_  _108_ (
    .A(_047_),
    .B(_043_),
    .Y(_051_)
  );
  \$_AND_  _109_ (
    .A(_051_),
    .B(_042_),
    .Y(_052_)
  );
  \$_AND_  _110_ (
    .A(_052_),
    .B(ie1[4]),
    .Y(_053_)
  );
  \$_AND_  _111_ (
    .A(_048_),
    .B(_042_),
    .Y(_054_)
  );
  \$_AND_  _112_ (
    .A(_054_),
    .B(ifg1[4]),
    .Y(_055_)
  );
  \$_OR_  _113_ (
    .A(_055_),
    .B(_053_),
    .Y(per_dout[4])
  );
  \$_AND_  _114_ (
    .A(_054_),
    .B(wdtifg),
    .Y(_056_)
  );
  \$_AND_  _115_ (
    .A(_052_),
    .B(ie1[0]),
    .Y(_057_)
  );
  \$_OR_  _116_ (
    .A(_057_),
    .B(cpu_id_hi_rd[11]),
    .Y(_058_)
  );
  \$_OR_  _117_ (
    .A(_058_),
    .B(_056_),
    .Y(per_dout[0])
  );
  \$_OR_  _118_ (
    .A(cpu_id_hi_rd[11]),
    .B(cpu_id_lo_rd[9]),
    .Y(per_dout[1])
  );
  \$_INV_  _119_ (
    .A(nmi_acc),
    .Y(_059_)
  );
  \$_INV_  _120_ (
    .A(_016_),
    .Y(_060_)
  );
  \$_OR_  _121_ (
    .A(per_addr[2]),
    .B(per_addr[13]),
    .Y(_061_)
  );
  \$_OR_  _122_ (
    .A(per_addr[4]),
    .B(per_addr[3]),
    .Y(_062_)
  );
  \$_OR_  _123_ (
    .A(_062_),
    .B(_061_),
    .Y(_063_)
  );
  \$_OR_  _124_ (
    .A(_063_),
    .B(_060_),
    .Y(_064_)
  );
  \$_OR_  _125_ (
    .A(per_addr[10]),
    .B(per_addr[9]),
    .Y(_065_)
  );
  \$_OR_  _126_ (
    .A(_065_),
    .B(per_addr[11]),
    .Y(_066_)
  );
  \$_OR_  _127_ (
    .A(per_addr[6]),
    .B(per_addr[5]),
    .Y(_003_)
  );
  \$_OR_  _128_ (
    .A(per_addr[8]),
    .B(per_addr[7]),
    .Y(_004_)
  );
  \$_OR_  _129_ (
    .A(_004_),
    .B(_003_),
    .Y(_005_)
  );
  \$_OR_  _130_ (
    .A(_005_),
    .B(_066_),
    .Y(_006_)
  );
  \$_OR_  _131_ (
    .A(_006_),
    .B(_064_),
    .Y(_007_)
  );
  \$_OR_  _132_ (
    .A(_007_),
    .B(_039_),
    .Y(_008_)
  );
  \$_INV_  _133_ (
    .A(_051_),
    .Y(_009_)
  );
  \$_OR_  _134_ (
    .A(_009_),
    .B(_008_),
    .Y(_010_)
  );
  \$_MUX_  _135_ (
    .A(per_din[4]),
    .B(ie1[4]),
    .S(_010_),
    .Y(_011_)
  );
  \$_AND_  _136_ (
    .A(_011_),
    .B(_059_),
    .Y(_000_)
  );
  \$_MUX_  _137_ (
    .A(per_din[0]),
    .B(ie1[0]),
    .S(_010_),
    .Y(_002_)
  );
  \$_INV_  _138_ (
    .A(nmi_dly),
    .Y(_012_)
  );
  \$_AND_  _139_ (
    .A(_012_),
    .B(nmi_s),
    .Y(_013_)
  );
  \$_MUX_  _140_ (
    .A(ifg1[4]),
    .B(per_din[4]),
    .S(_050_),
    .Y(_014_)
  );
  \$_OR_  _141_ (
    .A(_014_),
    .B(_013_),
    .Y(_001_)
  );
  \$_XOR_  _142_ (
    .A(nmi),
    .B(wdtnmies),
    .Y(nmi_capture)
  );
  \$_DFF_PP0_  \ie1_reg[4]  /* _143_ */ (
    .C(mclk),
    .D(_000_),
    .Q(ie1[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \ie1_reg[0]  /* _144_ */ (
    .C(mclk),
    .D(_002_),
    .Q(ie1[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \ifg1_reg[4]  /* _145_ */ (
    .C(mclk),
    .D(_001_),
    .Q(ifg1[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  nmi_dly_reg /* _146_ */ (
    .C(mclk),
    .D(nmi_s),
    .Q(nmi_dly),
    .R(puc_rst)
  );
  omsp_sync_cell sync_cell_nmi (
    .clk(mclk),
    .data_in(nmi_capture),
    .data_out(nmi_s),
    .rst(puc_rst)
  );
  assign cpu_id = 134414850;
  assign { cpu_id_hi_rd[15:12], cpu_id_hi_rd[10:0] } = { 13'b0000000000000, cpu_id_hi_rd[11], cpu_id_hi_rd[11] };
  assign { cpu_id_lo_rd[15:10], cpu_id_lo_rd[8:0] } = { 13'b0000000000000, cpu_id_lo_rd[9], 1'b0 };
  assign { ie1[7:5], ie1[3:1] } = 6'b000000;
  assign ie1_nxt = per_din[7:0];
  assign { ifg1[7:5], ifg1[3:0] } = { 6'b000000, wdtifg };
  assign ifg1_nxt = per_din[7:0];
  assign nmi_pol = nmi_capture;
  assign nmi_wkup = 1'b0;
  assign nmie = ie1[4];
  assign nmiifg = ifg1[4];
  assign { per_dout[15:5], per_dout[3:2] } = { 4'b0000, cpu_id_hi_rd[11], 1'b0, cpu_id_lo_rd[9], 6'b000000 };
  assign reg_addr = { 1'b0, per_addr[1:0] };
  assign { reg_rd[7:3], reg_rd[1] } = { 1'b0, cpu_id_hi_rd[11], 1'b0, cpu_id_lo_rd[9], 2'b00 };
  assign wdtie = ie1[0];
endmodule

module omsp_sync_cell(data_out, clk, data_in, rst);
  input clk;
  input data_in;
  output data_out;
  wire [1:0] data_sync;
  input rst;
  \$_DFF_PP0_  \data_sync_reg[0]  /* _0_ */ (
    .C(clk),
    .D(data_in),
    .Q(data_sync[0]),
    .R(rst)
  );
  \$_DFF_PP0_  data_out_reg /* _1_ */ (
    .C(clk),
    .D(data_sync[0]),
    .Q(data_out),
    .R(rst)
  );
  assign data_sync[1] = data_out;
endmodule

module omsp_sync_reset(rst_s, clk, rst_a);
  input clk;
  wire [1:0] data_sync;
  input rst_a;
  output rst_s;
  \$_DFF_PP1_  \data_sync_reg[0]  /* _0_ */ (
    .C(clk),
    .D(1'b0),
    .Q(data_sync[0]),
    .R(rst_a)
  );
  \$_DFF_PP1_  \data_sync_reg[1]  /* _1_ */ (
    .C(clk),
    .D(data_sync[0]),
    .Q(data_sync[1]),
    .R(rst_a)
  );
  assign rst_s = data_sync[1];
endmodule

module omsp_watchdog(per_dout, wdt_irq, wdt_reset, wdt_wkup, wdtifg, wdtnmies, aclk, aclk_en, dbg_freeze, mclk, per_addr, per_din, per_en, per_we, por, puc_rst, scan_enable, scan_mode, smclk, smclk_en, wdtie, wdtifg_irq_clr, wdtifg_sw_clr, wdtifg_sw_set);
  wire _000_;
  wire [15:0] _001_;
  wire [7:0] _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  input aclk;
  input aclk_en;
  input dbg_freeze;
  input mclk;
  wire mclk_wdtctl;
  input [13:0] per_addr;
  input [15:0] per_din;
  output [15:0] per_dout;
  input per_en;
  input [1:0] per_we;
  input por;
  input puc_rst;
  wire [1:0] reg_addr;
  wire [3:0] reg_rd;
  input scan_enable;
  input scan_mode;
  input smclk;
  input smclk_en;
  output wdt_irq;
  output wdt_reset;
  output wdt_wkup;
  wire [15:0] wdtcnt;
  wire [7:0] wdtctl;
  wire [15:0] wdtctl_rd;
  input wdtie;
  output wdtifg;
  input wdtifg_irq_clr;
  input wdtifg_sw_clr;
  input wdtifg_sw_set;
  output wdtnmies;
  wire wdttmsel;
  \$_INV_  _124_ (
    .A(per_addr[11]),
    .Y(_121_)
  );
  \$_AND_  _125_ (
    .A(_121_),
    .B(per_en),
    .Y(_122_)
  );
  \$_OR_  _126_ (
    .A(per_addr[13]),
    .B(per_addr[12]),
    .Y(_123_)
  );
  \$_OR_  _127_ (
    .A(per_addr[2]),
    .B(per_addr[1]),
    .Y(_004_)
  );
  \$_OR_  _128_ (
    .A(_004_),
    .B(_123_),
    .Y(_005_)
  );
  \$_INV_  _129_ (
    .A(_005_),
    .Y(_006_)
  );
  \$_AND_  _130_ (
    .A(_006_),
    .B(_122_),
    .Y(_007_)
  );
  \$_OR_  _131_ (
    .A(per_addr[10]),
    .B(per_addr[9]),
    .Y(_008_)
  );
  \$_INV_  _132_ (
    .A(_008_),
    .Y(_009_)
  );
  \$_AND_  _133_ (
    .A(per_addr[7]),
    .B(per_addr[4]),
    .Y(_010_)
  );
  \$_AND_  _134_ (
    .A(_010_),
    .B(_009_),
    .Y(_011_)
  );
  \$_OR_  _135_ (
    .A(per_addr[5]),
    .B(per_addr[3]),
    .Y(_012_)
  );
  \$_OR_  _136_ (
    .A(per_addr[8]),
    .B(per_addr[6]),
    .Y(_013_)
  );
  \$_OR_  _137_ (
    .A(_013_),
    .B(_012_),
    .Y(_014_)
  );
  \$_INV_  _138_ (
    .A(_014_),
    .Y(_015_)
  );
  \$_AND_  _139_ (
    .A(_015_),
    .B(_011_),
    .Y(_016_)
  );
  \$_AND_  _140_ (
    .A(_016_),
    .B(_007_),
    .Y(_017_)
  );
  \$_INV_  _141_ (
    .A(per_addr[0]),
    .Y(_018_)
  );
  \$_OR_  _142_ (
    .A(per_we[1]),
    .B(per_we[0]),
    .Y(_019_)
  );
  \$_INV_  _143_ (
    .A(_019_),
    .Y(_020_)
  );
  \$_AND_  _144_ (
    .A(_020_),
    .B(_018_),
    .Y(_021_)
  );
  \$_AND_  _145_ (
    .A(_021_),
    .B(_017_),
    .Y(per_dout[14])
  );
  \$_AND_  _146_ (
    .A(per_dout[14]),
    .B(wdtctl[0]),
    .Y(per_dout[0])
  );
  \$_AND_  _147_ (
    .A(per_dout[14]),
    .B(wdtctl[1]),
    .Y(per_dout[1])
  );
  \$_AND_  _148_ (
    .A(per_dout[14]),
    .B(wdtctl[2]),
    .Y(per_dout[2])
  );
  \$_AND_  _149_ (
    .A(per_dout[14]),
    .B(wdtctl[3]),
    .Y(per_dout[3])
  );
  \$_AND_  _150_ (
    .A(per_dout[14]),
    .B(wdtctl[4]),
    .Y(per_dout[4])
  );
  \$_AND_  _151_ (
    .A(per_dout[14]),
    .B(wdtctl[6]),
    .Y(per_dout[6])
  );
  \$_AND_  _152_ (
    .A(per_dout[14]),
    .B(wdtctl[7]),
    .Y(per_dout[7])
  );
  \$_AND_  _153_ (
    .A(wdtifg),
    .B(wdtctl[4]),
    .Y(_022_)
  );
  \$_AND_  _154_ (
    .A(_022_),
    .B(wdtie),
    .Y(wdt_irq)
  );
  \$_AND_  _155_ (
    .A(_019_),
    .B(_018_),
    .Y(_023_)
  );
  \$_AND_  _156_ (
    .A(_023_),
    .B(_017_),
    .Y(_024_)
  );
  \$_INV_  _157_ (
    .A(_024_),
    .Y(_025_)
  );
  \$_AND_  _158_ (
    .A(per_din[11]),
    .B(per_din[9]),
    .Y(_026_)
  );
  \$_AND_  _159_ (
    .A(per_din[14]),
    .B(per_din[12]),
    .Y(_027_)
  );
  \$_AND_  _160_ (
    .A(_027_),
    .B(_026_),
    .Y(_028_)
  );
  \$_OR_  _161_ (
    .A(per_din[10]),
    .B(per_din[8]),
    .Y(_029_)
  );
  \$_OR_  _162_ (
    .A(per_din[15]),
    .B(per_din[13]),
    .Y(_030_)
  );
  \$_OR_  _163_ (
    .A(_030_),
    .B(_029_),
    .Y(_031_)
  );
  \$_INV_  _164_ (
    .A(_031_),
    .Y(_032_)
  );
  \$_AND_  _165_ (
    .A(_032_),
    .B(_028_),
    .Y(_033_)
  );
  \$_OR_  _166_ (
    .A(_033_),
    .B(_025_),
    .Y(_034_)
  );
  \$_INV_  _167_ (
    .A(_034_),
    .Y(_035_)
  );
  \$_INV_  _168_ (
    .A(wdtctl[4]),
    .Y(_036_)
  );
  \$_INV_  _169_ (
    .A(wdtctl[0]),
    .Y(_037_)
  );
  \$_INV_  _170_ (
    .A(wdtctl[1]),
    .Y(_038_)
  );
  \$_OR_  _171_ (
    .A(_038_),
    .B(_037_),
    .Y(_039_)
  );
  \$_AND_  _172_ (
    .A(_038_),
    .B(_037_),
    .Y(_040_)
  );
  \$_AND_  _173_ (
    .A(wdtcnt[1]),
    .B(wdtcnt[0]),
    .Y(_041_)
  );
  \$_AND_  _174_ (
    .A(_041_),
    .B(wdtcnt[2]),
    .Y(_042_)
  );
  \$_AND_  _175_ (
    .A(_042_),
    .B(wdtcnt[3]),
    .Y(_043_)
  );
  \$_AND_  _176_ (
    .A(_043_),
    .B(wdtcnt[4]),
    .Y(_044_)
  );
  \$_AND_  _177_ (
    .A(_044_),
    .B(wdtcnt[5]),
    .Y(_045_)
  );
  \$_AND_  _178_ (
    .A(_045_),
    .B(wdtcnt[6]),
    .Y(_046_)
  );
  \$_AND_  _179_ (
    .A(_046_),
    .B(wdtcnt[7]),
    .Y(_047_)
  );
  \$_AND_  _180_ (
    .A(_047_),
    .B(wdtcnt[8]),
    .Y(_048_)
  );
  \$_AND_  _181_ (
    .A(_048_),
    .B(wdtcnt[9]),
    .Y(_049_)
  );
  \$_AND_  _182_ (
    .A(_049_),
    .B(wdtcnt[10]),
    .Y(_050_)
  );
  \$_AND_  _183_ (
    .A(_050_),
    .B(wdtcnt[11]),
    .Y(_051_)
  );
  \$_AND_  _184_ (
    .A(_051_),
    .B(wdtcnt[12]),
    .Y(_052_)
  );
  \$_AND_  _185_ (
    .A(_052_),
    .B(wdtcnt[13]),
    .Y(_053_)
  );
  \$_AND_  _186_ (
    .A(_053_),
    .B(wdtcnt[14]),
    .Y(_054_)
  );
  \$_XOR_  _187_ (
    .A(_054_),
    .B(wdtcnt[15]),
    .Y(_055_)
  );
  \$_AND_  _188_ (
    .A(_055_),
    .B(_040_),
    .Y(_056_)
  );
  \$_AND_  _189_ (
    .A(_038_),
    .B(wdtctl[0]),
    .Y(_057_)
  );
  \$_XOR_  _190_ (
    .A(_052_),
    .B(wdtcnt[13]),
    .Y(_058_)
  );
  \$_AND_  _191_ (
    .A(_058_),
    .B(_057_),
    .Y(_059_)
  );
  \$_AND_  _192_ (
    .A(wdtctl[1]),
    .B(_037_),
    .Y(_060_)
  );
  \$_XOR_  _193_ (
    .A(_048_),
    .B(wdtcnt[9]),
    .Y(_061_)
  );
  \$_AND_  _194_ (
    .A(_061_),
    .B(_060_),
    .Y(_062_)
  );
  \$_OR_  _195_ (
    .A(_062_),
    .B(_059_),
    .Y(_063_)
  );
  \$_OR_  _196_ (
    .A(_063_),
    .B(_056_),
    .Y(_064_)
  );
  \$_XOR_  _197_ (
    .A(_045_),
    .B(wdtcnt[6]),
    .Y(_065_)
  );
  \$_MUX_  _198_ (
    .A(_065_),
    .B(_064_),
    .S(_039_),
    .Y(_066_)
  );
  \$_MUX_  _199_ (
    .A(smclk_en),
    .B(aclk_en),
    .S(wdtctl[2]),
    .Y(_067_)
  );
  \$_OR_  _200_ (
    .A(dbg_freeze),
    .B(wdtctl[7]),
    .Y(_068_)
  );
  \$_INV_  _201_ (
    .A(_068_),
    .Y(_069_)
  );
  \$_AND_  _202_ (
    .A(_069_),
    .B(_067_),
    .Y(_070_)
  );
  \$_AND_  _203_ (
    .A(_070_),
    .B(_066_),
    .Y(_071_)
  );
  \$_OR_  _204_ (
    .A(_071_),
    .B(_035_),
    .Y(_072_)
  );
  \$_OR_  _205_ (
    .A(_072_),
    .B(wdtifg_sw_set),
    .Y(_073_)
  );
  \$_AND_  _206_ (
    .A(_073_),
    .B(_036_),
    .Y(_074_)
  );
  \$_OR_  _207_ (
    .A(_074_),
    .B(_035_),
    .Y(_000_)
  );
  \$_MUX_  _208_ (
    .A(wdtctl[0]),
    .B(per_din[0]),
    .S(_024_),
    .Y(_002_[0])
  );
  \$_MUX_  _209_ (
    .A(wdtctl[1]),
    .B(per_din[1]),
    .S(_024_),
    .Y(_002_[1])
  );
  \$_MUX_  _210_ (
    .A(wdtctl[2]),
    .B(per_din[2]),
    .S(_024_),
    .Y(_002_[2])
  );
  \$_AND_  _211_ (
    .A(_025_),
    .B(wdtctl[3]),
    .Y(_002_[3])
  );
  \$_MUX_  _212_ (
    .A(wdtctl[4]),
    .B(per_din[4]),
    .S(_024_),
    .Y(_002_[4])
  );
  \$_MUX_  _213_ (
    .A(wdtctl[6]),
    .B(per_din[6]),
    .S(_024_),
    .Y(_002_[6])
  );
  \$_MUX_  _214_ (
    .A(wdtctl[7]),
    .B(per_din[7]),
    .S(_024_),
    .Y(_002_[7])
  );
  \$_INV_  _215_ (
    .A(_040_),
    .Y(_075_)
  );
  \$_INV_  _216_ (
    .A(wdtcnt[15]),
    .Y(_076_)
  );
  \$_XOR_  _217_ (
    .A(_054_),
    .B(_076_),
    .Y(_077_)
  );
  \$_OR_  _218_ (
    .A(_077_),
    .B(_075_),
    .Y(_078_)
  );
  \$_INV_  _219_ (
    .A(_063_),
    .Y(_079_)
  );
  \$_AND_  _220_ (
    .A(_079_),
    .B(_078_),
    .Y(_080_)
  );
  \$_INV_  _221_ (
    .A(_065_),
    .Y(_081_)
  );
  \$_MUX_  _222_ (
    .A(_081_),
    .B(_080_),
    .S(_039_),
    .Y(_082_)
  );
  \$_INV_  _223_ (
    .A(_070_),
    .Y(_083_)
  );
  \$_OR_  _224_ (
    .A(_083_),
    .B(_082_),
    .Y(_084_)
  );
  \$_AND_  _225_ (
    .A(_084_),
    .B(_034_),
    .Y(_085_)
  );
  \$_INV_  _226_ (
    .A(per_din[3]),
    .Y(_086_)
  );
  \$_OR_  _227_ (
    .A(_025_),
    .B(_086_),
    .Y(_087_)
  );
  \$_AND_  _228_ (
    .A(_087_),
    .B(_085_),
    .Y(_088_)
  );
  \$_XOR_  _229_ (
    .A(_070_),
    .B(wdtcnt[0]),
    .Y(_089_)
  );
  \$_AND_  _230_ (
    .A(_089_),
    .B(_088_),
    .Y(_001_[0])
  );
  \$_XOR_  _231_ (
    .A(_049_),
    .B(wdtcnt[10]),
    .Y(_090_)
  );
  \$_MUX_  _232_ (
    .A(_090_),
    .B(wdtcnt[10]),
    .S(_083_),
    .Y(_091_)
  );
  \$_AND_  _233_ (
    .A(_091_),
    .B(_088_),
    .Y(_001_[10])
  );
  \$_XOR_  _234_ (
    .A(_050_),
    .B(wdtcnt[11]),
    .Y(_092_)
  );
  \$_MUX_  _235_ (
    .A(_092_),
    .B(wdtcnt[11]),
    .S(_083_),
    .Y(_093_)
  );
  \$_AND_  _236_ (
    .A(_093_),
    .B(_088_),
    .Y(_001_[11])
  );
  \$_XOR_  _237_ (
    .A(_051_),
    .B(wdtcnt[12]),
    .Y(_094_)
  );
  \$_MUX_  _238_ (
    .A(_094_),
    .B(wdtcnt[12]),
    .S(_083_),
    .Y(_095_)
  );
  \$_AND_  _239_ (
    .A(_095_),
    .B(_088_),
    .Y(_001_[12])
  );
  \$_MUX_  _240_ (
    .A(_058_),
    .B(wdtcnt[13]),
    .S(_083_),
    .Y(_096_)
  );
  \$_AND_  _241_ (
    .A(_096_),
    .B(_088_),
    .Y(_001_[13])
  );
  \$_XOR_  _242_ (
    .A(_053_),
    .B(wdtcnt[14]),
    .Y(_097_)
  );
  \$_MUX_  _243_ (
    .A(_097_),
    .B(wdtcnt[14]),
    .S(_083_),
    .Y(_098_)
  );
  \$_AND_  _244_ (
    .A(_098_),
    .B(_088_),
    .Y(_001_[14])
  );
  \$_MUX_  _245_ (
    .A(_055_),
    .B(wdtcnt[15]),
    .S(_083_),
    .Y(_099_)
  );
  \$_AND_  _246_ (
    .A(_099_),
    .B(_088_),
    .Y(_001_[15])
  );
  \$_XOR_  _247_ (
    .A(wdtcnt[1]),
    .B(wdtcnt[0]),
    .Y(_100_)
  );
  \$_MUX_  _248_ (
    .A(wdtcnt[1]),
    .B(_100_),
    .S(_070_),
    .Y(_101_)
  );
  \$_AND_  _249_ (
    .A(_101_),
    .B(_088_),
    .Y(_001_[1])
  );
  \$_XOR_  _250_ (
    .A(_041_),
    .B(wdtcnt[2]),
    .Y(_102_)
  );
  \$_MUX_  _251_ (
    .A(wdtcnt[2]),
    .B(_102_),
    .S(_070_),
    .Y(_103_)
  );
  \$_AND_  _252_ (
    .A(_103_),
    .B(_088_),
    .Y(_001_[2])
  );
  \$_XOR_  _253_ (
    .A(_042_),
    .B(wdtcnt[3]),
    .Y(_104_)
  );
  \$_MUX_  _254_ (
    .A(wdtcnt[3]),
    .B(_104_),
    .S(_070_),
    .Y(_105_)
  );
  \$_AND_  _255_ (
    .A(_105_),
    .B(_088_),
    .Y(_001_[3])
  );
  \$_XOR_  _256_ (
    .A(_043_),
    .B(wdtcnt[4]),
    .Y(_106_)
  );
  \$_MUX_  _257_ (
    .A(_106_),
    .B(wdtcnt[4]),
    .S(_083_),
    .Y(_107_)
  );
  \$_AND_  _258_ (
    .A(_107_),
    .B(_088_),
    .Y(_001_[4])
  );
  \$_XOR_  _259_ (
    .A(_044_),
    .B(wdtcnt[5]),
    .Y(_108_)
  );
  \$_MUX_  _260_ (
    .A(_108_),
    .B(wdtcnt[5]),
    .S(_083_),
    .Y(_109_)
  );
  \$_AND_  _261_ (
    .A(_109_),
    .B(_088_),
    .Y(_001_[5])
  );
  \$_MUX_  _262_ (
    .A(_065_),
    .B(wdtcnt[6]),
    .S(_083_),
    .Y(_110_)
  );
  \$_AND_  _263_ (
    .A(_110_),
    .B(_088_),
    .Y(_001_[6])
  );
  \$_XOR_  _264_ (
    .A(_046_),
    .B(wdtcnt[7]),
    .Y(_111_)
  );
  \$_MUX_  _265_ (
    .A(_111_),
    .B(wdtcnt[7]),
    .S(_083_),
    .Y(_112_)
  );
  \$_AND_  _266_ (
    .A(_112_),
    .B(_088_),
    .Y(_001_[7])
  );
  \$_XOR_  _267_ (
    .A(_047_),
    .B(wdtcnt[8]),
    .Y(_113_)
  );
  \$_MUX_  _268_ (
    .A(_113_),
    .B(wdtcnt[8]),
    .S(_083_),
    .Y(_114_)
  );
  \$_AND_  _269_ (
    .A(_114_),
    .B(_088_),
    .Y(_001_[8])
  );
  \$_MUX_  _270_ (
    .A(_061_),
    .B(wdtcnt[9]),
    .S(_083_),
    .Y(_115_)
  );
  \$_AND_  _271_ (
    .A(_115_),
    .B(_088_),
    .Y(_001_[9])
  );
  \$_INV_  _272_ (
    .A(wdtifg_irq_clr),
    .Y(_116_)
  );
  \$_OR_  _273_ (
    .A(_116_),
    .B(_036_),
    .Y(_117_)
  );
  \$_INV_  _274_ (
    .A(wdtifg_sw_clr),
    .Y(_118_)
  );
  \$_AND_  _275_ (
    .A(_118_),
    .B(wdtifg),
    .Y(_119_)
  );
  \$_AND_  _276_ (
    .A(_119_),
    .B(_117_),
    .Y(_120_)
  );
  \$_OR_  _277_ (
    .A(_120_),
    .B(_073_),
    .Y(_003_)
  );
  \$_DFF_PP0_  \wdtctl_reg[0]  /* _278_ */ (
    .C(mclk),
    .D(_002_[0]),
    .Q(wdtctl[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[1]  /* _279_ */ (
    .C(mclk),
    .D(_002_[1]),
    .Q(wdtctl[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[2]  /* _280_ */ (
    .C(mclk),
    .D(_002_[2]),
    .Q(wdtctl[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[3]  /* _281_ */ (
    .C(mclk),
    .D(_002_[3]),
    .Q(wdtctl[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[4]  /* _282_ */ (
    .C(mclk),
    .D(_002_[4]),
    .Q(wdtctl[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[6]  /* _283_ */ (
    .C(mclk),
    .D(_002_[6]),
    .Q(wdtctl[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtctl_reg[7]  /* _284_ */ (
    .C(mclk),
    .D(_002_[7]),
    .Q(wdtctl[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[0]  /* _285_ */ (
    .C(mclk),
    .D(_001_[0]),
    .Q(wdtcnt[0]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[10]  /* _286_ */ (
    .C(mclk),
    .D(_001_[10]),
    .Q(wdtcnt[10]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[11]  /* _287_ */ (
    .C(mclk),
    .D(_001_[11]),
    .Q(wdtcnt[11]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[12]  /* _288_ */ (
    .C(mclk),
    .D(_001_[12]),
    .Q(wdtcnt[12]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[13]  /* _289_ */ (
    .C(mclk),
    .D(_001_[13]),
    .Q(wdtcnt[13]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[14]  /* _290_ */ (
    .C(mclk),
    .D(_001_[14]),
    .Q(wdtcnt[14]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[15]  /* _291_ */ (
    .C(mclk),
    .D(_001_[15]),
    .Q(wdtcnt[15]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[1]  /* _292_ */ (
    .C(mclk),
    .D(_001_[1]),
    .Q(wdtcnt[1]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[2]  /* _293_ */ (
    .C(mclk),
    .D(_001_[2]),
    .Q(wdtcnt[2]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[3]  /* _294_ */ (
    .C(mclk),
    .D(_001_[3]),
    .Q(wdtcnt[3]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[4]  /* _295_ */ (
    .C(mclk),
    .D(_001_[4]),
    .Q(wdtcnt[4]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[5]  /* _296_ */ (
    .C(mclk),
    .D(_001_[5]),
    .Q(wdtcnt[5]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[6]  /* _297_ */ (
    .C(mclk),
    .D(_001_[6]),
    .Q(wdtcnt[6]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[7]  /* _298_ */ (
    .C(mclk),
    .D(_001_[7]),
    .Q(wdtcnt[7]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[8]  /* _299_ */ (
    .C(mclk),
    .D(_001_[8]),
    .Q(wdtcnt[8]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  \wdtcnt_reg[9]  /* _300_ */ (
    .C(mclk),
    .D(_001_[9]),
    .Q(wdtcnt[9]),
    .R(puc_rst)
  );
  \$_DFF_PP0_  wdtifg_reg /* _301_ */ (
    .C(mclk),
    .D(_003_),
    .Q(wdtifg),
    .R(por)
  );
  \$_DFF_PP0_  wdt_reset_reg /* _302_ */ (
    .C(mclk),
    .D(_000_),
    .Q(wdt_reset),
    .R(por)
  );
  assign mclk_wdtctl = mclk;
  assign { per_dout[15], per_dout[13:8], per_dout[5] } = { 1'b0, per_dout[14], 1'b0, per_dout[14], 2'b00, per_dout[14], per_dout[14] };
  assign reg_addr = { per_addr[0], 1'b0 };
  assign reg_rd = { 3'b000, per_dout[14] };
  assign wdt_wkup = 1'b0;
  assign wdtctl_rd = { 1'b0, per_dout[14], per_dout[14], 1'b0, per_dout[14], 2'b00, per_dout[14], per_dout[7:6], per_dout[14], per_dout[4:0] };
  assign wdtnmies = wdtctl[6];
  assign wdttmsel = wdtctl[4];
endmodule

module openMSP430(aclk, aclk_en, dbg_freeze, dbg_uart_txd, dco_enable, dco_wkup, dmem_addr, dmem_cen, dmem_din, dmem_wen, irq_acc, lfxt_enable, lfxt_wkup, mclk, per_addr, per_din, per_we, per_en, pmem_addr, pmem_cen, pmem_din, pmem_wen, puc_rst, smclk, smclk_en, cpu_en, dbg_en, dbg_uart_rxd, dco_clk, dmem_dout, irq, lfxt_clk, nmi, per_dout, pmem_dout, reset_n, scan_enable, scan_mode, wkup);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  output aclk;
  output aclk_en;
  input cpu_en;
  wire cpu_en_s;
  wire [31:0] cpu_id;
  wire cpuoff;
  wire dbg_clk;
  wire dbg_cpu_reset;
  input dbg_en;
  wire dbg_en_s;
  output dbg_freeze;
  wire dbg_halt_cmd;
  wire dbg_halt_st;
  wire [15:0] dbg_mem_addr;
  wire [15:0] dbg_mem_din;
  wire [15:0] dbg_mem_dout;
  wire dbg_mem_en;
  wire [1:0] dbg_mem_wr;
  wire [15:0] dbg_reg_din;
  wire dbg_reg_wr;
  wire dbg_rst;
  input dbg_uart_rxd;
  output dbg_uart_txd;
  input dco_clk;
  output dco_enable;
  output dco_wkup;
  wire decode_noirq;
  output [5:0] dmem_addr;
  output dmem_cen;
  output [15:0] dmem_din;
  input [15:0] dmem_dout;
  output [1:0] dmem_wen;
  wire [3:0] e_state;
  wire [15:0] eu_mab;
  wire eu_mb_en;
  wire [1:0] eu_mb_wr;
  wire [15:0] eu_mdb_in;
  wire [15:0] eu_mdb_out;
  wire exec_done;
  wire [15:0] fe_mab;
  wire fe_mb_en;
  wire [15:0] fe_mdb_in;
  wire fe_pmem_wait;
  wire gie;
  wire [7:0] inst_ad;
  wire [11:0] inst_alu;
  wire [7:0] inst_as;
  wire inst_bw;
  wire [15:0] inst_dest;
  wire [15:0] inst_dext;
  wire inst_irq_rst;
  wire [7:0] inst_jmp;
  wire inst_mov;
  wire [15:0] inst_sext;
  wire [7:0] inst_so;
  wire [15:0] inst_src;
  wire [2:0] inst_type;
  input [13:0] irq;
  output [13:0] irq_acc;
  input lfxt_clk;
  output lfxt_enable;
  output lfxt_wkup;
  output mclk;
  wire mclk_enable;
  wire mclk_wkup;
  input nmi;
  wire nmi_acc;
  wire nmi_pnd;
  wire nmi_wkup;
  wire oscoff;
  wire [15:0] pc;
  wire [15:0] pc_nxt;
  wire [15:0] pc_sw;
  wire pc_sw_wr;
  output [13:0] per_addr;
  output [15:0] per_din;
  input [15:0] per_dout;
  wire [15:0] per_dout_clk;
  wire [15:0] per_dout_mpy;
  wire [15:0] per_dout_or;
  wire [15:0] per_dout_sfr;
  wire [15:0] per_dout_wdog;
  output per_en;
  output [1:0] per_we;
  output [9:0] pmem_addr;
  output pmem_cen;
  output [15:0] pmem_din;
  input [15:0] pmem_dout;
  output [1:0] pmem_wen;
  wire por;
  wire puc_pnd_set;
  output puc_rst;
  input reset_n;
  input scan_enable;
  input scan_mode;
  wire scg0;
  wire scg1;
  output smclk;
  output smclk_en;
  wire wdt_irq;
  wire wdt_reset;
  wire wdt_wkup;
  wire wdtie;
  wire wdtifg;
  wire wdtifg_sw_clr;
  wire wdtifg_sw_set;
  wire wdtnmies;
  input wkup;
  \$_OR_  _048_ (
    .A(per_dout[0]),
    .B(per_dout_clk[0]),
    .Y(_045_)
  );
  \$_OR_  _049_ (
    .A(per_dout_wdog[0]),
    .B(per_dout_sfr[0]),
    .Y(_046_)
  );
  \$_OR_  _050_ (
    .A(_046_),
    .B(per_dout_mpy[0]),
    .Y(_047_)
  );
  \$_OR_  _051_ (
    .A(_047_),
    .B(_045_),
    .Y(per_dout_or[0])
  );
  \$_OR_  _052_ (
    .A(per_dout[10]),
    .B(per_dout_clk[10]),
    .Y(_000_)
  );
  \$_OR_  _053_ (
    .A(per_dout_wdog[10]),
    .B(per_dout_sfr[10]),
    .Y(_001_)
  );
  \$_OR_  _054_ (
    .A(_001_),
    .B(per_dout_mpy[10]),
    .Y(_002_)
  );
  \$_OR_  _055_ (
    .A(_002_),
    .B(_000_),
    .Y(per_dout_or[10])
  );
  \$_OR_  _056_ (
    .A(per_dout[11]),
    .B(per_dout_clk[11]),
    .Y(_003_)
  );
  \$_OR_  _057_ (
    .A(per_dout_wdog[11]),
    .B(per_dout_sfr[11]),
    .Y(_004_)
  );
  \$_OR_  _058_ (
    .A(_004_),
    .B(per_dout_mpy[11]),
    .Y(_005_)
  );
  \$_OR_  _059_ (
    .A(_005_),
    .B(_003_),
    .Y(per_dout_or[11])
  );
  \$_OR_  _060_ (
    .A(per_dout[12]),
    .B(per_dout_clk[12]),
    .Y(_006_)
  );
  \$_OR_  _061_ (
    .A(per_dout_wdog[12]),
    .B(per_dout_sfr[12]),
    .Y(_007_)
  );
  \$_OR_  _062_ (
    .A(_007_),
    .B(per_dout_mpy[12]),
    .Y(_008_)
  );
  \$_OR_  _063_ (
    .A(_008_),
    .B(_006_),
    .Y(per_dout_or[12])
  );
  \$_OR_  _064_ (
    .A(per_dout[13]),
    .B(per_dout_clk[13]),
    .Y(_009_)
  );
  \$_OR_  _065_ (
    .A(per_dout_wdog[13]),
    .B(per_dout_sfr[13]),
    .Y(_010_)
  );
  \$_OR_  _066_ (
    .A(_010_),
    .B(per_dout_mpy[13]),
    .Y(_011_)
  );
  \$_OR_  _067_ (
    .A(_011_),
    .B(_009_),
    .Y(per_dout_or[13])
  );
  \$_OR_  _068_ (
    .A(per_dout[14]),
    .B(per_dout_clk[14]),
    .Y(_012_)
  );
  \$_OR_  _069_ (
    .A(per_dout_wdog[14]),
    .B(per_dout_sfr[14]),
    .Y(_013_)
  );
  \$_OR_  _070_ (
    .A(_013_),
    .B(per_dout_mpy[14]),
    .Y(_014_)
  );
  \$_OR_  _071_ (
    .A(_014_),
    .B(_012_),
    .Y(per_dout_or[14])
  );
  \$_OR_  _072_ (
    .A(per_dout[15]),
    .B(per_dout_clk[15]),
    .Y(_015_)
  );
  \$_OR_  _073_ (
    .A(per_dout_wdog[15]),
    .B(per_dout_sfr[15]),
    .Y(_016_)
  );
  \$_OR_  _074_ (
    .A(_016_),
    .B(per_dout_mpy[15]),
    .Y(_017_)
  );
  \$_OR_  _075_ (
    .A(_017_),
    .B(_015_),
    .Y(per_dout_or[15])
  );
  \$_OR_  _076_ (
    .A(per_dout[1]),
    .B(per_dout_clk[1]),
    .Y(_018_)
  );
  \$_OR_  _077_ (
    .A(per_dout_wdog[1]),
    .B(per_dout_sfr[1]),
    .Y(_019_)
  );
  \$_OR_  _078_ (
    .A(_019_),
    .B(per_dout_mpy[1]),
    .Y(_020_)
  );
  \$_OR_  _079_ (
    .A(_020_),
    .B(_018_),
    .Y(per_dout_or[1])
  );
  \$_OR_  _080_ (
    .A(per_dout[2]),
    .B(per_dout_clk[2]),
    .Y(_021_)
  );
  \$_OR_  _081_ (
    .A(per_dout_wdog[2]),
    .B(per_dout_sfr[2]),
    .Y(_022_)
  );
  \$_OR_  _082_ (
    .A(_022_),
    .B(per_dout_mpy[2]),
    .Y(_023_)
  );
  \$_OR_  _083_ (
    .A(_023_),
    .B(_021_),
    .Y(per_dout_or[2])
  );
  \$_OR_  _084_ (
    .A(per_dout[3]),
    .B(per_dout_clk[3]),
    .Y(_024_)
  );
  \$_OR_  _085_ (
    .A(per_dout_wdog[3]),
    .B(per_dout_sfr[3]),
    .Y(_025_)
  );
  \$_OR_  _086_ (
    .A(_025_),
    .B(per_dout_mpy[3]),
    .Y(_026_)
  );
  \$_OR_  _087_ (
    .A(_026_),
    .B(_024_),
    .Y(per_dout_or[3])
  );
  \$_OR_  _088_ (
    .A(per_dout[4]),
    .B(per_dout_clk[4]),
    .Y(_027_)
  );
  \$_OR_  _089_ (
    .A(per_dout_wdog[4]),
    .B(per_dout_sfr[4]),
    .Y(_028_)
  );
  \$_OR_  _090_ (
    .A(_028_),
    .B(per_dout_mpy[4]),
    .Y(_029_)
  );
  \$_OR_  _091_ (
    .A(_029_),
    .B(_027_),
    .Y(per_dout_or[4])
  );
  \$_OR_  _092_ (
    .A(per_dout[5]),
    .B(per_dout_clk[5]),
    .Y(_030_)
  );
  \$_OR_  _093_ (
    .A(per_dout_wdog[5]),
    .B(per_dout_sfr[5]),
    .Y(_031_)
  );
  \$_OR_  _094_ (
    .A(_031_),
    .B(per_dout_mpy[5]),
    .Y(_032_)
  );
  \$_OR_  _095_ (
    .A(_032_),
    .B(_030_),
    .Y(per_dout_or[5])
  );
  \$_OR_  _096_ (
    .A(per_dout[6]),
    .B(per_dout_clk[6]),
    .Y(_033_)
  );
  \$_OR_  _097_ (
    .A(per_dout_wdog[6]),
    .B(per_dout_sfr[6]),
    .Y(_034_)
  );
  \$_OR_  _098_ (
    .A(_034_),
    .B(per_dout_mpy[6]),
    .Y(_035_)
  );
  \$_OR_  _099_ (
    .A(_035_),
    .B(_033_),
    .Y(per_dout_or[6])
  );
  \$_OR_  _100_ (
    .A(per_dout[7]),
    .B(per_dout_clk[7]),
    .Y(_036_)
  );
  \$_OR_  _101_ (
    .A(per_dout_wdog[7]),
    .B(per_dout_sfr[7]),
    .Y(_037_)
  );
  \$_OR_  _102_ (
    .A(_037_),
    .B(per_dout_mpy[7]),
    .Y(_038_)
  );
  \$_OR_  _103_ (
    .A(_038_),
    .B(_036_),
    .Y(per_dout_or[7])
  );
  \$_OR_  _104_ (
    .A(per_dout[8]),
    .B(per_dout_clk[8]),
    .Y(_039_)
  );
  \$_OR_  _105_ (
    .A(per_dout_wdog[8]),
    .B(per_dout_sfr[8]),
    .Y(_040_)
  );
  \$_OR_  _106_ (
    .A(_040_),
    .B(per_dout_mpy[8]),
    .Y(_041_)
  );
  \$_OR_  _107_ (
    .A(_041_),
    .B(_039_),
    .Y(per_dout_or[8])
  );
  \$_OR_  _108_ (
    .A(per_dout[9]),
    .B(per_dout_clk[9]),
    .Y(_042_)
  );
  \$_OR_  _109_ (
    .A(per_dout_wdog[9]),
    .B(per_dout_sfr[9]),
    .Y(_043_)
  );
  \$_OR_  _110_ (
    .A(_043_),
    .B(per_dout_mpy[9]),
    .Y(_044_)
  );
  \$_OR_  _111_ (
    .A(_044_),
    .B(_042_),
    .Y(per_dout_or[9])
  );
  omsp_clock_module clock_module_0 (
    .aclk(aclk),
    .aclk_en(aclk_en),
    .cpu_en(cpu_en),
    .cpu_en_s(cpu_en_s),
    .cpuoff(cpuoff),
    .dbg_clk(dbg_clk),
    .dbg_cpu_reset(dbg_cpu_reset),
    .dbg_en(dbg_en),
    .dbg_en_s(dbg_en_s),
    .dbg_rst(dbg_rst),
    .dco_clk(dco_clk),
    .dco_enable(dco_enable),
    .dco_wkup(dco_wkup),
    .lfxt_clk(lfxt_clk),
    .lfxt_enable(lfxt_enable),
    .lfxt_wkup(lfxt_wkup),
    .mclk(mclk),
    .mclk_enable(mclk_enable),
    .mclk_wkup(mclk_wkup),
    .oscoff(oscoff),
    .per_addr(per_addr),
    .per_din(per_din),
    .per_dout(per_dout_clk),
    .per_en(per_en),
    .per_we(per_we),
    .por(por),
    .puc_pnd_set(puc_pnd_set),
    .puc_rst(puc_rst),
    .reset_n(reset_n),
    .scan_enable(scan_enable),
    .scan_mode(scan_mode),
    .scg0(scg0),
    .scg1(scg1),
    .smclk(smclk),
    .smclk_en(smclk_en),
    .wdt_reset(wdt_reset)
  );
  omsp_dbg dbg_0 (
    .cpu_en_s(cpu_en_s),
    .cpu_id(cpu_id),
    .dbg_clk(dbg_clk),
    .dbg_cpu_reset(dbg_cpu_reset),
    .dbg_en_s(dbg_en_s),
    .dbg_freeze(dbg_freeze),
    .dbg_halt_cmd(dbg_halt_cmd),
    .dbg_halt_st(dbg_halt_st),
    .dbg_mem_addr(dbg_mem_addr),
    .dbg_mem_din(dbg_mem_din),
    .dbg_mem_dout(dbg_mem_dout),
    .dbg_mem_en(dbg_mem_en),
    .dbg_mem_wr(dbg_mem_wr),
    .dbg_reg_din(dbg_reg_din),
    .dbg_reg_wr(dbg_reg_wr),
    .dbg_rst(dbg_rst),
    .dbg_uart_rxd(dbg_uart_rxd),
    .dbg_uart_txd(dbg_uart_txd),
    .decode_noirq(decode_noirq),
    .eu_mab(eu_mab),
    .eu_mb_en(eu_mb_en),
    .eu_mb_wr(eu_mb_wr),
    .eu_mdb_in(eu_mdb_in),
    .eu_mdb_out(eu_mdb_out),
    .exec_done(exec_done),
    .fe_mb_en(fe_mb_en),
    .fe_mdb_in(fe_mdb_in),
    .pc(pc),
    .puc_pnd_set(puc_pnd_set)
  );
  omsp_execution_unit execution_unit_0 (
    .cpuoff(cpuoff),
    .dbg_halt_st(dbg_halt_st),
    .dbg_mem_dout(dbg_mem_dout),
    .dbg_reg_din(dbg_reg_din),
    .dbg_reg_wr(dbg_reg_wr),
    .e_state(e_state),
    .exec_done(exec_done),
    .gie(gie),
    .inst_ad(inst_ad),
    .inst_alu(inst_alu),
    .inst_as(inst_as),
    .inst_bw(inst_bw),
    .inst_dest(inst_dest),
    .inst_dext(inst_dext),
    .inst_irq_rst(inst_irq_rst),
    .inst_jmp(inst_jmp),
    .inst_mov(inst_mov),
    .inst_sext(inst_sext),
    .inst_so(inst_so),
    .inst_src(inst_src),
    .inst_type(inst_type),
    .mab(eu_mab),
    .mb_en(eu_mb_en),
    .mb_wr(eu_mb_wr),
    .mclk(mclk),
    .mdb_in(eu_mdb_in),
    .mdb_out(eu_mdb_out),
    .oscoff(oscoff),
    .pc(pc),
    .pc_nxt(pc_nxt),
    .pc_sw(pc_sw),
    .pc_sw_wr(pc_sw_wr),
    .puc_rst(puc_rst),
    .scan_enable(scan_enable),
    .scg0(scg0),
    .scg1(scg1)
  );
  omsp_frontend frontend_0 (
    .cpu_en_s(cpu_en_s),
    .cpuoff(cpuoff),
    .dbg_halt_cmd(dbg_halt_cmd),
    .dbg_halt_st(dbg_halt_st),
    .dbg_reg_sel(dbg_mem_addr[3:0]),
    .decode_noirq(decode_noirq),
    .e_state(e_state),
    .exec_done(exec_done),
    .fe_pmem_wait(fe_pmem_wait),
    .gie(gie),
    .inst_ad(inst_ad),
    .inst_alu(inst_alu),
    .inst_as(inst_as),
    .inst_bw(inst_bw),
    .inst_dest(inst_dest),
    .inst_dext(inst_dext),
    .inst_irq_rst(inst_irq_rst),
    .inst_jmp(inst_jmp),
    .inst_mov(inst_mov),
    .inst_sext(inst_sext),
    .inst_so(inst_so),
    .inst_src(inst_src),
    .inst_type(inst_type),
    .irq(irq),
    .irq_acc(irq_acc),
    .mab(fe_mab),
    .mb_en(fe_mb_en),
    .mclk(mclk),
    .mclk_enable(mclk_enable),
    .mclk_wkup(mclk_wkup),
    .mdb_in(fe_mdb_in),
    .nmi_acc(nmi_acc),
    .nmi_pnd(nmi_pnd),
    .nmi_wkup(nmi_wkup),
    .pc(pc),
    .pc_nxt(pc_nxt),
    .pc_sw(pc_sw),
    .pc_sw_wr(pc_sw_wr),
    .puc_rst(puc_rst),
    .scan_enable(scan_enable),
    .wdt_irq(wdt_irq),
    .wdt_wkup(wdt_wkup),
    .wkup(wkup)
  );
  omsp_mem_backbone mem_backbone_0 (
    .dbg_halt_st(dbg_halt_st),
    .dbg_mem_addr(dbg_mem_addr),
    .dbg_mem_din(dbg_mem_din),
    .dbg_mem_dout(dbg_mem_dout),
    .dbg_mem_en(dbg_mem_en),
    .dbg_mem_wr(dbg_mem_wr),
    .dmem_addr(dmem_addr),
    .dmem_cen(dmem_cen),
    .dmem_din(dmem_din),
    .dmem_dout(dmem_dout),
    .dmem_wen(dmem_wen),
    .eu_mab(eu_mab[15:1]),
    .eu_mb_en(eu_mb_en),
    .eu_mb_wr(eu_mb_wr),
    .eu_mdb_in(eu_mdb_in),
    .eu_mdb_out(eu_mdb_out),
    .fe_mab(fe_mab[15:1]),
    .fe_mb_en(fe_mb_en),
    .fe_mdb_in(fe_mdb_in),
    .fe_pmem_wait(fe_pmem_wait),
    .mclk(mclk),
    .per_addr(per_addr),
    .per_din(per_din),
    .per_dout(per_dout_or),
    .per_en(per_en),
    .per_we(per_we),
    .pmem_addr(pmem_addr),
    .pmem_cen(pmem_cen),
    .pmem_din(pmem_din),
    .pmem_dout(pmem_dout),
    .pmem_wen(pmem_wen),
    .puc_rst(puc_rst),
    .scan_enable(scan_enable)
  );
  omsp_multiplier multiplier_0 (
    .mclk(mclk),
    .per_addr(per_addr),
    .per_din(per_din),
    .per_dout(per_dout_mpy),
    .per_en(per_en),
    .per_we(per_we),
    .puc_rst(puc_rst),
    .scan_enable(scan_enable)
  );
  omsp_sfr sfr_0 (
    .cpu_id(cpu_id),
    .mclk(mclk),
    .nmi(nmi),
    .nmi_acc(nmi_acc),
    .nmi_pnd(nmi_pnd),
    .nmi_wkup(nmi_wkup),
    .per_addr(per_addr),
    .per_din(per_din),
    .per_dout(per_dout_sfr),
    .per_en(per_en),
    .per_we(per_we),
    .puc_rst(puc_rst),
    .scan_mode(scan_mode),
    .wdtie(wdtie),
    .wdtifg(wdtifg),
    .wdtifg_sw_clr(wdtifg_sw_clr),
    .wdtifg_sw_set(wdtifg_sw_set),
    .wdtnmies(wdtnmies)
  );
  omsp_watchdog watchdog_0 (
    .aclk(aclk),
    .aclk_en(aclk_en),
    .dbg_freeze(dbg_freeze),
    .mclk(mclk),
    .per_addr(per_addr),
    .per_din(per_din),
    .per_dout(per_dout_wdog),
    .per_en(per_en),
    .per_we(per_we),
    .por(por),
    .puc_rst(puc_rst),
    .scan_enable(scan_enable),
    .scan_mode(scan_mode),
    .smclk(smclk),
    .smclk_en(smclk_en),
    .wdt_irq(wdt_irq),
    .wdt_reset(wdt_reset),
    .wdt_wkup(wdt_wkup),
    .wdtie(wdtie),
    .wdtifg(wdtifg),
    .wdtifg_irq_clr(irq_acc[10]),
    .wdtifg_sw_clr(wdtifg_sw_clr),
    .wdtifg_sw_set(wdtifg_sw_set),
    .wdtnmies(wdtnmies)
  );
endmodule
