/*
:name: string_len
:description: string.len()  tests
:tags: 6.16.1
*/
module top();
	string a = "Test";
	int b = a.len();
endmodule
