/*
:name: class_test_29
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo extends Base implements Pkg::Bar, Baz; endclass