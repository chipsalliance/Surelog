/*
:name: class_test_34
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class zzyyy;
extern function void set_port(dbg_pkg::analysis_port #(1,N) apb);
endclass