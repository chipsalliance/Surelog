/*
:name: class_member_test_23
:description: Test
:tags: 8.3
*/
class myclass;
extern function void subr(mypkg::foo y[M]);
endclass