///////////////////////////////////////////////////////
//     Copyright (c) 2011 Xilinx Inc.
// 
//    Licensed under the Apache License, Version 2.0 (the "License");
//    you may not use this file except in compliance with the License.
//    You may obtain a copy of the License at
// 
//        http://www.apache.org/licenses/LICENSE-2.0
// 
//    Unless required by applicable law or agreed to in writing, software
//    distributed under the License is distributed on an "AS IS" BASIS,
//    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//    See the License for the specific language governing permissions and
//    limitations under the License.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     :  13.1
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : PCIE_2_1.uniprim.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Generated by :	/home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
//  Revision:		1.0
//  01/18/13 - 695630 - added drp monitor
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module PCIE_2_1 (
  CFGAERECRCCHECKEN,
  CFGAERECRCGENEN,
  CFGAERROOTERRCORRERRRECEIVED,
  CFGAERROOTERRCORRERRREPORTINGEN,
  CFGAERROOTERRFATALERRRECEIVED,
  CFGAERROOTERRFATALERRREPORTINGEN,
  CFGAERROOTERRNONFATALERRRECEIVED,
  CFGAERROOTERRNONFATALERRREPORTINGEN,
  CFGBRIDGESERREN,
  CFGCOMMANDBUSMASTERENABLE,
  CFGCOMMANDINTERRUPTDISABLE,
  CFGCOMMANDIOENABLE,
  CFGCOMMANDMEMENABLE,
  CFGCOMMANDSERREN,
  CFGDEVCONTROL2ARIFORWARDEN,
  CFGDEVCONTROL2ATOMICEGRESSBLOCK,
  CFGDEVCONTROL2ATOMICREQUESTEREN,
  CFGDEVCONTROL2CPLTIMEOUTDIS,
  CFGDEVCONTROL2CPLTIMEOUTVAL,
  CFGDEVCONTROL2IDOCPLEN,
  CFGDEVCONTROL2IDOREQEN,
  CFGDEVCONTROL2LTREN,
  CFGDEVCONTROL2TLPPREFIXBLOCK,
  CFGDEVCONTROLAUXPOWEREN,
  CFGDEVCONTROLCORRERRREPORTINGEN,
  CFGDEVCONTROLENABLERO,
  CFGDEVCONTROLEXTTAGEN,
  CFGDEVCONTROLFATALERRREPORTINGEN,
  CFGDEVCONTROLMAXPAYLOAD,
  CFGDEVCONTROLMAXREADREQ,
  CFGDEVCONTROLNONFATALREPORTINGEN,
  CFGDEVCONTROLNOSNOOPEN,
  CFGDEVCONTROLPHANTOMEN,
  CFGDEVCONTROLURERRREPORTINGEN,
  CFGDEVSTATUSCORRERRDETECTED,
  CFGDEVSTATUSFATALERRDETECTED,
  CFGDEVSTATUSNONFATALERRDETECTED,
  CFGDEVSTATUSURDETECTED,
  CFGERRAERHEADERLOGSETN,
  CFGERRCPLRDYN,
  CFGINTERRUPTDO,
  CFGINTERRUPTMMENABLE,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFM,
  CFGINTERRUPTRDYN,
  CFGLINKCONTROLASPMCONTROL,
  CFGLINKCONTROLAUTOBANDWIDTHINTEN,
  CFGLINKCONTROLBANDWIDTHINTEN,
  CFGLINKCONTROLCLOCKPMEN,
  CFGLINKCONTROLCOMMONCLOCK,
  CFGLINKCONTROLEXTENDEDSYNC,
  CFGLINKCONTROLHWAUTOWIDTHDIS,
  CFGLINKCONTROLLINKDISABLE,
  CFGLINKCONTROLRCB,
  CFGLINKCONTROLRETRAINLINK,
  CFGLINKSTATUSAUTOBANDWIDTHSTATUS,
  CFGLINKSTATUSBANDWIDTHSTATUS,
  CFGLINKSTATUSCURRENTSPEED,
  CFGLINKSTATUSDLLACTIVE,
  CFGLINKSTATUSLINKTRAINING,
  CFGLINKSTATUSNEGOTIATEDWIDTH,
  CFGMGMTDO,
  CFGMGMTRDWRDONEN,
  CFGMSGDATA,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDASSERTINTA,
  CFGMSGRECEIVEDASSERTINTB,
  CFGMSGRECEIVEDASSERTINTC,
  CFGMSGRECEIVEDASSERTINTD,
  CFGMSGRECEIVEDDEASSERTINTA,
  CFGMSGRECEIVEDDEASSERTINTB,
  CFGMSGRECEIVEDDEASSERTINTC,
  CFGMSGRECEIVEDDEASSERTINTD,
  CFGMSGRECEIVEDERRCOR,
  CFGMSGRECEIVEDERRFATAL,
  CFGMSGRECEIVEDERRNONFATAL,
  CFGMSGRECEIVEDPMASNAK,
  CFGMSGRECEIVEDPMETO,
  CFGMSGRECEIVEDPMETOACK,
  CFGMSGRECEIVEDPMPME,
  CFGMSGRECEIVEDSETSLOTPOWERLIMIT,
  CFGMSGRECEIVEDUNLOCK,
  CFGPCIELINKSTATE,
  CFGPMCSRPMEEN,
  CFGPMCSRPMESTATUS,
  CFGPMCSRPOWERSTATE,
  CFGPMRCVASREQL1N,
  CFGPMRCVENTERL1N,
  CFGPMRCVENTERL23N,
  CFGPMRCVREQACKN,
  CFGROOTCONTROLPMEINTEN,
  CFGROOTCONTROLSYSERRCORRERREN,
  CFGROOTCONTROLSYSERRFATALERREN,
  CFGROOTCONTROLSYSERRNONFATALERREN,
  CFGSLOTCONTROLELECTROMECHILCTLPULSE,
  CFGTRANSACTION,
  CFGTRANSACTIONADDR,
  CFGTRANSACTIONTYPE,
  CFGVCTCVCMAP,
  DBGSCLRA,
  DBGSCLRB,
  DBGSCLRC,
  DBGSCLRD,
  DBGSCLRE,
  DBGSCLRF,
  DBGSCLRG,
  DBGSCLRH,
  DBGSCLRI,
  DBGSCLRJ,
  DBGSCLRK,
  DBGVECA,
  DBGVECB,
  DBGVECC,
  DRPDO,
  DRPRDY,
  LL2BADDLLPERR,
  LL2BADTLPERR,
  LL2LINKSTATUS,
  LL2PROTOCOLERR,
  LL2RECEIVERERR,
  LL2REPLAYROERR,
  LL2REPLAYTOERR,
  LL2SUSPENDOK,
  LL2TFCINIT1SEQ,
  LL2TFCINIT2SEQ,
  LL2TXIDLE,
  LNKCLKEN,
  MIMRXRADDR,
  MIMRXREN,
  MIMRXWADDR,
  MIMRXWDATA,
  MIMRXWEN,
  MIMTXRADDR,
  MIMTXREN,
  MIMTXWADDR,
  MIMTXWDATA,
  MIMTXWEN,
  PIPERX0POLARITY,
  PIPERX1POLARITY,
  PIPERX2POLARITY,
  PIPERX3POLARITY,
  PIPERX4POLARITY,
  PIPERX5POLARITY,
  PIPERX6POLARITY,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0ELECIDLE,
  PIPETX0POWERDOWN,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1ELECIDLE,
  PIPETX1POWERDOWN,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2ELECIDLE,
  PIPETX2POWERDOWN,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3ELECIDLE,
  PIPETX3POWERDOWN,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4ELECIDLE,
  PIPETX4POWERDOWN,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5ELECIDLE,
  PIPETX5POWERDOWN,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6ELECIDLE,
  PIPETX6POWERDOWN,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7ELECIDLE,
  PIPETX7POWERDOWN,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PL2L0REQ,
  PL2LINKUP,
  PL2RECEIVERERR,
  PL2RECOVERY,
  PL2RXELECIDLE,
  PL2RXPMSTATE,
  PL2SUSPENDOK,
  PLDBGVEC,
  PLDIRECTEDCHANGEDONE,
  PLINITIALLINKWIDTH,
  PLLANEREVERSALMODE,
  PLLINKGEN2CAP,
  PLLINKPARTNERGEN2SUPPORTED,
  PLLINKUPCFGCAP,
  PLLTSSMSTATE,
  PLPHYLNKUPN,
  PLRECEIVEDHOTRST,
  PLRXPMSTATE,
  PLSELLNKRATE,
  PLSELLNKWIDTH,
  PLTXPMSTATE,
  RECEIVEDFUNCLVLRSTN,
  TL2ASPMSUSPENDCREDITCHECKOK,
  TL2ASPMSUSPENDREQ,
  TL2ERRFCPE,
  TL2ERRHDR,
  TL2ERRMALFORMED,
  TL2ERRRXOVERFLOW,
  TL2PPMSUSPENDOK,
  TRNFCCPLD,
  TRNFCCPLH,
  TRNFCNPD,
  TRNFCNPH,
  TRNFCPD,
  TRNFCPH,
  TRNLNKUP,
  TRNRBARHIT,
  TRNRD,
  TRNRDLLPDATA,
  TRNRDLLPSRCRDY,
  TRNRECRCERR,
  TRNREOF,
  TRNRERRFWD,
  TRNRREM,
  TRNRSOF,
  TRNRSRCDSC,
  TRNRSRCRDY,
  TRNTBUFAV,
  TRNTCFGREQ,
  TRNTDLLPDSTRDY,
  TRNTDSTRDY,
  TRNTERRDROP,
  USERRSTN,

  CFGAERINTERRUPTMSGNUM,
  CFGDEVID,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGERRACSN,
  CFGERRAERHEADERLOG,
  CFGERRATOMICEGRESSBLOCKEDN,
  CFGERRCORN,
  CFGERRCPLABORTN,
  CFGERRCPLTIMEOUTN,
  CFGERRCPLUNEXPECTN,
  CFGERRECRCN,
  CFGERRINTERNALCORN,
  CFGERRINTERNALUNCORN,
  CFGERRLOCKEDN,
  CFGERRMALFORMEDN,
  CFGERRMCBLOCKEDN,
  CFGERRNORECOVERYN,
  CFGERRPOISONEDN,
  CFGERRPOSTEDN,
  CFGERRTLPCPLHEADER,
  CFGERRURN,
  CFGFORCECOMMONCLOCKOFF,
  CFGFORCEEXTENDEDSYNCON,
  CFGFORCEMPS,
  CFGINTERRUPTASSERTN,
  CFGINTERRUPTDI,
  CFGINTERRUPTN,
  CFGINTERRUPTSTATN,
  CFGMGMTBYTEENN,
  CFGMGMTDI,
  CFGMGMTDWADDR,
  CFGMGMTRDENN,
  CFGMGMTWRENN,
  CFGMGMTWRREADONLYN,
  CFGMGMTWRRW1CASRWN,
  CFGPCIECAPINTERRUPTMSGNUM,
  CFGPMFORCESTATE,
  CFGPMFORCESTATEENN,
  CFGPMHALTASPML0SN,
  CFGPMHALTASPML1N,
  CFGPMSENDPMETON,
  CFGPMTURNOFFOKN,
  CFGPMWAKEN,
  CFGPORTNUMBER,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENDID,
  CFGTRNPENDINGN,
  CFGVENDID,
  CMRSTN,
  CMSTICKYRSTN,
  DBGMODE,
  DBGSUBMODE,
  DLRSTN,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  FUNCLVLRSTN,
  LL2SENDASREQL1,
  LL2SENDENTERL1,
  LL2SENDENTERL23,
  LL2SENDPMACK,
  LL2SUSPENDNOW,
  LL2TLPRCV,
  MIMRXRDATA,
  MIMTXRDATA,
  PIPECLK,
  PIPERX0CHANISALIGNED,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0ELECIDLE,
  PIPERX0PHYSTATUS,
  PIPERX0STATUS,
  PIPERX0VALID,
  PIPERX1CHANISALIGNED,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1ELECIDLE,
  PIPERX1PHYSTATUS,
  PIPERX1STATUS,
  PIPERX1VALID,
  PIPERX2CHANISALIGNED,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2ELECIDLE,
  PIPERX2PHYSTATUS,
  PIPERX2STATUS,
  PIPERX2VALID,
  PIPERX3CHANISALIGNED,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3ELECIDLE,
  PIPERX3PHYSTATUS,
  PIPERX3STATUS,
  PIPERX3VALID,
  PIPERX4CHANISALIGNED,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4ELECIDLE,
  PIPERX4PHYSTATUS,
  PIPERX4STATUS,
  PIPERX4VALID,
  PIPERX5CHANISALIGNED,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5ELECIDLE,
  PIPERX5PHYSTATUS,
  PIPERX5STATUS,
  PIPERX5VALID,
  PIPERX6CHANISALIGNED,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6ELECIDLE,
  PIPERX6PHYSTATUS,
  PIPERX6STATUS,
  PIPERX6VALID,
  PIPERX7CHANISALIGNED,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7ELECIDLE,
  PIPERX7PHYSTATUS,
  PIPERX7STATUS,
  PIPERX7VALID,
  PL2DIRECTEDLSTATE,
  PLDBGMODE,
  PLDIRECTEDLINKAUTON,
  PLDIRECTEDLINKCHANGE,
  PLDIRECTEDLINKSPEED,
  PLDIRECTEDLINKWIDTH,
  PLDIRECTEDLTSSMNEW,
  PLDIRECTEDLTSSMNEWVLD,
  PLDIRECTEDLTSSMSTALL,
  PLDOWNSTREAMDEEMPHSOURCE,
  PLRSTN,
  PLTRANSMITHOTRST,
  PLUPSTREAMPREFERDEEMPH,
  SYSRSTN,
  TL2ASPMSUSPENDCREDITCHECK,
  TL2PPMSUSPENDREQ,
  TLRSTN,
  TRNFCSEL,
  TRNRDSTRDY,
  TRNRFCPRET,
  TRNRNPOK,
  TRNRNPREQ,
  TRNTCFGGNT,
  TRNTD,
  TRNTDLLPDATA,
  TRNTDLLPSRCRDY,
  TRNTECRCGEN,
  TRNTEOF,
  TRNTERRFWD,
  TRNTREM,
  TRNTSOF,
  TRNTSRCDSC,
  TRNTSRCRDY,
  TRNTSTR,
  USERCLK,
  USERCLK2
);

  `ifdef XIL_TIMING //Simprim 
  parameter LOC = "UNPLACED";
  `endif
  parameter [11:0] AER_BASE_PTR = 12'h140;
  parameter AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
  parameter AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
  parameter [15:0] AER_CAP_ID = 16'h0001;
  parameter AER_CAP_MULTIHEADER = "FALSE";
  parameter [11:0] AER_CAP_NEXTPTR = 12'h178;
  parameter AER_CAP_ON = "FALSE";
  parameter [23:0] AER_CAP_OPTIONAL_ERR_SUPPORT = 24'h000000;
  parameter AER_CAP_PERMIT_ROOTERR_UPDATE = "TRUE";
  parameter [3:0] AER_CAP_VERSION = 4'h2;
  parameter ALLOW_X8_GEN2 = "FALSE";
  parameter [31:0] BAR0 = 32'hFFFFFF00;
  parameter [31:0] BAR1 = 32'hFFFF0000;
  parameter [31:0] BAR2 = 32'hFFFF000C;
  parameter [31:0] BAR3 = 32'hFFFFFFFF;
  parameter [31:0] BAR4 = 32'h00000000;
  parameter [31:0] BAR5 = 32'h00000000;
  parameter [7:0] CAPABILITIES_PTR = 8'h40;
  parameter [31:0] CARDBUS_CIS_POINTER = 32'h00000000;
  parameter integer CFG_ECRC_ERR_CPLSTAT = 0;
  parameter [23:0] CLASS_CODE = 24'h000000;
  parameter CMD_INTX_IMPLEMENTED = "TRUE";
  parameter CPL_TIMEOUT_DISABLE_SUPPORTED = "FALSE";
  parameter [3:0] CPL_TIMEOUT_RANGES_SUPPORTED = 4'h0;
  parameter [6:0] CRM_MODULE_RSTS = 7'h00;
  parameter DEV_CAP2_ARI_FORWARDING_SUPPORTED = "FALSE";
  parameter DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED = "FALSE";
  parameter DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED = "FALSE";
  parameter DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED = "FALSE";
  parameter DEV_CAP2_CAS128_COMPLETER_SUPPORTED = "FALSE";
  parameter DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED = "FALSE";
  parameter DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED = "FALSE";
  parameter DEV_CAP2_LTR_MECHANISM_SUPPORTED = "FALSE";
  parameter [1:0] DEV_CAP2_MAX_ENDEND_TLP_PREFIXES = 2'h0;
  parameter DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING = "FALSE";
  parameter [1:0] DEV_CAP2_TPH_COMPLETER_SUPPORTED = 2'h0;
  parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE = "TRUE";
  parameter DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE = "TRUE";
  parameter integer DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
  parameter integer DEV_CAP_ENDPOINT_L1_LATENCY = 0;
  parameter DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
  parameter DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "FALSE";
  parameter integer DEV_CAP_MAX_PAYLOAD_SUPPORTED = 2;
  parameter integer DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT = 0;
  parameter DEV_CAP_ROLE_BASED_ERROR = "TRUE";
  parameter integer DEV_CAP_RSVD_14_12 = 0;
  parameter integer DEV_CAP_RSVD_17_16 = 0;
  parameter integer DEV_CAP_RSVD_31_29 = 0;
  parameter DEV_CONTROL_AUX_POWER_SUPPORTED = "FALSE";
  parameter DEV_CONTROL_EXT_TAG_DEFAULT = "FALSE";
  parameter DISABLE_ASPM_L1_TIMER = "FALSE";
  parameter DISABLE_BAR_FILTERING = "FALSE";
  parameter DISABLE_ERR_MSG = "FALSE";
  parameter DISABLE_ID_CHECK = "FALSE";
  parameter DISABLE_LANE_REVERSAL = "FALSE";
  parameter DISABLE_LOCKED_FILTER = "FALSE";
  parameter DISABLE_PPM_FILTER = "FALSE";
  parameter DISABLE_RX_POISONED_RESP = "FALSE";
  parameter DISABLE_RX_TC_FILTER = "FALSE";
  parameter DISABLE_SCRAMBLING = "FALSE";
  parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
  parameter [11:0] DSN_BASE_PTR = 12'h100;
  parameter [15:0] DSN_CAP_ID = 16'h0003;
  parameter [11:0] DSN_CAP_NEXTPTR = 12'h10C;
  parameter DSN_CAP_ON = "TRUE";
  parameter [3:0] DSN_CAP_VERSION = 4'h1;
  parameter [10:0] ENABLE_MSG_ROUTE = 11'h000;
  parameter ENABLE_RX_TD_ECRC_TRIM = "FALSE";
  parameter ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED = "FALSE";
  parameter ENTER_RVRY_EI_L0 = "TRUE";
  parameter EXIT_LOOPBACK_ON_EI = "TRUE";
  parameter [31:0] EXPANSION_ROM = 32'hFFFFF001;
  parameter [5:0] EXT_CFG_CAP_PTR = 6'h3F;
  parameter [9:0] EXT_CFG_XP_CAP_PTR = 10'h3FF;
  parameter [7:0] HEADER_TYPE = 8'h00;
  parameter [4:0] INFER_EI = 5'h00;
  parameter [7:0] INTERRUPT_PIN = 8'h01;
  parameter INTERRUPT_STAT_AUTO = "TRUE";
  parameter IS_SWITCH = "FALSE";
  parameter [9:0] LAST_CONFIG_DWORD = 10'h3FF;
  parameter LINK_CAP_ASPM_OPTIONALITY = "TRUE";
  parameter integer LINK_CAP_ASPM_SUPPORT = 1;
  parameter LINK_CAP_CLOCK_POWER_MANAGEMENT = "FALSE";
  parameter LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP = "FALSE";
  parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
  parameter integer LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
  parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
  parameter integer LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
  parameter LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP = "FALSE";
  parameter [3:0] LINK_CAP_MAX_LINK_SPEED = 4'h1;
  parameter [5:0] LINK_CAP_MAX_LINK_WIDTH = 6'h08;
  parameter integer LINK_CAP_RSVD_23 = 0;
  parameter LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE = "FALSE";
  parameter integer LINK_CONTROL_RCB = 0;
  parameter LINK_CTRL2_DEEMPHASIS = "FALSE";
  parameter LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE = "FALSE";
  parameter [3:0] LINK_CTRL2_TARGET_LINK_SPEED = 4'h2;
  parameter LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
  parameter [14:0] LL_ACK_TIMEOUT = 15'h0000;
  parameter LL_ACK_TIMEOUT_EN = "FALSE";
  parameter integer LL_ACK_TIMEOUT_FUNC = 0;
  parameter [14:0] LL_REPLAY_TIMEOUT = 15'h0000;
  parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
  parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
  parameter [5:0] LTSSM_MAX_LINK_WIDTH = 6'h01;
  parameter MPS_FORCE = "FALSE";
  parameter [7:0] MSIX_BASE_PTR = 8'h9C;
  parameter [7:0] MSIX_CAP_ID = 8'h11;
  parameter [7:0] MSIX_CAP_NEXTPTR = 8'h00;
  parameter MSIX_CAP_ON = "FALSE";
  parameter integer MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter [7:0] MSI_BASE_PTR = 8'h48;
  parameter MSI_CAP_64_BIT_ADDR_CAPABLE = "TRUE";
  parameter [7:0] MSI_CAP_ID = 8'h05;
  parameter integer MSI_CAP_MULTIMSGCAP = 0;
  parameter integer MSI_CAP_MULTIMSG_EXTENSION = 0;
  parameter [7:0] MSI_CAP_NEXTPTR = 8'h60;
  parameter MSI_CAP_ON = "FALSE";
  parameter MSI_CAP_PER_VECTOR_MASKING_CAPABLE = "TRUE";
  parameter integer N_FTS_COMCLK_GEN1 = 255;
  parameter integer N_FTS_COMCLK_GEN2 = 255;
  parameter integer N_FTS_GEN1 = 255;
  parameter integer N_FTS_GEN2 = 255;
  parameter [7:0] PCIE_BASE_PTR = 8'h60;
  parameter [7:0] PCIE_CAP_CAPABILITY_ID = 8'h10;
  parameter [3:0] PCIE_CAP_CAPABILITY_VERSION = 4'h2;
  parameter [3:0] PCIE_CAP_DEVICE_PORT_TYPE = 4'h0;
  parameter [7:0] PCIE_CAP_NEXTPTR = 8'h9C;
  parameter PCIE_CAP_ON = "TRUE";
  parameter integer PCIE_CAP_RSVD_15_14 = 0;
  parameter PCIE_CAP_SLOT_IMPLEMENTED = "FALSE";
  parameter integer PCIE_REVISION = 2;
  parameter integer PL_AUTO_CONFIG = 0;
  parameter PL_FAST_TRAIN = "FALSE";
  parameter [14:0] PM_ASPML0S_TIMEOUT = 15'h0000;
  parameter PM_ASPML0S_TIMEOUT_EN = "FALSE";
  parameter integer PM_ASPML0S_TIMEOUT_FUNC = 0;
  parameter PM_ASPM_FASTEXIT = "FALSE";
  parameter [7:0] PM_BASE_PTR = 8'h40;
  parameter integer PM_CAP_AUXCURRENT = 0;
  parameter PM_CAP_D1SUPPORT = "TRUE";
  parameter PM_CAP_D2SUPPORT = "TRUE";
  parameter PM_CAP_DSI = "FALSE";
  parameter [7:0] PM_CAP_ID = 8'h01;
  parameter [7:0] PM_CAP_NEXTPTR = 8'h48;
  parameter PM_CAP_ON = "TRUE";
  parameter [4:0] PM_CAP_PMESUPPORT = 5'h0F;
  parameter PM_CAP_PME_CLOCK = "FALSE";
  parameter integer PM_CAP_RSVD_04 = 0;
  parameter integer PM_CAP_VERSION = 3;
  parameter PM_CSR_B2B3 = "FALSE";
  parameter PM_CSR_BPCCEN = "FALSE";
  parameter PM_CSR_NOSOFTRST = "TRUE";
  parameter [7:0] PM_DATA0 = 8'h01;
  parameter [7:0] PM_DATA1 = 8'h01;
  parameter [7:0] PM_DATA2 = 8'h01;
  parameter [7:0] PM_DATA3 = 8'h01;
  parameter [7:0] PM_DATA4 = 8'h01;
  parameter [7:0] PM_DATA5 = 8'h01;
  parameter [7:0] PM_DATA6 = 8'h01;
  parameter [7:0] PM_DATA7 = 8'h01;
  parameter [1:0] PM_DATA_SCALE0 = 2'h1;
  parameter [1:0] PM_DATA_SCALE1 = 2'h1;
  parameter [1:0] PM_DATA_SCALE2 = 2'h1;
  parameter [1:0] PM_DATA_SCALE3 = 2'h1;
  parameter [1:0] PM_DATA_SCALE4 = 2'h1;
  parameter [1:0] PM_DATA_SCALE5 = 2'h1;
  parameter [1:0] PM_DATA_SCALE6 = 2'h1;
  parameter [1:0] PM_DATA_SCALE7 = 2'h1;
  parameter PM_MF = "FALSE";
  parameter [11:0] RBAR_BASE_PTR = 12'h178;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR0 = 5'h00;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR1 = 5'h00;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR2 = 5'h00;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR3 = 5'h00;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR4 = 5'h00;
  parameter [4:0] RBAR_CAP_CONTROL_ENCODEDBAR5 = 5'h00;
  parameter [15:0] RBAR_CAP_ID = 16'h0015;
  parameter [2:0] RBAR_CAP_INDEX0 = 3'h0;
  parameter [2:0] RBAR_CAP_INDEX1 = 3'h0;
  parameter [2:0] RBAR_CAP_INDEX2 = 3'h0;
  parameter [2:0] RBAR_CAP_INDEX3 = 3'h0;
  parameter [2:0] RBAR_CAP_INDEX4 = 3'h0;
  parameter [2:0] RBAR_CAP_INDEX5 = 3'h0;
  parameter [11:0] RBAR_CAP_NEXTPTR = 12'h000;
  parameter RBAR_CAP_ON = "FALSE";
  parameter [31:0] RBAR_CAP_SUP0 = 32'h00000000;
  parameter [31:0] RBAR_CAP_SUP1 = 32'h00000000;
  parameter [31:0] RBAR_CAP_SUP2 = 32'h00000000;
  parameter [31:0] RBAR_CAP_SUP3 = 32'h00000000;
  parameter [31:0] RBAR_CAP_SUP4 = 32'h00000000;
  parameter [31:0] RBAR_CAP_SUP5 = 32'h00000000;
  parameter [3:0] RBAR_CAP_VERSION = 4'h1;
  parameter [2:0] RBAR_NUM = 3'h1;
  parameter integer RECRC_CHK = 0;
  parameter RECRC_CHK_TRIM = "FALSE";
  parameter ROOT_CAP_CRS_SW_VISIBILITY = "FALSE";
  parameter [1:0] RP_AUTO_SPD = 2'h1;
  parameter [4:0] RP_AUTO_SPD_LOOPCNT = 5'h1F;
  parameter SELECT_DLL_IF = "FALSE";
  parameter SIM_VERSION = "1.0";
  parameter SLOT_CAP_ATT_BUTTON_PRESENT = "FALSE";
  parameter SLOT_CAP_ATT_INDICATOR_PRESENT = "FALSE";
  parameter SLOT_CAP_ELEC_INTERLOCK_PRESENT = "FALSE";
  parameter SLOT_CAP_HOTPLUG_CAPABLE = "FALSE";
  parameter SLOT_CAP_HOTPLUG_SURPRISE = "FALSE";
  parameter SLOT_CAP_MRL_SENSOR_PRESENT = "FALSE";
  parameter SLOT_CAP_NO_CMD_COMPLETED_SUPPORT = "FALSE";
  parameter [12:0] SLOT_CAP_PHYSICAL_SLOT_NUM = 13'h0000;
  parameter SLOT_CAP_POWER_CONTROLLER_PRESENT = "FALSE";
  parameter SLOT_CAP_POWER_INDICATOR_PRESENT = "FALSE";
  parameter integer SLOT_CAP_SLOT_POWER_LIMIT_SCALE = 0;
  parameter [7:0] SLOT_CAP_SLOT_POWER_LIMIT_VALUE = 8'h00;
  parameter integer SPARE_BIT0 = 0;
  parameter integer SPARE_BIT1 = 0;
  parameter integer SPARE_BIT2 = 0;
  parameter integer SPARE_BIT3 = 0;
  parameter integer SPARE_BIT4 = 0;
  parameter integer SPARE_BIT5 = 0;
  parameter integer SPARE_BIT6 = 0;
  parameter integer SPARE_BIT7 = 0;
  parameter integer SPARE_BIT8 = 0;
  parameter [7:0] SPARE_BYTE0 = 8'h00;
  parameter [7:0] SPARE_BYTE1 = 8'h00;
  parameter [7:0] SPARE_BYTE2 = 8'h00;
  parameter [7:0] SPARE_BYTE3 = 8'h00;
  parameter [31:0] SPARE_WORD0 = 32'h00000000;
  parameter [31:0] SPARE_WORD1 = 32'h00000000;
  parameter [31:0] SPARE_WORD2 = 32'h00000000;
  parameter [31:0] SPARE_WORD3 = 32'h00000000;
  parameter SSL_MESSAGE_AUTO = "FALSE";
  parameter TECRC_EP_INV = "FALSE";
  parameter TL_RBYPASS = "FALSE";
  parameter integer TL_RX_RAM_RADDR_LATENCY = 0;
  parameter integer TL_RX_RAM_RDATA_LATENCY = 2;
  parameter integer TL_RX_RAM_WRITE_LATENCY = 0;
  parameter TL_TFC_DISABLE = "FALSE";
  parameter TL_TX_CHECKS_DISABLE = "FALSE";
  parameter integer TL_TX_RAM_RADDR_LATENCY = 0;
  parameter integer TL_TX_RAM_RDATA_LATENCY = 2;
  parameter integer TL_TX_RAM_WRITE_LATENCY = 0;
  parameter TRN_DW = "FALSE";
  parameter TRN_NP_FC = "FALSE";
  parameter UPCONFIG_CAPABLE = "TRUE";
  parameter UPSTREAM_FACING = "TRUE";
  parameter UR_ATOMIC = "TRUE";
  parameter UR_CFG1 = "TRUE";
  parameter UR_INV_REQ = "TRUE";
  parameter UR_PRS_RESPONSE = "TRUE";
  parameter USER_CLK2_DIV2 = "FALSE";
  parameter integer USER_CLK_FREQ = 3;
  parameter USE_RID_PINS = "FALSE";
  parameter VC0_CPL_INFINITE = "TRUE";
  parameter [12:0] VC0_RX_RAM_LIMIT = 13'h03FF;
  parameter integer VC0_TOTAL_CREDITS_CD = 127;
  parameter integer VC0_TOTAL_CREDITS_CH = 31;
  parameter integer VC0_TOTAL_CREDITS_NPD = 24;
  parameter integer VC0_TOTAL_CREDITS_NPH = 12;
  parameter integer VC0_TOTAL_CREDITS_PD = 288;
  parameter integer VC0_TOTAL_CREDITS_PH = 32;
  parameter integer VC0_TX_LASTPACKET = 31;
  parameter [11:0] VC_BASE_PTR = 12'h10C;
  parameter [15:0] VC_CAP_ID = 16'h0002;
  parameter [11:0] VC_CAP_NEXTPTR = 12'h000;
  parameter VC_CAP_ON = "FALSE";
  parameter VC_CAP_REJECT_SNOOP_TRANSACTIONS = "FALSE";
  parameter [3:0] VC_CAP_VERSION = 4'h1;
  parameter [11:0] VSEC_BASE_PTR = 12'h128;
  parameter [15:0] VSEC_CAP_HDR_ID = 16'h1234;
  parameter [11:0] VSEC_CAP_HDR_LENGTH = 12'h018;
  parameter [3:0] VSEC_CAP_HDR_REVISION = 4'h1;
  parameter [15:0] VSEC_CAP_ID = 16'h000B;
  parameter VSEC_CAP_IS_LINK_VISIBLE = "TRUE";
  parameter [11:0] VSEC_CAP_NEXTPTR = 12'h140;
  parameter VSEC_CAP_ON = "FALSE";
  parameter [3:0] VSEC_CAP_VERSION = 4'h1;
  
  localparam in_delay = 0;
  localparam out_delay = 0;
  localparam INCLK_DELAY = 0;
  localparam OUTCLK_DELAY = 0;

  output CFGAERECRCCHECKEN;
  output CFGAERECRCGENEN;
  output CFGAERROOTERRCORRERRRECEIVED;
  output CFGAERROOTERRCORRERRREPORTINGEN;
  output CFGAERROOTERRFATALERRRECEIVED;
  output CFGAERROOTERRFATALERRREPORTINGEN;
  output CFGAERROOTERRNONFATALERRRECEIVED;
  output CFGAERROOTERRNONFATALERRREPORTINGEN;
  output CFGBRIDGESERREN;
  output CFGCOMMANDBUSMASTERENABLE;
  output CFGCOMMANDINTERRUPTDISABLE;
  output CFGCOMMANDIOENABLE;
  output CFGCOMMANDMEMENABLE;
  output CFGCOMMANDSERREN;
  output CFGDEVCONTROL2ARIFORWARDEN;
  output CFGDEVCONTROL2ATOMICEGRESSBLOCK;
  output CFGDEVCONTROL2ATOMICREQUESTEREN;
  output CFGDEVCONTROL2CPLTIMEOUTDIS;
  output CFGDEVCONTROL2IDOCPLEN;
  output CFGDEVCONTROL2IDOREQEN;
  output CFGDEVCONTROL2LTREN;
  output CFGDEVCONTROL2TLPPREFIXBLOCK;
  output CFGDEVCONTROLAUXPOWEREN;
  output CFGDEVCONTROLCORRERRREPORTINGEN;
  output CFGDEVCONTROLENABLERO;
  output CFGDEVCONTROLEXTTAGEN;
  output CFGDEVCONTROLFATALERRREPORTINGEN;
  output CFGDEVCONTROLNONFATALREPORTINGEN;
  output CFGDEVCONTROLNOSNOOPEN;
  output CFGDEVCONTROLPHANTOMEN;
  output CFGDEVCONTROLURERRREPORTINGEN;
  output CFGDEVSTATUSCORRERRDETECTED;
  output CFGDEVSTATUSFATALERRDETECTED;
  output CFGDEVSTATUSNONFATALERRDETECTED;
  output CFGDEVSTATUSURDETECTED;
  output CFGERRAERHEADERLOGSETN;
  output CFGERRCPLRDYN;
  output CFGINTERRUPTMSIENABLE;
  output CFGINTERRUPTMSIXENABLE;
  output CFGINTERRUPTMSIXFM;
  output CFGINTERRUPTRDYN;
  output CFGLINKCONTROLAUTOBANDWIDTHINTEN;
  output CFGLINKCONTROLBANDWIDTHINTEN;
  output CFGLINKCONTROLCLOCKPMEN;
  output CFGLINKCONTROLCOMMONCLOCK;
  output CFGLINKCONTROLEXTENDEDSYNC;
  output CFGLINKCONTROLHWAUTOWIDTHDIS;
  output CFGLINKCONTROLLINKDISABLE;
  output CFGLINKCONTROLRCB;
  output CFGLINKCONTROLRETRAINLINK;
  output CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
  output CFGLINKSTATUSBANDWIDTHSTATUS;
  output CFGLINKSTATUSDLLACTIVE;
  output CFGLINKSTATUSLINKTRAINING;
  output CFGMGMTRDWRDONEN;
  output CFGMSGRECEIVED;
  output CFGMSGRECEIVEDASSERTINTA;
  output CFGMSGRECEIVEDASSERTINTB;
  output CFGMSGRECEIVEDASSERTINTC;
  output CFGMSGRECEIVEDASSERTINTD;
  output CFGMSGRECEIVEDDEASSERTINTA;
  output CFGMSGRECEIVEDDEASSERTINTB;
  output CFGMSGRECEIVEDDEASSERTINTC;
  output CFGMSGRECEIVEDDEASSERTINTD;
  output CFGMSGRECEIVEDERRCOR;
  output CFGMSGRECEIVEDERRFATAL;
  output CFGMSGRECEIVEDERRNONFATAL;
  output CFGMSGRECEIVEDPMASNAK;
  output CFGMSGRECEIVEDPMETO;
  output CFGMSGRECEIVEDPMETOACK;
  output CFGMSGRECEIVEDPMPME;
  output CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
  output CFGMSGRECEIVEDUNLOCK;
  output CFGPMCSRPMEEN;
  output CFGPMCSRPMESTATUS;
  output CFGPMRCVASREQL1N;
  output CFGPMRCVENTERL1N;
  output CFGPMRCVENTERL23N;
  output CFGPMRCVREQACKN;
  output CFGROOTCONTROLPMEINTEN;
  output CFGROOTCONTROLSYSERRCORRERREN;
  output CFGROOTCONTROLSYSERRFATALERREN;
  output CFGROOTCONTROLSYSERRNONFATALERREN;
  output CFGSLOTCONTROLELECTROMECHILCTLPULSE;
  output CFGTRANSACTION;
  output CFGTRANSACTIONTYPE;
  output DBGSCLRA;
  output DBGSCLRB;
  output DBGSCLRC;
  output DBGSCLRD;
  output DBGSCLRE;
  output DBGSCLRF;
  output DBGSCLRG;
  output DBGSCLRH;
  output DBGSCLRI;
  output DBGSCLRJ;
  output DBGSCLRK;
  output DRPRDY;
  output LL2BADDLLPERR;
  output LL2BADTLPERR;
  output LL2PROTOCOLERR;
  output LL2RECEIVERERR;
  output LL2REPLAYROERR;
  output LL2REPLAYTOERR;
  output LL2SUSPENDOK;
  output LL2TFCINIT1SEQ;
  output LL2TFCINIT2SEQ;
  output LL2TXIDLE;
  output LNKCLKEN;
  output MIMRXREN;
  output MIMRXWEN;
  output MIMTXREN;
  output MIMTXWEN;
  output PIPERX0POLARITY;
  output PIPERX1POLARITY;
  output PIPERX2POLARITY;
  output PIPERX3POLARITY;
  output PIPERX4POLARITY;
  output PIPERX5POLARITY;
  output PIPERX6POLARITY;
  output PIPERX7POLARITY;
  output PIPETX0COMPLIANCE;
  output PIPETX0ELECIDLE;
  output PIPETX1COMPLIANCE;
  output PIPETX1ELECIDLE;
  output PIPETX2COMPLIANCE;
  output PIPETX2ELECIDLE;
  output PIPETX3COMPLIANCE;
  output PIPETX3ELECIDLE;
  output PIPETX4COMPLIANCE;
  output PIPETX4ELECIDLE;
  output PIPETX5COMPLIANCE;
  output PIPETX5ELECIDLE;
  output PIPETX6COMPLIANCE;
  output PIPETX6ELECIDLE;
  output PIPETX7COMPLIANCE;
  output PIPETX7ELECIDLE;
  output PIPETXDEEMPH;
  output PIPETXRATE;
  output PIPETXRCVRDET;
  output PIPETXRESET;
  output PL2L0REQ;
  output PL2LINKUP;
  output PL2RECEIVERERR;
  output PL2RECOVERY;
  output PL2RXELECIDLE;
  output PL2SUSPENDOK;
  output PLDIRECTEDCHANGEDONE;
  output PLLINKGEN2CAP;
  output PLLINKPARTNERGEN2SUPPORTED;
  output PLLINKUPCFGCAP;
  output PLPHYLNKUPN;
  output PLRECEIVEDHOTRST;
  output PLSELLNKRATE;
  output RECEIVEDFUNCLVLRSTN;
  output TL2ASPMSUSPENDCREDITCHECKOK;
  output TL2ASPMSUSPENDREQ;
  output TL2ERRFCPE;
  output TL2ERRMALFORMED;
  output TL2ERRRXOVERFLOW;
  output TL2PPMSUSPENDOK;
  output TRNLNKUP;
  output TRNRECRCERR;
  output TRNREOF;
  output TRNRERRFWD;
  output TRNRSOF;
  output TRNRSRCDSC;
  output TRNRSRCRDY;
  output TRNTCFGREQ;
  output TRNTDLLPDSTRDY;
  output TRNTERRDROP;
  output USERRSTN;
  output [11:0] DBGVECC;
  output [11:0] PLDBGVEC;
  output [11:0] TRNFCCPLD;
  output [11:0] TRNFCNPD;
  output [11:0] TRNFCPD;
  output [127:0] TRNRD;
  output [12:0] MIMRXRADDR;
  output [12:0] MIMRXWADDR;
  output [12:0] MIMTXRADDR;
  output [12:0] MIMTXWADDR;
  output [15:0] CFGMSGDATA;
  output [15:0] DRPDO;
  output [15:0] PIPETX0DATA;
  output [15:0] PIPETX1DATA;
  output [15:0] PIPETX2DATA;
  output [15:0] PIPETX3DATA;
  output [15:0] PIPETX4DATA;
  output [15:0] PIPETX5DATA;
  output [15:0] PIPETX6DATA;
  output [15:0] PIPETX7DATA;
  output [1:0] CFGLINKCONTROLASPMCONTROL;
  output [1:0] CFGLINKSTATUSCURRENTSPEED;
  output [1:0] CFGPMCSRPOWERSTATE;
  output [1:0] PIPETX0CHARISK;
  output [1:0] PIPETX0POWERDOWN;
  output [1:0] PIPETX1CHARISK;
  output [1:0] PIPETX1POWERDOWN;
  output [1:0] PIPETX2CHARISK;
  output [1:0] PIPETX2POWERDOWN;
  output [1:0] PIPETX3CHARISK;
  output [1:0] PIPETX3POWERDOWN;
  output [1:0] PIPETX4CHARISK;
  output [1:0] PIPETX4POWERDOWN;
  output [1:0] PIPETX5CHARISK;
  output [1:0] PIPETX5POWERDOWN;
  output [1:0] PIPETX6CHARISK;
  output [1:0] PIPETX6POWERDOWN;
  output [1:0] PIPETX7CHARISK;
  output [1:0] PIPETX7POWERDOWN;
  output [1:0] PL2RXPMSTATE;
  output [1:0] PLLANEREVERSALMODE;
  output [1:0] PLRXPMSTATE;
  output [1:0] PLSELLNKWIDTH;
  output [1:0] TRNRDLLPSRCRDY;
  output [1:0] TRNRREM;
  output [2:0] CFGDEVCONTROLMAXPAYLOAD;
  output [2:0] CFGDEVCONTROLMAXREADREQ;
  output [2:0] CFGINTERRUPTMMENABLE;
  output [2:0] CFGPCIELINKSTATE;
  output [2:0] PIPETXMARGIN;
  output [2:0] PLINITIALLINKWIDTH;
  output [2:0] PLTXPMSTATE;
  output [31:0] CFGMGMTDO;
  output [3:0] CFGDEVCONTROL2CPLTIMEOUTVAL;
  output [3:0] CFGLINKSTATUSNEGOTIATEDWIDTH;
  output [3:0] TRNTDSTRDY;
  output [4:0] LL2LINKSTATUS;
  output [5:0] PLLTSSMSTATE;
  output [5:0] TRNTBUFAV;
  output [63:0] DBGVECA;
  output [63:0] DBGVECB;
  output [63:0] TL2ERRHDR;
  output [63:0] TRNRDLLPDATA;
  output [67:0] MIMRXWDATA;
  output [68:0] MIMTXWDATA;
  output [6:0] CFGTRANSACTIONADDR;
  output [6:0] CFGVCTCVCMAP;
  output [7:0] CFGINTERRUPTDO;
  output [7:0] TRNFCCPLH;
  output [7:0] TRNFCNPH;
  output [7:0] TRNFCPH;
  output [7:0] TRNRBARHIT;

  input CFGERRACSN;
  input CFGERRATOMICEGRESSBLOCKEDN;
  input CFGERRCORN;
  input CFGERRCPLABORTN;
  input CFGERRCPLTIMEOUTN;
  input CFGERRCPLUNEXPECTN;
  input CFGERRECRCN;
  input CFGERRINTERNALCORN;
  input CFGERRINTERNALUNCORN;
  input CFGERRLOCKEDN;
  input CFGERRMALFORMEDN;
  input CFGERRMCBLOCKEDN;
  input CFGERRNORECOVERYN;
  input CFGERRPOISONEDN;
  input CFGERRPOSTEDN;
  input CFGERRURN;
  input CFGFORCECOMMONCLOCKOFF;
  input CFGFORCEEXTENDEDSYNCON;
  input CFGINTERRUPTASSERTN;
  input CFGINTERRUPTN;
  input CFGINTERRUPTSTATN;
  input CFGMGMTRDENN;
  input CFGMGMTWRENN;
  input CFGMGMTWRREADONLYN;
  input CFGMGMTWRRW1CASRWN;
  input CFGPMFORCESTATEENN;
  input CFGPMHALTASPML0SN;
  input CFGPMHALTASPML1N;
  input CFGPMSENDPMETON;
  input CFGPMTURNOFFOKN;
  input CFGPMWAKEN;
  input CFGTRNPENDINGN;
  input CMRSTN;
  input CMSTICKYRSTN;
  input DBGSUBMODE;
  input DLRSTN;
  input DRPCLK;
  input DRPEN;
  input DRPWE;
  input FUNCLVLRSTN;
  input LL2SENDASREQL1;
  input LL2SENDENTERL1;
  input LL2SENDENTERL23;
  input LL2SENDPMACK;
  input LL2SUSPENDNOW;
  input LL2TLPRCV;
  input PIPECLK;
  input PIPERX0CHANISALIGNED;
  input PIPERX0ELECIDLE;
  input PIPERX0PHYSTATUS;
  input PIPERX0VALID;
  input PIPERX1CHANISALIGNED;
  input PIPERX1ELECIDLE;
  input PIPERX1PHYSTATUS;
  input PIPERX1VALID;
  input PIPERX2CHANISALIGNED;
  input PIPERX2ELECIDLE;
  input PIPERX2PHYSTATUS;
  input PIPERX2VALID;
  input PIPERX3CHANISALIGNED;
  input PIPERX3ELECIDLE;
  input PIPERX3PHYSTATUS;
  input PIPERX3VALID;
  input PIPERX4CHANISALIGNED;
  input PIPERX4ELECIDLE;
  input PIPERX4PHYSTATUS;
  input PIPERX4VALID;
  input PIPERX5CHANISALIGNED;
  input PIPERX5ELECIDLE;
  input PIPERX5PHYSTATUS;
  input PIPERX5VALID;
  input PIPERX6CHANISALIGNED;
  input PIPERX6ELECIDLE;
  input PIPERX6PHYSTATUS;
  input PIPERX6VALID;
  input PIPERX7CHANISALIGNED;
  input PIPERX7ELECIDLE;
  input PIPERX7PHYSTATUS;
  input PIPERX7VALID;
  input PLDIRECTEDLINKAUTON;
  input PLDIRECTEDLINKSPEED;
  input PLDIRECTEDLTSSMNEWVLD;
  input PLDIRECTEDLTSSMSTALL;
  input PLDOWNSTREAMDEEMPHSOURCE;
  input PLRSTN;
  input PLTRANSMITHOTRST;
  input PLUPSTREAMPREFERDEEMPH;
  input SYSRSTN;
  input TL2ASPMSUSPENDCREDITCHECK;
  input TL2PPMSUSPENDREQ;
  input TLRSTN;
  input TRNRDSTRDY;
  input TRNRFCPRET;
  input TRNRNPOK;
  input TRNRNPREQ;
  input TRNTCFGGNT;
  input TRNTDLLPSRCRDY;
  input TRNTECRCGEN;
  input TRNTEOF;
  input TRNTERRFWD;
  input TRNTSOF;
  input TRNTSRCDSC;
  input TRNTSRCRDY;
  input TRNTSTR;
  input USERCLK2;
  input USERCLK;
  input [127:0] CFGERRAERHEADERLOG;
  input [127:0] TRNTD;
  input [15:0] CFGDEVID;
  input [15:0] CFGSUBSYSID;
  input [15:0] CFGSUBSYSVENDID;
  input [15:0] CFGVENDID;
  input [15:0] DRPDI;
  input [15:0] PIPERX0DATA;
  input [15:0] PIPERX1DATA;
  input [15:0] PIPERX2DATA;
  input [15:0] PIPERX3DATA;
  input [15:0] PIPERX4DATA;
  input [15:0] PIPERX5DATA;
  input [15:0] PIPERX6DATA;
  input [15:0] PIPERX7DATA;
  input [1:0] CFGPMFORCESTATE;
  input [1:0] DBGMODE;
  input [1:0] PIPERX0CHARISK;
  input [1:0] PIPERX1CHARISK;
  input [1:0] PIPERX2CHARISK;
  input [1:0] PIPERX3CHARISK;
  input [1:0] PIPERX4CHARISK;
  input [1:0] PIPERX5CHARISK;
  input [1:0] PIPERX6CHARISK;
  input [1:0] PIPERX7CHARISK;
  input [1:0] PLDIRECTEDLINKCHANGE;
  input [1:0] PLDIRECTEDLINKWIDTH;
  input [1:0] TRNTREM;
  input [2:0] CFGDSFUNCTIONNUMBER;
  input [2:0] CFGFORCEMPS;
  input [2:0] PIPERX0STATUS;
  input [2:0] PIPERX1STATUS;
  input [2:0] PIPERX2STATUS;
  input [2:0] PIPERX3STATUS;
  input [2:0] PIPERX4STATUS;
  input [2:0] PIPERX5STATUS;
  input [2:0] PIPERX6STATUS;
  input [2:0] PIPERX7STATUS;
  input [2:0] PLDBGMODE;
  input [2:0] TRNFCSEL;
  input [31:0] CFGMGMTDI;
  input [31:0] TRNTDLLPDATA;
  input [3:0] CFGMGMTBYTEENN;
  input [47:0] CFGERRTLPCPLHEADER;
  input [4:0] CFGAERINTERRUPTMSGNUM;
  input [4:0] CFGDSDEVICENUMBER;
  input [4:0] CFGPCIECAPINTERRUPTMSGNUM;
  input [4:0] PL2DIRECTEDLSTATE;
  input [5:0] PLDIRECTEDLTSSMNEW;
  input [63:0] CFGDSN;
  input [67:0] MIMRXRDATA;
  input [68:0] MIMTXRDATA;
  input [7:0] CFGDSBUSNUMBER;
  input [7:0] CFGINTERRUPTDI;
  input [7:0] CFGPORTNUMBER;
  input [7:0] CFGREVID;
  input [8:0] DRPADDR;
  input [9:0] CFGMGMTDWADDR;

  reg SIM_VERSION_BINARY;
  reg [0:0] AER_CAP_ECRC_CHECK_CAPABLE_BINARY;
  reg [0:0] AER_CAP_ECRC_GEN_CAPABLE_BINARY;
  reg [0:0] AER_CAP_MULTIHEADER_BINARY;
  reg [0:0] AER_CAP_ON_BINARY;
  reg [0:0] AER_CAP_PERMIT_ROOTERR_UPDATE_BINARY;
  reg [0:0] ALLOW_X8_GEN2_BINARY;
  reg [0:0] CMD_INTX_IMPLEMENTED_BINARY;
  reg [0:0] CPL_TIMEOUT_DISABLE_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_ARI_FORWARDING_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_CAS128_COMPLETER_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_LTR_MECHANISM_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING_BINARY;
  reg [0:0] DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE_BINARY;
  reg [0:0] DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE_BINARY;
  reg [0:0] DEV_CAP_EXT_TAG_SUPPORTED_BINARY;
  reg [0:0] DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY;
  reg [0:0] DEV_CAP_ROLE_BASED_ERROR_BINARY;
  reg [0:0] DEV_CONTROL_AUX_POWER_SUPPORTED_BINARY;
  reg [0:0] DEV_CONTROL_EXT_TAG_DEFAULT_BINARY;
  reg [0:0] DISABLE_ASPM_L1_TIMER_BINARY;
  reg [0:0] DISABLE_BAR_FILTERING_BINARY;
  reg [0:0] DISABLE_ERR_MSG_BINARY;
  reg [0:0] DISABLE_ID_CHECK_BINARY;
  reg [0:0] DISABLE_LANE_REVERSAL_BINARY;
  reg [0:0] DISABLE_LOCKED_FILTER_BINARY;
  reg [0:0] DISABLE_PPM_FILTER_BINARY;
  reg [0:0] DISABLE_RX_POISONED_RESP_BINARY;
  reg [0:0] DISABLE_RX_TC_FILTER_BINARY;
  reg [0:0] DISABLE_SCRAMBLING_BINARY;
  reg [0:0] DSN_CAP_ON_BINARY;
  reg [0:0] ENABLE_RX_TD_ECRC_TRIM_BINARY;
  reg [0:0] ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED_BINARY;
  reg [0:0] ENTER_RVRY_EI_L0_BINARY;
  reg [0:0] EXIT_LOOPBACK_ON_EI_BINARY;
  reg [0:0] INTERRUPT_STAT_AUTO_BINARY;
  reg [0:0] IS_SWITCH_BINARY;
  reg [0:0] LINK_CAP_ASPM_OPTIONALITY_BINARY;
  reg [0:0] LINK_CAP_CLOCK_POWER_MANAGEMENT_BINARY;
  reg [0:0] LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP_BINARY;
  reg [0:0] LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP_BINARY;
  reg [0:0] LINK_CAP_RSVD_23_BINARY;
  reg [0:0] LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE_BINARY;
  reg [0:0] LINK_CONTROL_RCB_BINARY;
  reg [0:0] LINK_CTRL2_DEEMPHASIS_BINARY;
  reg [0:0] LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE_BINARY;
  reg [0:0] LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY;
  reg [0:0] LL_ACK_TIMEOUT_EN_BINARY;
  reg [0:0] LL_REPLAY_TIMEOUT_EN_BINARY;
  reg [0:0] MPS_FORCE_BINARY;
  reg [0:0] MSIX_CAP_ON_BINARY;
  reg [0:0] MSI_CAP_64_BIT_ADDR_CAPABLE_BINARY;
  reg [0:0] MSI_CAP_MULTIMSG_EXTENSION_BINARY;
  reg [0:0] MSI_CAP_ON_BINARY;
  reg [0:0] MSI_CAP_PER_VECTOR_MASKING_CAPABLE_BINARY;
  reg [0:0] PCIE_CAP_ON_BINARY;
  reg [0:0] PCIE_CAP_SLOT_IMPLEMENTED_BINARY;
  reg [0:0] PL_FAST_TRAIN_BINARY;
  reg [0:0] PM_ASPML0S_TIMEOUT_EN_BINARY;
  reg [0:0] PM_ASPM_FASTEXIT_BINARY;
  reg [0:0] PM_CAP_D1SUPPORT_BINARY;
  reg [0:0] PM_CAP_D2SUPPORT_BINARY;
  reg [0:0] PM_CAP_DSI_BINARY;
  reg [0:0] PM_CAP_ON_BINARY;
  reg [0:0] PM_CAP_PME_CLOCK_BINARY;
  reg [0:0] PM_CAP_RSVD_04_BINARY;
  reg [0:0] PM_CSR_B2B3_BINARY;
  reg [0:0] PM_CSR_BPCCEN_BINARY;
  reg [0:0] PM_CSR_NOSOFTRST_BINARY;
  reg [0:0] PM_MF_BINARY;
  reg [0:0] RBAR_CAP_ON_BINARY;
  reg [0:0] RECRC_CHK_TRIM_BINARY;
  reg [0:0] ROOT_CAP_CRS_SW_VISIBILITY_BINARY;
  reg [0:0] SELECT_DLL_IF_BINARY;
  reg [0:0] SLOT_CAP_ATT_BUTTON_PRESENT_BINARY;
  reg [0:0] SLOT_CAP_ATT_INDICATOR_PRESENT_BINARY;
  reg [0:0] SLOT_CAP_ELEC_INTERLOCK_PRESENT_BINARY;
  reg [0:0] SLOT_CAP_HOTPLUG_CAPABLE_BINARY;
  reg [0:0] SLOT_CAP_HOTPLUG_SURPRISE_BINARY;
  reg [0:0] SLOT_CAP_MRL_SENSOR_PRESENT_BINARY;
  reg [0:0] SLOT_CAP_NO_CMD_COMPLETED_SUPPORT_BINARY;
  reg [0:0] SLOT_CAP_POWER_CONTROLLER_PRESENT_BINARY;
  reg [0:0] SLOT_CAP_POWER_INDICATOR_PRESENT_BINARY;
  reg [0:0] SPARE_BIT0_BINARY;
  reg [0:0] SPARE_BIT1_BINARY;
  reg [0:0] SPARE_BIT2_BINARY;
  reg [0:0] SPARE_BIT3_BINARY;
  reg [0:0] SPARE_BIT4_BINARY;
  reg [0:0] SPARE_BIT5_BINARY;
  reg [0:0] SPARE_BIT6_BINARY;
  reg [0:0] SPARE_BIT7_BINARY;
  reg [0:0] SPARE_BIT8_BINARY;
  reg [0:0] SSL_MESSAGE_AUTO_BINARY;
  reg [0:0] TECRC_EP_INV_BINARY;
  reg [0:0] TL_RBYPASS_BINARY;
  reg [0:0] TL_RX_RAM_RADDR_LATENCY_BINARY;
  reg [0:0] TL_RX_RAM_WRITE_LATENCY_BINARY;
  reg [0:0] TL_TFC_DISABLE_BINARY;
  reg [0:0] TL_TX_CHECKS_DISABLE_BINARY;
  reg [0:0] TL_TX_RAM_RADDR_LATENCY_BINARY;
  reg [0:0] TL_TX_RAM_WRITE_LATENCY_BINARY;
  reg [0:0] TRN_DW_BINARY;
  reg [0:0] TRN_NP_FC_BINARY;
  reg [0:0] UPCONFIG_CAPABLE_BINARY;
  reg [0:0] UPSTREAM_FACING_BINARY;
  reg [0:0] UR_ATOMIC_BINARY;
  reg [0:0] UR_CFG1_BINARY;
  reg [0:0] UR_INV_REQ_BINARY;
  reg [0:0] UR_PRS_RESPONSE_BINARY;
  reg [0:0] USER_CLK2_DIV2_BINARY;
  reg [0:0] USE_RID_PINS_BINARY;
  reg [0:0] VC0_CPL_INFINITE_BINARY;
  reg [0:0] VC_CAP_ON_BINARY;
  reg [0:0] VC_CAP_REJECT_SNOOP_TRANSACTIONS_BINARY;
  reg [0:0] VSEC_CAP_IS_LINK_VISIBLE_BINARY;
  reg [0:0] VSEC_CAP_ON_BINARY;
  reg [10:0] VC0_TOTAL_CREDITS_CD_BINARY;
  reg [10:0] VC0_TOTAL_CREDITS_NPD_BINARY;
  reg [10:0] VC0_TOTAL_CREDITS_PD_BINARY;
  reg [1:0] CFG_ECRC_ERR_CPLSTAT_BINARY;
  reg [1:0] DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT_BINARY;
  reg [1:0] DEV_CAP_RSVD_17_16_BINARY;
  reg [1:0] LINK_CAP_ASPM_SUPPORT_BINARY;
  reg [1:0] LL_ACK_TIMEOUT_FUNC_BINARY;
  reg [1:0] LL_REPLAY_TIMEOUT_FUNC_BINARY;
  reg [1:0] PCIE_CAP_RSVD_15_14_BINARY;
  reg [1:0] PM_ASPML0S_TIMEOUT_FUNC_BINARY;
  reg [1:0] RECRC_CHK_BINARY;
  reg [1:0] SLOT_CAP_SLOT_POWER_LIMIT_SCALE_BINARY;
  reg [1:0] TL_RX_RAM_RDATA_LATENCY_BINARY;
  reg [1:0] TL_TX_RAM_RDATA_LATENCY_BINARY;
  reg [2:0] DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY;
  reg [2:0] DEV_CAP_ENDPOINT_L1_LATENCY_BINARY;
  reg [2:0] DEV_CAP_MAX_PAYLOAD_SUPPORTED_BINARY;
  reg [2:0] DEV_CAP_RSVD_14_12_BINARY;
  reg [2:0] DEV_CAP_RSVD_31_29_BINARY;
  reg [2:0] LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] PL_AUTO_CONFIG_BINARY;
  reg [2:0] PM_CAP_AUXCURRENT_BINARY;
  reg [2:0] PM_CAP_VERSION_BINARY;
  reg [2:0] USER_CLK_FREQ_BINARY;
  reg [3:0] PCIE_REVISION_BINARY;
  reg [4:0] VC0_TX_LASTPACKET_BINARY;
  reg [6:0] VC0_TOTAL_CREDITS_CH_BINARY;
  reg [6:0] VC0_TOTAL_CREDITS_NPH_BINARY;
  reg [6:0] VC0_TOTAL_CREDITS_PH_BINARY;
  reg [7:0] N_FTS_COMCLK_GEN1_BINARY;
  reg [7:0] N_FTS_COMCLK_GEN2_BINARY;
  reg [7:0] N_FTS_GEN1_BINARY;
  reg [7:0] N_FTS_GEN2_BINARY;

//  tri0 GSR = glbl.GSR;
  reg notifier;

  initial begin
    case (AER_CAP_ECRC_CHECK_CAPABLE)
      "FALSE" : AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b0;
      "TRUE" : AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AER_CAP_ECRC_CHECK_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AER_CAP_ECRC_CHECK_CAPABLE);
        #1 $finish;
      end
    endcase

    case (AER_CAP_ECRC_GEN_CAPABLE)
      "FALSE" : AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b0;
      "TRUE" : AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AER_CAP_ECRC_GEN_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AER_CAP_ECRC_GEN_CAPABLE);
        #1 $finish;
      end
    endcase

    case (AER_CAP_MULTIHEADER)
      "FALSE" : AER_CAP_MULTIHEADER_BINARY = 1'b0;
      "TRUE" : AER_CAP_MULTIHEADER_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AER_CAP_MULTIHEADER on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AER_CAP_MULTIHEADER);
        #1 $finish;
      end
    endcase

    case (AER_CAP_ON)
      "FALSE" : AER_CAP_ON_BINARY = 1'b0;
      "TRUE" : AER_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AER_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AER_CAP_ON);
        #1 $finish;
      end
    endcase

    case (AER_CAP_PERMIT_ROOTERR_UPDATE)
      "TRUE" : AER_CAP_PERMIT_ROOTERR_UPDATE_BINARY = 1'b1;
      "FALSE" : AER_CAP_PERMIT_ROOTERR_UPDATE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute AER_CAP_PERMIT_ROOTERR_UPDATE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", AER_CAP_PERMIT_ROOTERR_UPDATE);
        #1 $finish;
      end
    endcase

    case (ALLOW_X8_GEN2)
      "FALSE" : ALLOW_X8_GEN2_BINARY = 1'b0;
      "TRUE" : ALLOW_X8_GEN2_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ALLOW_X8_GEN2 on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ALLOW_X8_GEN2);
        #1 $finish;
      end
    endcase

    case (CMD_INTX_IMPLEMENTED)
      "TRUE" : CMD_INTX_IMPLEMENTED_BINARY = 1'b1;
      "FALSE" : CMD_INTX_IMPLEMENTED_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CMD_INTX_IMPLEMENTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", CMD_INTX_IMPLEMENTED);
        #1 $finish;
      end
    endcase

    case (CPL_TIMEOUT_DISABLE_SUPPORTED)
      "FALSE" : CPL_TIMEOUT_DISABLE_SUPPORTED_BINARY = 1'b0;
      "TRUE" : CPL_TIMEOUT_DISABLE_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute CPL_TIMEOUT_DISABLE_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", CPL_TIMEOUT_DISABLE_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_ARI_FORWARDING_SUPPORTED)
      "FALSE" : DEV_CAP2_ARI_FORWARDING_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_ARI_FORWARDING_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_ARI_FORWARDING_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_ARI_FORWARDING_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED)
      "FALSE" : DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED)
      "FALSE" : DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED)
      "FALSE" : DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_CAS128_COMPLETER_SUPPORTED)
      "FALSE" : DEV_CAP2_CAS128_COMPLETER_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_CAS128_COMPLETER_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_CAS128_COMPLETER_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_CAS128_COMPLETER_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED)
      "FALSE" : DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED)
      "FALSE" : DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_LTR_MECHANISM_SUPPORTED)
      "FALSE" : DEV_CAP2_LTR_MECHANISM_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_LTR_MECHANISM_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_LTR_MECHANISM_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_LTR_MECHANISM_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING)
      "FALSE" : DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING_BINARY = 1'b0;
      "TRUE" : DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING);
        #1 $finish;
      end
    endcase

    case (DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE)
      "TRUE" : DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE_BINARY = 1'b1;
      "FALSE" : DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE);
        #1 $finish;
      end
    endcase

    case (DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE)
      "TRUE" : DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE_BINARY = 1'b1;
      "FALSE" : DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE);
        #1 $finish;
      end
    endcase

    case (DEV_CAP_EXT_TAG_SUPPORTED)
      "TRUE" : DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b1;
      "FALSE" : DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP_EXT_TAG_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEV_CAP_EXT_TAG_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
      "FALSE" : DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b0;
      "TRUE" : DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE);
        #1 $finish;
      end
    endcase

    case (DEV_CAP_ROLE_BASED_ERROR)
      "TRUE" : DEV_CAP_ROLE_BASED_ERROR_BINARY = 1'b1;
      "FALSE" : DEV_CAP_ROLE_BASED_ERROR_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CAP_ROLE_BASED_ERROR on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DEV_CAP_ROLE_BASED_ERROR);
        #1 $finish;
      end
    endcase

    case (DEV_CONTROL_AUX_POWER_SUPPORTED)
      "FALSE" : DEV_CONTROL_AUX_POWER_SUPPORTED_BINARY = 1'b0;
      "TRUE" : DEV_CONTROL_AUX_POWER_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CONTROL_AUX_POWER_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CONTROL_AUX_POWER_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (DEV_CONTROL_EXT_TAG_DEFAULT)
      "FALSE" : DEV_CONTROL_EXT_TAG_DEFAULT_BINARY = 1'b0;
      "TRUE" : DEV_CONTROL_EXT_TAG_DEFAULT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DEV_CONTROL_EXT_TAG_DEFAULT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DEV_CONTROL_EXT_TAG_DEFAULT);
        #1 $finish;
      end
    endcase

    case (DISABLE_ASPM_L1_TIMER)
      "FALSE" : DISABLE_ASPM_L1_TIMER_BINARY = 1'b0;
      "TRUE" : DISABLE_ASPM_L1_TIMER_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_ASPM_L1_TIMER on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_ASPM_L1_TIMER);
        #1 $finish;
      end
    endcase

    case (DISABLE_BAR_FILTERING)
      "FALSE" : DISABLE_BAR_FILTERING_BINARY = 1'b0;
      "TRUE" : DISABLE_BAR_FILTERING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_BAR_FILTERING on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_BAR_FILTERING);
        #1 $finish;
      end
    endcase

    case (DISABLE_ERR_MSG)
      "FALSE" : DISABLE_ERR_MSG_BINARY = 1'b0;
      "TRUE" : DISABLE_ERR_MSG_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_ERR_MSG on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_ERR_MSG);
        #1 $finish;
      end
    endcase

    case (DISABLE_ID_CHECK)
      "FALSE" : DISABLE_ID_CHECK_BINARY = 1'b0;
      "TRUE" : DISABLE_ID_CHECK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_ID_CHECK on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_ID_CHECK);
        #1 $finish;
      end
    endcase

    case (DISABLE_LANE_REVERSAL)
      "FALSE" : DISABLE_LANE_REVERSAL_BINARY = 1'b0;
      "TRUE" : DISABLE_LANE_REVERSAL_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_LANE_REVERSAL on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_LANE_REVERSAL);
        #1 $finish;
      end
    endcase

    case (DISABLE_LOCKED_FILTER)
      "FALSE" : DISABLE_LOCKED_FILTER_BINARY = 1'b0;
      "TRUE" : DISABLE_LOCKED_FILTER_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_LOCKED_FILTER on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_LOCKED_FILTER);
        #1 $finish;
      end
    endcase

    case (DISABLE_PPM_FILTER)
      "FALSE" : DISABLE_PPM_FILTER_BINARY = 1'b0;
      "TRUE" : DISABLE_PPM_FILTER_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_PPM_FILTER on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_PPM_FILTER);
        #1 $finish;
      end
    endcase

    case (DISABLE_RX_POISONED_RESP)
      "FALSE" : DISABLE_RX_POISONED_RESP_BINARY = 1'b0;
      "TRUE" : DISABLE_RX_POISONED_RESP_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_RX_POISONED_RESP on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_RX_POISONED_RESP);
        #1 $finish;
      end
    endcase

    case (DISABLE_RX_TC_FILTER)
      "FALSE" : DISABLE_RX_TC_FILTER_BINARY = 1'b0;
      "TRUE" : DISABLE_RX_TC_FILTER_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_RX_TC_FILTER on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_RX_TC_FILTER);
        #1 $finish;
      end
    endcase

    case (DISABLE_SCRAMBLING)
      "FALSE" : DISABLE_SCRAMBLING_BINARY = 1'b0;
      "TRUE" : DISABLE_SCRAMBLING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute DISABLE_SCRAMBLING on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", DISABLE_SCRAMBLING);
        #1 $finish;
      end
    endcase

    case (DSN_CAP_ON)
      "TRUE" : DSN_CAP_ON_BINARY = 1'b1;
      "FALSE" : DSN_CAP_ON_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute DSN_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", DSN_CAP_ON);
        #1 $finish;
      end
    endcase

    case (ENABLE_RX_TD_ECRC_TRIM)
      "FALSE" : ENABLE_RX_TD_ECRC_TRIM_BINARY = 1'b0;
      "TRUE" : ENABLE_RX_TD_ECRC_TRIM_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ENABLE_RX_TD_ECRC_TRIM on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ENABLE_RX_TD_ECRC_TRIM);
        #1 $finish;
      end
    endcase

    case (ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED)
      "FALSE" : ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED_BINARY = 1'b0;
      "TRUE" : ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED);
        #1 $finish;
      end
    endcase

    case (ENTER_RVRY_EI_L0)
      "TRUE" : ENTER_RVRY_EI_L0_BINARY = 1'b1;
      "FALSE" : ENTER_RVRY_EI_L0_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute ENTER_RVRY_EI_L0 on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", ENTER_RVRY_EI_L0);
        #1 $finish;
      end
    endcase

    case (EXIT_LOOPBACK_ON_EI)
      "TRUE" : EXIT_LOOPBACK_ON_EI_BINARY = 1'b1;
      "FALSE" : EXIT_LOOPBACK_ON_EI_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute EXIT_LOOPBACK_ON_EI on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", EXIT_LOOPBACK_ON_EI);
        #1 $finish;
      end
    endcase

    case (INTERRUPT_STAT_AUTO)
      "TRUE" : INTERRUPT_STAT_AUTO_BINARY = 1'b1;
      "FALSE" : INTERRUPT_STAT_AUTO_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute INTERRUPT_STAT_AUTO on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", INTERRUPT_STAT_AUTO);
        #1 $finish;
      end
    endcase

    case (IS_SWITCH)
      "FALSE" : IS_SWITCH_BINARY = 1'b0;
      "TRUE" : IS_SWITCH_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute IS_SWITCH on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", IS_SWITCH);
        #1 $finish;
      end
    endcase

    case (LINK_CAP_ASPM_OPTIONALITY)
      "TRUE" : LINK_CAP_ASPM_OPTIONALITY_BINARY = 1'b1;
      "FALSE" : LINK_CAP_ASPM_OPTIONALITY_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CAP_ASPM_OPTIONALITY on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", LINK_CAP_ASPM_OPTIONALITY);
        #1 $finish;
      end
    endcase

    case (LINK_CAP_CLOCK_POWER_MANAGEMENT)
      "FALSE" : LINK_CAP_CLOCK_POWER_MANAGEMENT_BINARY = 1'b0;
      "TRUE" : LINK_CAP_CLOCK_POWER_MANAGEMENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CAP_CLOCK_POWER_MANAGEMENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CAP_CLOCK_POWER_MANAGEMENT);
        #1 $finish;
      end
    endcase

    case (LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP)
      "FALSE" : LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP_BINARY = 1'b0;
      "TRUE" : LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP);
        #1 $finish;
      end
    endcase

    case (LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP)
      "FALSE" : LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP_BINARY = 1'b0;
      "TRUE" : LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP);
        #1 $finish;
      end
    endcase

    case (LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE)
      "FALSE" : LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE_BINARY = 1'b0;
      "TRUE" : LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE);
        #1 $finish;
      end
    endcase

    case (LINK_CTRL2_DEEMPHASIS)
      "FALSE" : LINK_CTRL2_DEEMPHASIS_BINARY = 1'b0;
      "TRUE" : LINK_CTRL2_DEEMPHASIS_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CTRL2_DEEMPHASIS on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CTRL2_DEEMPHASIS);
        #1 $finish;
      end
    endcase

    case (LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE)
      "FALSE" : LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE_BINARY = 1'b0;
      "TRUE" : LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE);
        #1 $finish;
      end
    endcase

    case (LINK_STATUS_SLOT_CLOCK_CONFIG)
      "TRUE" : LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b1;
      "FALSE" : LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute LINK_STATUS_SLOT_CLOCK_CONFIG on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", LINK_STATUS_SLOT_CLOCK_CONFIG);
        #1 $finish;
      end
    endcase

    case (LL_ACK_TIMEOUT_EN)
      "FALSE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_EN on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_ACK_TIMEOUT_EN);
        #1 $finish;
      end
    endcase

    case (LL_REPLAY_TIMEOUT_EN)
      "FALSE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_EN on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_REPLAY_TIMEOUT_EN);
        #1 $finish;
      end
    endcase

    case (MPS_FORCE)
      "FALSE" : MPS_FORCE_BINARY = 1'b0;
      "TRUE" : MPS_FORCE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute MPS_FORCE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", MPS_FORCE);
        #1 $finish;
      end
    endcase

    case (MSIX_CAP_ON)
      "FALSE" : MSIX_CAP_ON_BINARY = 1'b0;
      "TRUE" : MSIX_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute MSIX_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", MSIX_CAP_ON);
        #1 $finish;
      end
    endcase

    case (MSI_CAP_64_BIT_ADDR_CAPABLE)
      "TRUE" : MSI_CAP_64_BIT_ADDR_CAPABLE_BINARY = 1'b1;
      "FALSE" : MSI_CAP_64_BIT_ADDR_CAPABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute MSI_CAP_64_BIT_ADDR_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", MSI_CAP_64_BIT_ADDR_CAPABLE);
        #1 $finish;
      end
    endcase

    case (MSI_CAP_ON)
      "FALSE" : MSI_CAP_ON_BINARY = 1'b0;
      "TRUE" : MSI_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute MSI_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", MSI_CAP_ON);
        #1 $finish;
      end
    endcase

    case (MSI_CAP_PER_VECTOR_MASKING_CAPABLE)
      "TRUE" : MSI_CAP_PER_VECTOR_MASKING_CAPABLE_BINARY = 1'b1;
      "FALSE" : MSI_CAP_PER_VECTOR_MASKING_CAPABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute MSI_CAP_PER_VECTOR_MASKING_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", MSI_CAP_PER_VECTOR_MASKING_CAPABLE);
        #1 $finish;
      end
    endcase

    case (PCIE_CAP_ON)
      "TRUE" : PCIE_CAP_ON_BINARY = 1'b1;
      "FALSE" : PCIE_CAP_ON_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PCIE_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PCIE_CAP_ON);
        #1 $finish;
      end
    endcase

    case (PCIE_CAP_SLOT_IMPLEMENTED)
      "FALSE" : PCIE_CAP_SLOT_IMPLEMENTED_BINARY = 1'b0;
      "TRUE" : PCIE_CAP_SLOT_IMPLEMENTED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PCIE_CAP_SLOT_IMPLEMENTED on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PCIE_CAP_SLOT_IMPLEMENTED);
        #1 $finish;
      end
    endcase

    case (PL_FAST_TRAIN)
      "FALSE" : PL_FAST_TRAIN_BINARY = 1'b0;
      "TRUE" : PL_FAST_TRAIN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_FAST_TRAIN on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_FAST_TRAIN);
        #1 $finish;
      end
    endcase

    case (PM_ASPML0S_TIMEOUT_EN)
      "FALSE" : PM_ASPML0S_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : PM_ASPML0S_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_ASPML0S_TIMEOUT_EN on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_ASPML0S_TIMEOUT_EN);
        #1 $finish;
      end
    endcase

    case (PM_ASPM_FASTEXIT)
      "FALSE" : PM_ASPM_FASTEXIT_BINARY = 1'b0;
      "TRUE" : PM_ASPM_FASTEXIT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_ASPM_FASTEXIT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_ASPM_FASTEXIT);
        #1 $finish;
      end
    endcase

    case (PM_CAP_D1SUPPORT)
      "TRUE" : PM_CAP_D1SUPPORT_BINARY = 1'b1;
      "FALSE" : PM_CAP_D1SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CAP_D1SUPPORT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_CAP_D1SUPPORT);
        #1 $finish;
      end
    endcase

    case (PM_CAP_D2SUPPORT)
      "TRUE" : PM_CAP_D2SUPPORT_BINARY = 1'b1;
      "FALSE" : PM_CAP_D2SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CAP_D2SUPPORT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_CAP_D2SUPPORT);
        #1 $finish;
      end
    endcase

    case (PM_CAP_DSI)
      "FALSE" : PM_CAP_DSI_BINARY = 1'b0;
      "TRUE" : PM_CAP_DSI_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CAP_DSI on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_CAP_DSI);
        #1 $finish;
      end
    endcase

    case (PM_CAP_ON)
      "TRUE" : PM_CAP_ON_BINARY = 1'b1;
      "FALSE" : PM_CAP_ON_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_CAP_ON);
        #1 $finish;
      end
    endcase

    case (PM_CAP_PME_CLOCK)
      "FALSE" : PM_CAP_PME_CLOCK_BINARY = 1'b0;
      "TRUE" : PM_CAP_PME_CLOCK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CAP_PME_CLOCK on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_CAP_PME_CLOCK);
        #1 $finish;
      end
    endcase

    case (PM_CSR_B2B3)
      "FALSE" : PM_CSR_B2B3_BINARY = 1'b0;
      "TRUE" : PM_CSR_B2B3_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CSR_B2B3 on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_CSR_B2B3);
        #1 $finish;
      end
    endcase

    case (PM_CSR_BPCCEN)
      "FALSE" : PM_CSR_BPCCEN_BINARY = 1'b0;
      "TRUE" : PM_CSR_BPCCEN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CSR_BPCCEN on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_CSR_BPCCEN);
        #1 $finish;
      end
    endcase

    case (PM_CSR_NOSOFTRST)
      "TRUE" : PM_CSR_NOSOFTRST_BINARY = 1'b1;
      "FALSE" : PM_CSR_NOSOFTRST_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_CSR_NOSOFTRST on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_CSR_NOSOFTRST);
        #1 $finish;
      end
    endcase

    case (PM_MF)
      "FALSE" : PM_MF_BINARY = 1'b0;
      "TRUE" : PM_MF_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_MF on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PM_MF);
        #1 $finish;
      end
    endcase

    case (RBAR_CAP_ON)
      "FALSE" : RBAR_CAP_ON_BINARY = 1'b0;
      "TRUE" : RBAR_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RBAR_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", RBAR_CAP_ON);
        #1 $finish;
      end
    endcase

    case (RECRC_CHK_TRIM)
      "FALSE" : RECRC_CHK_TRIM_BINARY = 1'b0;
      "TRUE" : RECRC_CHK_TRIM_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute RECRC_CHK_TRIM on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", RECRC_CHK_TRIM);
        #1 $finish;
      end
    endcase

    case (ROOT_CAP_CRS_SW_VISIBILITY)
      "FALSE" : ROOT_CAP_CRS_SW_VISIBILITY_BINARY = 1'b0;
      "TRUE" : ROOT_CAP_CRS_SW_VISIBILITY_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ROOT_CAP_CRS_SW_VISIBILITY on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ROOT_CAP_CRS_SW_VISIBILITY);
        #1 $finish;
      end
    endcase

    case (SELECT_DLL_IF)
      "FALSE" : SELECT_DLL_IF_BINARY = 1'b0;
      "TRUE" : SELECT_DLL_IF_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SELECT_DLL_IF on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SELECT_DLL_IF);
        #1 $finish;
      end
    endcase

    case (SIM_VERSION)
      "1.0" : SIM_VERSION_BINARY = 0;
      "1.1" : SIM_VERSION_BINARY = 0;
      "1.2" : SIM_VERSION_BINARY = 0;
      "1.3" : SIM_VERSION_BINARY = 0;
      "2.0" : SIM_VERSION_BINARY = 0;
      "3.0" : SIM_VERSION_BINARY = 0;
      "4.0" : SIM_VERSION_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_VERSION on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are 1.0, 1.1, 1.2, 1.3, 2.0, 3.0, or 4.0.", SIM_VERSION);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_ATT_BUTTON_PRESENT)
      "FALSE" : SLOT_CAP_ATT_BUTTON_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_ATT_BUTTON_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_ATT_BUTTON_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_ATT_BUTTON_PRESENT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_ATT_INDICATOR_PRESENT)
      "FALSE" : SLOT_CAP_ATT_INDICATOR_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_ATT_INDICATOR_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_ATT_INDICATOR_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_ATT_INDICATOR_PRESENT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_ELEC_INTERLOCK_PRESENT)
      "FALSE" : SLOT_CAP_ELEC_INTERLOCK_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_ELEC_INTERLOCK_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_ELEC_INTERLOCK_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_ELEC_INTERLOCK_PRESENT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_HOTPLUG_CAPABLE)
      "FALSE" : SLOT_CAP_HOTPLUG_CAPABLE_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_HOTPLUG_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_HOTPLUG_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_HOTPLUG_CAPABLE);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_HOTPLUG_SURPRISE)
      "FALSE" : SLOT_CAP_HOTPLUG_SURPRISE_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_HOTPLUG_SURPRISE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_HOTPLUG_SURPRISE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_HOTPLUG_SURPRISE);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_MRL_SENSOR_PRESENT)
      "FALSE" : SLOT_CAP_MRL_SENSOR_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_MRL_SENSOR_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_MRL_SENSOR_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_MRL_SENSOR_PRESENT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_NO_CMD_COMPLETED_SUPPORT)
      "FALSE" : SLOT_CAP_NO_CMD_COMPLETED_SUPPORT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_NO_CMD_COMPLETED_SUPPORT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_NO_CMD_COMPLETED_SUPPORT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_NO_CMD_COMPLETED_SUPPORT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_POWER_CONTROLLER_PRESENT)
      "FALSE" : SLOT_CAP_POWER_CONTROLLER_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_POWER_CONTROLLER_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_POWER_CONTROLLER_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_POWER_CONTROLLER_PRESENT);
        #1 $finish;
      end
    endcase

    case (SLOT_CAP_POWER_INDICATOR_PRESENT)
      "FALSE" : SLOT_CAP_POWER_INDICATOR_PRESENT_BINARY = 1'b0;
      "TRUE" : SLOT_CAP_POWER_INDICATOR_PRESENT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SLOT_CAP_POWER_INDICATOR_PRESENT on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SLOT_CAP_POWER_INDICATOR_PRESENT);
        #1 $finish;
      end
    endcase

    case (SSL_MESSAGE_AUTO)
      "FALSE" : SSL_MESSAGE_AUTO_BINARY = 1'b0;
      "TRUE" : SSL_MESSAGE_AUTO_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SSL_MESSAGE_AUTO on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SSL_MESSAGE_AUTO);
        #1 $finish;
      end
    endcase

    case (TECRC_EP_INV)
      "FALSE" : TECRC_EP_INV_BINARY = 1'b0;
      "TRUE" : TECRC_EP_INV_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TECRC_EP_INV on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TECRC_EP_INV);
        #1 $finish;
      end
    endcase

    case (TL_RBYPASS)
      "FALSE" : TL_RBYPASS_BINARY = 1'b0;
      "TRUE" : TL_RBYPASS_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_RBYPASS on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_RBYPASS);
        #1 $finish;
      end
    endcase

    case (TL_TFC_DISABLE)
      "FALSE" : TL_TFC_DISABLE_BINARY = 1'b0;
      "TRUE" : TL_TFC_DISABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_TFC_DISABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_TFC_DISABLE);
        #1 $finish;
      end
    endcase

    case (TL_TX_CHECKS_DISABLE)
      "FALSE" : TL_TX_CHECKS_DISABLE_BINARY = 1'b0;
      "TRUE" : TL_TX_CHECKS_DISABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_TX_CHECKS_DISABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_TX_CHECKS_DISABLE);
        #1 $finish;
      end
    endcase

    case (TRN_DW)
      "FALSE" : TRN_DW_BINARY = 1'b0;
      "TRUE" : TRN_DW_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TRN_DW on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TRN_DW);
        #1 $finish;
      end
    endcase

    case (TRN_NP_FC)
      "FALSE" : TRN_NP_FC_BINARY = 1'b0;
      "TRUE" : TRN_NP_FC_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TRN_NP_FC on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TRN_NP_FC);
        #1 $finish;
      end
    endcase

    case (UPCONFIG_CAPABLE)
      "TRUE" : UPCONFIG_CAPABLE_BINARY = 1'b1;
      "FALSE" : UPCONFIG_CAPABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UPCONFIG_CAPABLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UPCONFIG_CAPABLE);
        #1 $finish;
      end
    endcase

    case (UPSTREAM_FACING)
      "TRUE" : UPSTREAM_FACING_BINARY = 1'b1;
      "FALSE" : UPSTREAM_FACING_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UPSTREAM_FACING on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UPSTREAM_FACING);
        #1 $finish;
      end
    endcase

    case (UR_ATOMIC)
      "TRUE" : UR_ATOMIC_BINARY = 1'b1;
      "FALSE" : UR_ATOMIC_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UR_ATOMIC on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UR_ATOMIC);
        #1 $finish;
      end
    endcase

    case (UR_CFG1)
      "TRUE" : UR_CFG1_BINARY = 1'b1;
      "FALSE" : UR_CFG1_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UR_CFG1 on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UR_CFG1);
        #1 $finish;
      end
    endcase

    case (UR_INV_REQ)
      "TRUE" : UR_INV_REQ_BINARY = 1'b1;
      "FALSE" : UR_INV_REQ_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UR_INV_REQ on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UR_INV_REQ);
        #1 $finish;
      end
    endcase

    case (UR_PRS_RESPONSE)
      "TRUE" : UR_PRS_RESPONSE_BINARY = 1'b1;
      "FALSE" : UR_PRS_RESPONSE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute UR_PRS_RESPONSE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", UR_PRS_RESPONSE);
        #1 $finish;
      end
    endcase

    case (USER_CLK2_DIV2)
      "FALSE" : USER_CLK2_DIV2_BINARY = 1'b0;
      "TRUE" : USER_CLK2_DIV2_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute USER_CLK2_DIV2 on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", USER_CLK2_DIV2);
        #1 $finish;
      end
    endcase

    case (USE_RID_PINS)
      "FALSE" : USE_RID_PINS_BINARY = 1'b0;
      "TRUE" : USE_RID_PINS_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute USE_RID_PINS on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", USE_RID_PINS);
        #1 $finish;
      end
    endcase

    case (VC0_CPL_INFINITE)
      "TRUE" : VC0_CPL_INFINITE_BINARY = 1'b1;
      "FALSE" : VC0_CPL_INFINITE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VC0_CPL_INFINITE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VC0_CPL_INFINITE);
        #1 $finish;
      end
    endcase

    case (VC_CAP_ON)
      "FALSE" : VC_CAP_ON_BINARY = 1'b0;
      "TRUE" : VC_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VC_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VC_CAP_ON);
        #1 $finish;
      end
    endcase

    case (VC_CAP_REJECT_SNOOP_TRANSACTIONS)
      "FALSE" : VC_CAP_REJECT_SNOOP_TRANSACTIONS_BINARY = 1'b0;
      "TRUE" : VC_CAP_REJECT_SNOOP_TRANSACTIONS_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VC_CAP_REJECT_SNOOP_TRANSACTIONS on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VC_CAP_REJECT_SNOOP_TRANSACTIONS);
        #1 $finish;
      end
    endcase

    case (VSEC_CAP_IS_LINK_VISIBLE)
      "TRUE" : VSEC_CAP_IS_LINK_VISIBLE_BINARY = 1'b1;
      "FALSE" : VSEC_CAP_IS_LINK_VISIBLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VSEC_CAP_IS_LINK_VISIBLE on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VSEC_CAP_IS_LINK_VISIBLE);
        #1 $finish;
      end
    endcase

    case (VSEC_CAP_ON)
      "FALSE" : VSEC_CAP_ON_BINARY = 1'b0;
      "TRUE" : VSEC_CAP_ON_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VSEC_CAP_ON on X_PCIE_2_1 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VSEC_CAP_ON);
        #1 $finish;
      end
    endcase

    if ((CFG_ECRC_ERR_CPLSTAT >= 0) && (CFG_ECRC_ERR_CPLSTAT <= 3))
      CFG_ECRC_ERR_CPLSTAT_BINARY = CFG_ECRC_ERR_CPLSTAT;
    else begin
      $display("Attribute Syntax Error : The Attribute CFG_ECRC_ERR_CPLSTAT on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", CFG_ECRC_ERR_CPLSTAT);
      #1 $finish;
    end

    if ((DEV_CAP_ENDPOINT_L0S_LATENCY >= 0) && (DEV_CAP_ENDPOINT_L0S_LATENCY <= 7))
      DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY = DEV_CAP_ENDPOINT_L0S_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_ENDPOINT_L0S_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", DEV_CAP_ENDPOINT_L0S_LATENCY);
      #1 $finish;
    end

    if ((DEV_CAP_ENDPOINT_L1_LATENCY >= 0) && (DEV_CAP_ENDPOINT_L1_LATENCY <= 7))
      DEV_CAP_ENDPOINT_L1_LATENCY_BINARY = DEV_CAP_ENDPOINT_L1_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_ENDPOINT_L1_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", DEV_CAP_ENDPOINT_L1_LATENCY);
      #1 $finish;
    end

    if ((DEV_CAP_MAX_PAYLOAD_SUPPORTED >= 0) && (DEV_CAP_MAX_PAYLOAD_SUPPORTED <= 7))
      DEV_CAP_MAX_PAYLOAD_SUPPORTED_BINARY = DEV_CAP_MAX_PAYLOAD_SUPPORTED;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_MAX_PAYLOAD_SUPPORTED on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", DEV_CAP_MAX_PAYLOAD_SUPPORTED);
      #1 $finish;
    end

    if ((DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT >= 0) && (DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT <= 3))
      DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT_BINARY = DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT);
      #1 $finish;
    end

    if ((DEV_CAP_RSVD_14_12 >= 0) && (DEV_CAP_RSVD_14_12 <= 7))
      DEV_CAP_RSVD_14_12_BINARY = DEV_CAP_RSVD_14_12;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_RSVD_14_12 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", DEV_CAP_RSVD_14_12);
      #1 $finish;
    end

    if ((DEV_CAP_RSVD_17_16 >= 0) && (DEV_CAP_RSVD_17_16 <= 3))
      DEV_CAP_RSVD_17_16_BINARY = DEV_CAP_RSVD_17_16;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_RSVD_17_16 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", DEV_CAP_RSVD_17_16);
      #1 $finish;
    end

    if ((DEV_CAP_RSVD_31_29 >= 0) && (DEV_CAP_RSVD_31_29 <= 7))
      DEV_CAP_RSVD_31_29_BINARY = DEV_CAP_RSVD_31_29;
    else begin
      $display("Attribute Syntax Error : The Attribute DEV_CAP_RSVD_31_29 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", DEV_CAP_RSVD_31_29);
      #1 $finish;
    end

    if ((LINK_CAP_ASPM_SUPPORT >= 0) && (LINK_CAP_ASPM_SUPPORT <= 3))
      LINK_CAP_ASPM_SUPPORT_BINARY = LINK_CAP_ASPM_SUPPORT;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_ASPM_SUPPORT on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LINK_CAP_ASPM_SUPPORT);
      #1 $finish;
    end

    if ((LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY = LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1);
      #1 $finish;
    end

    if ((LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY = LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2);
      #1 $finish;
    end

    if ((LINK_CAP_L0S_EXIT_LATENCY_GEN1 >= 0) && (LINK_CAP_L0S_EXIT_LATENCY_GEN1 <= 7))
      LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY = LINK_CAP_L0S_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L0S_EXIT_LATENCY_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L0S_EXIT_LATENCY_GEN1);
      #1 $finish;
    end

    if ((LINK_CAP_L0S_EXIT_LATENCY_GEN2 >= 0) && (LINK_CAP_L0S_EXIT_LATENCY_GEN2 <= 7))
      LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY = LINK_CAP_L0S_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L0S_EXIT_LATENCY_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L0S_EXIT_LATENCY_GEN2);
      #1 $finish;
    end

    if ((LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY = LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1);
      #1 $finish;
    end

    if ((LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY = LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2);
      #1 $finish;
    end

    if ((LINK_CAP_L1_EXIT_LATENCY_GEN1 >= 0) && (LINK_CAP_L1_EXIT_LATENCY_GEN1 <= 7))
      LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY = LINK_CAP_L1_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L1_EXIT_LATENCY_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L1_EXIT_LATENCY_GEN1);
      #1 $finish;
    end

    if ((LINK_CAP_L1_EXIT_LATENCY_GEN2 >= 0) && (LINK_CAP_L1_EXIT_LATENCY_GEN2 <= 7))
      LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY = LINK_CAP_L1_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_L1_EXIT_LATENCY_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", LINK_CAP_L1_EXIT_LATENCY_GEN2);
      #1 $finish;
    end

    if ((LINK_CAP_RSVD_23 >= 0) && (LINK_CAP_RSVD_23 <= 1))
      LINK_CAP_RSVD_23_BINARY = LINK_CAP_RSVD_23;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CAP_RSVD_23 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", LINK_CAP_RSVD_23);
      #1 $finish;
    end

    if ((LINK_CONTROL_RCB >= 0) && (LINK_CONTROL_RCB <= 1))
      LINK_CONTROL_RCB_BINARY = LINK_CONTROL_RCB;
    else begin
      $display("Attribute Syntax Error : The Attribute LINK_CONTROL_RCB on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", LINK_CONTROL_RCB);
      #1 $finish;
    end

    if ((LL_ACK_TIMEOUT_FUNC >= 0) && (LL_ACK_TIMEOUT_FUNC <= 3))
      LL_ACK_TIMEOUT_FUNC_BINARY = LL_ACK_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_FUNC on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_ACK_TIMEOUT_FUNC);
      #1 $finish;
    end

    if ((LL_REPLAY_TIMEOUT_FUNC >= 0) && (LL_REPLAY_TIMEOUT_FUNC <= 3))
      LL_REPLAY_TIMEOUT_FUNC_BINARY = LL_REPLAY_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_FUNC on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_REPLAY_TIMEOUT_FUNC);
      #1 $finish;
    end

    if ((MSIX_CAP_PBA_BIR >= 0) && (MSIX_CAP_PBA_BIR <= 7))
      MSIX_CAP_PBA_BIR_BINARY = MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute MSIX_CAP_PBA_BIR on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", MSIX_CAP_PBA_BIR);
      #1 $finish;
    end

    if ((MSIX_CAP_TABLE_BIR >= 0) && (MSIX_CAP_TABLE_BIR <= 7))
      MSIX_CAP_TABLE_BIR_BINARY = MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute MSIX_CAP_TABLE_BIR on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", MSIX_CAP_TABLE_BIR);
      #1 $finish;
    end

    if ((MSI_CAP_MULTIMSGCAP >= 0) && (MSI_CAP_MULTIMSGCAP <= 7))
      MSI_CAP_MULTIMSGCAP_BINARY = MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute MSI_CAP_MULTIMSGCAP on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", MSI_CAP_MULTIMSGCAP);
      #1 $finish;
    end

    if ((MSI_CAP_MULTIMSG_EXTENSION >= 0) && (MSI_CAP_MULTIMSG_EXTENSION <= 1))
      MSI_CAP_MULTIMSG_EXTENSION_BINARY = MSI_CAP_MULTIMSG_EXTENSION;
    else begin
      $display("Attribute Syntax Error : The Attribute MSI_CAP_MULTIMSG_EXTENSION on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", MSI_CAP_MULTIMSG_EXTENSION);
      #1 $finish;
    end

    if ((N_FTS_COMCLK_GEN1 >= 0) && (N_FTS_COMCLK_GEN1 <= 255))
      N_FTS_COMCLK_GEN1_BINARY = N_FTS_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute N_FTS_COMCLK_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", N_FTS_COMCLK_GEN1);
      #1 $finish;
    end

    if ((N_FTS_COMCLK_GEN2 >= 0) && (N_FTS_COMCLK_GEN2 <= 255))
      N_FTS_COMCLK_GEN2_BINARY = N_FTS_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute N_FTS_COMCLK_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", N_FTS_COMCLK_GEN2);
      #1 $finish;
    end

    if ((N_FTS_GEN1 >= 0) && (N_FTS_GEN1 <= 255))
      N_FTS_GEN1_BINARY = N_FTS_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute N_FTS_GEN1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", N_FTS_GEN1);
      #1 $finish;
    end

    if ((N_FTS_GEN2 >= 0) && (N_FTS_GEN2 <= 255))
      N_FTS_GEN2_BINARY = N_FTS_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute N_FTS_GEN2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", N_FTS_GEN2);
      #1 $finish;
    end

    if ((PCIE_CAP_RSVD_15_14 >= 0) && (PCIE_CAP_RSVD_15_14 <= 3))
      PCIE_CAP_RSVD_15_14_BINARY = PCIE_CAP_RSVD_15_14;
    else begin
      $display("Attribute Syntax Error : The Attribute PCIE_CAP_RSVD_15_14 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", PCIE_CAP_RSVD_15_14);
      #1 $finish;
    end

    if ((PCIE_REVISION >= 0) && (PCIE_REVISION <= 15))
      PCIE_REVISION_BINARY = PCIE_REVISION;
    else begin
      $display("Attribute Syntax Error : The Attribute PCIE_REVISION on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 15.", PCIE_REVISION);
      #1 $finish;
    end

    if ((PL_AUTO_CONFIG >= 0) && (PL_AUTO_CONFIG <= 7))
      PL_AUTO_CONFIG_BINARY = PL_AUTO_CONFIG;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_AUTO_CONFIG on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PL_AUTO_CONFIG);
      #1 $finish;
    end

    if ((PM_ASPML0S_TIMEOUT_FUNC >= 0) && (PM_ASPML0S_TIMEOUT_FUNC <= 3))
      PM_ASPML0S_TIMEOUT_FUNC_BINARY = PM_ASPML0S_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute PM_ASPML0S_TIMEOUT_FUNC on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", PM_ASPML0S_TIMEOUT_FUNC);
      #1 $finish;
    end

    if ((PM_CAP_AUXCURRENT >= 0) && (PM_CAP_AUXCURRENT <= 7))
      PM_CAP_AUXCURRENT_BINARY = PM_CAP_AUXCURRENT;
    else begin
      $display("Attribute Syntax Error : The Attribute PM_CAP_AUXCURRENT on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PM_CAP_AUXCURRENT);
      #1 $finish;
    end

    if ((PM_CAP_RSVD_04 >= 0) && (PM_CAP_RSVD_04 <= 1))
      PM_CAP_RSVD_04_BINARY = PM_CAP_RSVD_04;
    else begin
      $display("Attribute Syntax Error : The Attribute PM_CAP_RSVD_04 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", PM_CAP_RSVD_04);
      #1 $finish;
    end

    if ((PM_CAP_VERSION >= 0) && (PM_CAP_VERSION <= 7))
      PM_CAP_VERSION_BINARY = PM_CAP_VERSION;
    else begin
      $display("Attribute Syntax Error : The Attribute PM_CAP_VERSION on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PM_CAP_VERSION);
      #1 $finish;
    end

    if ((RECRC_CHK >= 0) && (RECRC_CHK <= 3))
      RECRC_CHK_BINARY = RECRC_CHK;
    else begin
      $display("Attribute Syntax Error : The Attribute RECRC_CHK on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", RECRC_CHK);
      #1 $finish;
    end

    if ((SLOT_CAP_SLOT_POWER_LIMIT_SCALE >= 0) && (SLOT_CAP_SLOT_POWER_LIMIT_SCALE <= 3))
      SLOT_CAP_SLOT_POWER_LIMIT_SCALE_BINARY = SLOT_CAP_SLOT_POWER_LIMIT_SCALE;
    else begin
      $display("Attribute Syntax Error : The Attribute SLOT_CAP_SLOT_POWER_LIMIT_SCALE on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", SLOT_CAP_SLOT_POWER_LIMIT_SCALE);
      #1 $finish;
    end

    if ((SPARE_BIT0 >= 0) && (SPARE_BIT0 <= 1))
      SPARE_BIT0_BINARY = SPARE_BIT0;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT0 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT0);
      #1 $finish;
    end

    if ((SPARE_BIT1 >= 0) && (SPARE_BIT1 <= 1))
      SPARE_BIT1_BINARY = SPARE_BIT1;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT1 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT1);
      #1 $finish;
    end

    if ((SPARE_BIT2 >= 0) && (SPARE_BIT2 <= 1))
      SPARE_BIT2_BINARY = SPARE_BIT2;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT2 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT2);
      #1 $finish;
    end

    if ((SPARE_BIT3 >= 0) && (SPARE_BIT3 <= 1))
      SPARE_BIT3_BINARY = SPARE_BIT3;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT3 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT3);
      #1 $finish;
    end

    if ((SPARE_BIT4 >= 0) && (SPARE_BIT4 <= 1))
      SPARE_BIT4_BINARY = SPARE_BIT4;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT4 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT4);
      #1 $finish;
    end

    if ((SPARE_BIT5 >= 0) && (SPARE_BIT5 <= 1))
      SPARE_BIT5_BINARY = SPARE_BIT5;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT5 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT5);
      #1 $finish;
    end

    if ((SPARE_BIT6 >= 0) && (SPARE_BIT6 <= 1))
      SPARE_BIT6_BINARY = SPARE_BIT6;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT6 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT6);
      #1 $finish;
    end

    if ((SPARE_BIT7 >= 0) && (SPARE_BIT7 <= 1))
      SPARE_BIT7_BINARY = SPARE_BIT7;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT7 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT7);
      #1 $finish;
    end

    if ((SPARE_BIT8 >= 0) && (SPARE_BIT8 <= 1))
      SPARE_BIT8_BINARY = SPARE_BIT8;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT8 on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT8);
      #1 $finish;
    end

    if ((TL_RX_RAM_RADDR_LATENCY >= 0) && (TL_RX_RAM_RADDR_LATENCY <= 1))
      TL_RX_RAM_RADDR_LATENCY_BINARY = TL_RX_RAM_RADDR_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_RX_RAM_RADDR_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", TL_RX_RAM_RADDR_LATENCY);
      #1 $finish;
    end

    if ((TL_RX_RAM_RDATA_LATENCY >= 0) && (TL_RX_RAM_RDATA_LATENCY <= 3))
      TL_RX_RAM_RDATA_LATENCY_BINARY = TL_RX_RAM_RDATA_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_RX_RAM_RDATA_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", TL_RX_RAM_RDATA_LATENCY);
      #1 $finish;
    end

    if ((TL_RX_RAM_WRITE_LATENCY >= 0) && (TL_RX_RAM_WRITE_LATENCY <= 1))
      TL_RX_RAM_WRITE_LATENCY_BINARY = TL_RX_RAM_WRITE_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_RX_RAM_WRITE_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", TL_RX_RAM_WRITE_LATENCY);
      #1 $finish;
    end

    if ((TL_TX_RAM_RADDR_LATENCY >= 0) && (TL_TX_RAM_RADDR_LATENCY <= 1))
      TL_TX_RAM_RADDR_LATENCY_BINARY = TL_TX_RAM_RADDR_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_TX_RAM_RADDR_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", TL_TX_RAM_RADDR_LATENCY);
      #1 $finish;
    end

    if ((TL_TX_RAM_RDATA_LATENCY >= 0) && (TL_TX_RAM_RDATA_LATENCY <= 3))
      TL_TX_RAM_RDATA_LATENCY_BINARY = TL_TX_RAM_RDATA_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_TX_RAM_RDATA_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", TL_TX_RAM_RDATA_LATENCY);
      #1 $finish;
    end

    if ((TL_TX_RAM_WRITE_LATENCY >= 0) && (TL_TX_RAM_WRITE_LATENCY <= 1))
      TL_TX_RAM_WRITE_LATENCY_BINARY = TL_TX_RAM_WRITE_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute TL_TX_RAM_WRITE_LATENCY on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", TL_TX_RAM_WRITE_LATENCY);
      #1 $finish;
    end

    if ((USER_CLK_FREQ >= 0) && (USER_CLK_FREQ <= 7))
      USER_CLK_FREQ_BINARY = USER_CLK_FREQ;
    else begin
      $display("Attribute Syntax Error : The Attribute USER_CLK_FREQ on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", USER_CLK_FREQ);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_CD >= 0) && (VC0_TOTAL_CREDITS_CD <= 2047))
      VC0_TOTAL_CREDITS_CD_BINARY = VC0_TOTAL_CREDITS_CD;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_CD on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 2047.", VC0_TOTAL_CREDITS_CD);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_CH >= 0) && (VC0_TOTAL_CREDITS_CH <= 127))
      VC0_TOTAL_CREDITS_CH_BINARY = VC0_TOTAL_CREDITS_CH;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_CH on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 127.", VC0_TOTAL_CREDITS_CH);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_NPD >= 0) && (VC0_TOTAL_CREDITS_NPD <= 2047))
      VC0_TOTAL_CREDITS_NPD_BINARY = VC0_TOTAL_CREDITS_NPD;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_NPD on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 2047.", VC0_TOTAL_CREDITS_NPD);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_NPH >= 0) && (VC0_TOTAL_CREDITS_NPH <= 127))
      VC0_TOTAL_CREDITS_NPH_BINARY = VC0_TOTAL_CREDITS_NPH;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_NPH on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 127.", VC0_TOTAL_CREDITS_NPH);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_PD >= 0) && (VC0_TOTAL_CREDITS_PD <= 2047))
      VC0_TOTAL_CREDITS_PD_BINARY = VC0_TOTAL_CREDITS_PD;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_PD on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 2047.", VC0_TOTAL_CREDITS_PD);
      #1 $finish;
    end

    if ((VC0_TOTAL_CREDITS_PH >= 0) && (VC0_TOTAL_CREDITS_PH <= 127))
      VC0_TOTAL_CREDITS_PH_BINARY = VC0_TOTAL_CREDITS_PH;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TOTAL_CREDITS_PH on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 127.", VC0_TOTAL_CREDITS_PH);
      #1 $finish;
    end

    if ((VC0_TX_LASTPACKET >= 0) && (VC0_TX_LASTPACKET <= 31))
      VC0_TX_LASTPACKET_BINARY = VC0_TX_LASTPACKET;
    else begin
      $display("Attribute Syntax Error : The Attribute VC0_TX_LASTPACKET on X_PCIE_2_1 instance %m is set to %d.  Legal values for this attribute are  0 to 31.", VC0_TX_LASTPACKET);
      #1 $finish;
    end

  end

  wire [11:0] delay_DBGVECC;
  wire [11:0] delay_PLDBGVEC;
  wire [11:0] delay_TRNFCCPLD;
  wire [11:0] delay_TRNFCNPD;
  wire [11:0] delay_TRNFCPD;
  wire [127:0] delay_TRNRD;
  wire [12:0] delay_MIMRXRADDR;
  wire [12:0] delay_MIMRXWADDR;
  wire [12:0] delay_MIMTXRADDR;
  wire [12:0] delay_MIMTXWADDR;
  wire [15:0] delay_CFGMSGDATA;
  wire [15:0] delay_DRPDO;
  wire [15:0] delay_PIPETX0DATA;
  wire [15:0] delay_PIPETX1DATA;
  wire [15:0] delay_PIPETX2DATA;
  wire [15:0] delay_PIPETX3DATA;
  wire [15:0] delay_PIPETX4DATA;
  wire [15:0] delay_PIPETX5DATA;
  wire [15:0] delay_PIPETX6DATA;
  wire [15:0] delay_PIPETX7DATA;
  wire [1:0] delay_CFGLINKCONTROLASPMCONTROL;
  wire [1:0] delay_CFGLINKSTATUSCURRENTSPEED;
  wire [1:0] delay_CFGPMCSRPOWERSTATE;
  wire [1:0] delay_PIPETX0CHARISK;
  wire [1:0] delay_PIPETX0POWERDOWN;
  wire [1:0] delay_PIPETX1CHARISK;
  wire [1:0] delay_PIPETX1POWERDOWN;
  wire [1:0] delay_PIPETX2CHARISK;
  wire [1:0] delay_PIPETX2POWERDOWN;
  wire [1:0] delay_PIPETX3CHARISK;
  wire [1:0] delay_PIPETX3POWERDOWN;
  wire [1:0] delay_PIPETX4CHARISK;
  wire [1:0] delay_PIPETX4POWERDOWN;
  wire [1:0] delay_PIPETX5CHARISK;
  wire [1:0] delay_PIPETX5POWERDOWN;
  wire [1:0] delay_PIPETX6CHARISK;
  wire [1:0] delay_PIPETX6POWERDOWN;
  wire [1:0] delay_PIPETX7CHARISK;
  wire [1:0] delay_PIPETX7POWERDOWN;
  wire [1:0] delay_PL2RXPMSTATE;
  wire [1:0] delay_PLLANEREVERSALMODE;
  wire [1:0] delay_PLRXPMSTATE;
  wire [1:0] delay_PLSELLNKWIDTH;
  wire [1:0] delay_TRNRDLLPSRCRDY;
  wire [1:0] delay_TRNRREM;
  wire [2:0] delay_CFGDEVCONTROLMAXPAYLOAD;
  wire [2:0] delay_CFGDEVCONTROLMAXREADREQ;
  wire [2:0] delay_CFGINTERRUPTMMENABLE;
  wire [2:0] delay_CFGPCIELINKSTATE;
  wire [2:0] delay_PIPETXMARGIN;
  wire [2:0] delay_PLINITIALLINKWIDTH;
  wire [2:0] delay_PLTXPMSTATE;
  wire [31:0] delay_CFGMGMTDO;
  wire [3:0] delay_CFGDEVCONTROL2CPLTIMEOUTVAL;
  wire [3:0] delay_CFGLINKSTATUSNEGOTIATEDWIDTH;
  wire [3:0] delay_TRNTDSTRDY;
  wire [4:0] delay_LL2LINKSTATUS;
  wire [5:0] delay_PLLTSSMSTATE;
  wire [5:0] delay_TRNTBUFAV;
  wire [63:0] delay_DBGVECA;
  wire [63:0] delay_DBGVECB;
  wire [63:0] delay_TL2ERRHDR;
  wire [63:0] delay_TRNRDLLPDATA;
  wire [67:0] delay_MIMRXWDATA;
  wire [68:0] delay_MIMTXWDATA;
  wire [6:0] delay_CFGTRANSACTIONADDR;
  wire [6:0] delay_CFGVCTCVCMAP;
  wire [7:0] delay_CFGINTERRUPTDO;
  wire [7:0] delay_TRNFCCPLH;
  wire [7:0] delay_TRNFCNPH;
  wire [7:0] delay_TRNFCPH;
  wire [7:0] delay_TRNRBARHIT;
  wire delay_CFGAERECRCCHECKEN;
  wire delay_CFGAERECRCGENEN;
  wire delay_CFGAERROOTERRCORRERRRECEIVED;
  wire delay_CFGAERROOTERRCORRERRREPORTINGEN;
  wire delay_CFGAERROOTERRFATALERRRECEIVED;
  wire delay_CFGAERROOTERRFATALERRREPORTINGEN;
  wire delay_CFGAERROOTERRNONFATALERRRECEIVED;
  wire delay_CFGAERROOTERRNONFATALERRREPORTINGEN;
  wire delay_CFGBRIDGESERREN;
  wire delay_CFGCOMMANDBUSMASTERENABLE;
  wire delay_CFGCOMMANDINTERRUPTDISABLE;
  wire delay_CFGCOMMANDIOENABLE;
  wire delay_CFGCOMMANDMEMENABLE;
  wire delay_CFGCOMMANDSERREN;
  wire delay_CFGDEVCONTROL2ARIFORWARDEN;
  wire delay_CFGDEVCONTROL2ATOMICEGRESSBLOCK;
  wire delay_CFGDEVCONTROL2ATOMICREQUESTEREN;
  wire delay_CFGDEVCONTROL2CPLTIMEOUTDIS;
  wire delay_CFGDEVCONTROL2IDOCPLEN;
  wire delay_CFGDEVCONTROL2IDOREQEN;
  wire delay_CFGDEVCONTROL2LTREN;
  wire delay_CFGDEVCONTROL2TLPPREFIXBLOCK;
  wire delay_CFGDEVCONTROLAUXPOWEREN;
  wire delay_CFGDEVCONTROLCORRERRREPORTINGEN;
  wire delay_CFGDEVCONTROLENABLERO;
  wire delay_CFGDEVCONTROLEXTTAGEN;
  wire delay_CFGDEVCONTROLFATALERRREPORTINGEN;
  wire delay_CFGDEVCONTROLNONFATALREPORTINGEN;
  wire delay_CFGDEVCONTROLNOSNOOPEN;
  wire delay_CFGDEVCONTROLPHANTOMEN;
  wire delay_CFGDEVCONTROLURERRREPORTINGEN;
  wire delay_CFGDEVSTATUSCORRERRDETECTED;
  wire delay_CFGDEVSTATUSFATALERRDETECTED;
  wire delay_CFGDEVSTATUSNONFATALERRDETECTED;
  wire delay_CFGDEVSTATUSURDETECTED;
  wire delay_CFGERRAERHEADERLOGSETN;
  wire delay_CFGERRCPLRDYN;
  wire delay_CFGINTERRUPTMSIENABLE;
  wire delay_CFGINTERRUPTMSIXENABLE;
  wire delay_CFGINTERRUPTMSIXFM;
  wire delay_CFGINTERRUPTRDYN;
  wire delay_CFGLINKCONTROLAUTOBANDWIDTHINTEN;
  wire delay_CFGLINKCONTROLBANDWIDTHINTEN;
  wire delay_CFGLINKCONTROLCLOCKPMEN;
  wire delay_CFGLINKCONTROLCOMMONCLOCK;
  wire delay_CFGLINKCONTROLEXTENDEDSYNC;
  wire delay_CFGLINKCONTROLHWAUTOWIDTHDIS;
  wire delay_CFGLINKCONTROLLINKDISABLE;
  wire delay_CFGLINKCONTROLRCB;
  wire delay_CFGLINKCONTROLRETRAINLINK;
  wire delay_CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
  wire delay_CFGLINKSTATUSBANDWIDTHSTATUS;
  wire delay_CFGLINKSTATUSDLLACTIVE;
  wire delay_CFGLINKSTATUSLINKTRAINING;
  wire delay_CFGMGMTRDWRDONEN;
  wire delay_CFGMSGRECEIVED;
  wire delay_CFGMSGRECEIVEDASSERTINTA;
  wire delay_CFGMSGRECEIVEDASSERTINTB;
  wire delay_CFGMSGRECEIVEDASSERTINTC;
  wire delay_CFGMSGRECEIVEDASSERTINTD;
  wire delay_CFGMSGRECEIVEDDEASSERTINTA;
  wire delay_CFGMSGRECEIVEDDEASSERTINTB;
  wire delay_CFGMSGRECEIVEDDEASSERTINTC;
  wire delay_CFGMSGRECEIVEDDEASSERTINTD;
  wire delay_CFGMSGRECEIVEDERRCOR;
  wire delay_CFGMSGRECEIVEDERRFATAL;
  wire delay_CFGMSGRECEIVEDERRNONFATAL;
  wire delay_CFGMSGRECEIVEDPMASNAK;
  wire delay_CFGMSGRECEIVEDPMETO;
  wire delay_CFGMSGRECEIVEDPMETOACK;
  wire delay_CFGMSGRECEIVEDPMPME;
  wire delay_CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
  wire delay_CFGMSGRECEIVEDUNLOCK;
  wire delay_CFGPMCSRPMEEN;
  wire delay_CFGPMCSRPMESTATUS;
  wire delay_CFGPMRCVASREQL1N;
  wire delay_CFGPMRCVENTERL1N;
  wire delay_CFGPMRCVENTERL23N;
  wire delay_CFGPMRCVREQACKN;
  wire delay_CFGROOTCONTROLPMEINTEN;
  wire delay_CFGROOTCONTROLSYSERRCORRERREN;
  wire delay_CFGROOTCONTROLSYSERRFATALERREN;
  wire delay_CFGROOTCONTROLSYSERRNONFATALERREN;
  wire delay_CFGSLOTCONTROLELECTROMECHILCTLPULSE;
  wire delay_CFGTRANSACTION;
  wire delay_CFGTRANSACTIONTYPE;
  wire delay_DBGSCLRA;
  wire delay_DBGSCLRB;
  wire delay_DBGSCLRC;
  wire delay_DBGSCLRD;
  wire delay_DBGSCLRE;
  wire delay_DBGSCLRF;
  wire delay_DBGSCLRG;
  wire delay_DBGSCLRH;
  wire delay_DBGSCLRI;
  wire delay_DBGSCLRJ;
  wire delay_DBGSCLRK;
  wire delay_DRPRDY;
  wire delay_LL2BADDLLPERR;
  wire delay_LL2BADTLPERR;
  wire delay_LL2PROTOCOLERR;
  wire delay_LL2RECEIVERERR;
  wire delay_LL2REPLAYROERR;
  wire delay_LL2REPLAYTOERR;
  wire delay_LL2SUSPENDOK;
  wire delay_LL2TFCINIT1SEQ;
  wire delay_LL2TFCINIT2SEQ;
  wire delay_LL2TXIDLE;
  wire delay_LNKCLKEN;
  wire delay_MIMRXREN;
  wire delay_MIMRXWEN;
  wire delay_MIMTXREN;
  wire delay_MIMTXWEN;
  wire delay_PIPERX0POLARITY;
  wire delay_PIPERX1POLARITY;
  wire delay_PIPERX2POLARITY;
  wire delay_PIPERX3POLARITY;
  wire delay_PIPERX4POLARITY;
  wire delay_PIPERX5POLARITY;
  wire delay_PIPERX6POLARITY;
  wire delay_PIPERX7POLARITY;
  wire delay_PIPETX0COMPLIANCE;
  wire delay_PIPETX0ELECIDLE;
  wire delay_PIPETX1COMPLIANCE;
  wire delay_PIPETX1ELECIDLE;
  wire delay_PIPETX2COMPLIANCE;
  wire delay_PIPETX2ELECIDLE;
  wire delay_PIPETX3COMPLIANCE;
  wire delay_PIPETX3ELECIDLE;
  wire delay_PIPETX4COMPLIANCE;
  wire delay_PIPETX4ELECIDLE;
  wire delay_PIPETX5COMPLIANCE;
  wire delay_PIPETX5ELECIDLE;
  wire delay_PIPETX6COMPLIANCE;
  wire delay_PIPETX6ELECIDLE;
  wire delay_PIPETX7COMPLIANCE;
  wire delay_PIPETX7ELECIDLE;
  wire delay_PIPETXDEEMPH;
  wire delay_PIPETXRATE;
  wire delay_PIPETXRCVRDET;
  wire delay_PIPETXRESET;
  wire delay_PL2L0REQ;
  wire delay_PL2LINKUP;
  wire delay_PL2RECEIVERERR;
  wire delay_PL2RECOVERY;
  wire delay_PL2RXELECIDLE;
  wire delay_PL2SUSPENDOK;
  wire delay_PLDIRECTEDCHANGEDONE;
  wire delay_PLLINKGEN2CAP;
  wire delay_PLLINKPARTNERGEN2SUPPORTED;
  wire delay_PLLINKUPCFGCAP;
  wire delay_PLPHYLNKUPN;
  wire delay_PLRECEIVEDHOTRST;
  wire delay_PLSELLNKRATE;
  wire delay_RECEIVEDFUNCLVLRSTN;
  wire delay_TL2ASPMSUSPENDCREDITCHECKOK;
  wire delay_TL2ASPMSUSPENDREQ;
  wire delay_TL2ERRFCPE;
  wire delay_TL2ERRMALFORMED;
  wire delay_TL2ERRRXOVERFLOW;
  wire delay_TL2PPMSUSPENDOK;
  wire delay_TRNLNKUP;
  wire delay_TRNRECRCERR;
  wire delay_TRNREOF;
  wire delay_TRNRERRFWD;
  wire delay_TRNRSOF;
  wire delay_TRNRSRCDSC;
  wire delay_TRNRSRCRDY;
  wire delay_TRNTCFGREQ;
  wire delay_TRNTDLLPDSTRDY;
  wire delay_TRNTERRDROP;
  wire delay_USERRSTN;

  wire [127:0] delay_CFGERRAERHEADERLOG;
  wire [127:0] delay_TRNTD;
  wire [15:0] delay_CFGDEVID;
  wire [15:0] delay_CFGSUBSYSID;
  wire [15:0] delay_CFGSUBSYSVENDID;
  wire [15:0] delay_CFGVENDID;
  wire [15:0] delay_DRPDI;
  wire [15:0] delay_PIPERX0DATA;
  wire [15:0] delay_PIPERX1DATA;
  wire [15:0] delay_PIPERX2DATA;
  wire [15:0] delay_PIPERX3DATA;
  wire [15:0] delay_PIPERX4DATA;
  wire [15:0] delay_PIPERX5DATA;
  wire [15:0] delay_PIPERX6DATA;
  wire [15:0] delay_PIPERX7DATA;
  wire [1:0] delay_CFGPMFORCESTATE;
  wire [1:0] delay_DBGMODE;
  wire [1:0] delay_PIPERX0CHARISK;
  wire [1:0] delay_PIPERX1CHARISK;
  wire [1:0] delay_PIPERX2CHARISK;
  wire [1:0] delay_PIPERX3CHARISK;
  wire [1:0] delay_PIPERX4CHARISK;
  wire [1:0] delay_PIPERX5CHARISK;
  wire [1:0] delay_PIPERX6CHARISK;
  wire [1:0] delay_PIPERX7CHARISK;
  wire [1:0] delay_PLDIRECTEDLINKCHANGE;
  wire [1:0] delay_PLDIRECTEDLINKWIDTH;
  wire [1:0] delay_TRNTREM;
  wire [2:0] delay_CFGDSFUNCTIONNUMBER;
  wire [2:0] delay_CFGFORCEMPS;
  wire [2:0] delay_PIPERX0STATUS;
  wire [2:0] delay_PIPERX1STATUS;
  wire [2:0] delay_PIPERX2STATUS;
  wire [2:0] delay_PIPERX3STATUS;
  wire [2:0] delay_PIPERX4STATUS;
  wire [2:0] delay_PIPERX5STATUS;
  wire [2:0] delay_PIPERX6STATUS;
  wire [2:0] delay_PIPERX7STATUS;
  wire [2:0] delay_PLDBGMODE;
  wire [2:0] delay_TRNFCSEL;
  wire [31:0] delay_CFGMGMTDI;
  wire [31:0] delay_TRNTDLLPDATA;
  wire [3:0] delay_CFGMGMTBYTEENN;
  wire [47:0] delay_CFGERRTLPCPLHEADER;
  wire [4:0] delay_CFGAERINTERRUPTMSGNUM;
  wire [4:0] delay_CFGDSDEVICENUMBER;
  wire [4:0] delay_CFGPCIECAPINTERRUPTMSGNUM;
  wire [4:0] delay_PL2DIRECTEDLSTATE;
  wire [5:0] delay_PLDIRECTEDLTSSMNEW;
  wire [63:0] delay_CFGDSN;
  wire [67:0] delay_MIMRXRDATA;
  wire [68:0] delay_MIMTXRDATA;
  wire [7:0] delay_CFGDSBUSNUMBER;
  wire [7:0] delay_CFGINTERRUPTDI;
  wire [7:0] delay_CFGPORTNUMBER;
  wire [7:0] delay_CFGREVID;
  wire [8:0] delay_DRPADDR;
  wire [9:0] delay_CFGMGMTDWADDR;
  wire delay_CFGERRACSN;
  wire delay_CFGERRATOMICEGRESSBLOCKEDN;
  wire delay_CFGERRCORN;
  wire delay_CFGERRCPLABORTN;
  wire delay_CFGERRCPLTIMEOUTN;
  wire delay_CFGERRCPLUNEXPECTN;
  wire delay_CFGERRECRCN;
  wire delay_CFGERRINTERNALCORN;
  wire delay_CFGERRINTERNALUNCORN;
  wire delay_CFGERRLOCKEDN;
  wire delay_CFGERRMALFORMEDN;
  wire delay_CFGERRMCBLOCKEDN;
  wire delay_CFGERRNORECOVERYN;
  wire delay_CFGERRPOISONEDN;
  wire delay_CFGERRPOSTEDN;
  wire delay_CFGERRURN;
  wire delay_CFGFORCECOMMONCLOCKOFF;
  wire delay_CFGFORCEEXTENDEDSYNCON;
  wire delay_CFGINTERRUPTASSERTN;
  wire delay_CFGINTERRUPTN;
  wire delay_CFGINTERRUPTSTATN;
  wire delay_CFGMGMTRDENN;
  wire delay_CFGMGMTWRENN;
  wire delay_CFGMGMTWRREADONLYN;
  wire delay_CFGMGMTWRRW1CASRWN;
  wire delay_CFGPMFORCESTATEENN;
  wire delay_CFGPMHALTASPML0SN;
  wire delay_CFGPMHALTASPML1N;
  wire delay_CFGPMSENDPMETON;
  wire delay_CFGPMTURNOFFOKN;
  wire delay_CFGPMWAKEN;
  wire delay_CFGTRNPENDINGN;
  wire delay_CMRSTN;
  wire delay_CMSTICKYRSTN;
  wire delay_DBGSUBMODE;
  wire delay_DLRSTN;
  wire delay_DRPCLK;
  wire delay_DRPEN;
  wire delay_DRPWE;
  wire delay_FUNCLVLRSTN;
  wire delay_LL2SENDASREQL1;
  wire delay_LL2SENDENTERL1;
  wire delay_LL2SENDENTERL23;
  wire delay_LL2SENDPMACK;
  wire delay_LL2SUSPENDNOW;
  wire delay_LL2TLPRCV;
  wire delay_PIPECLK;
  wire delay_PIPERX0CHANISALIGNED;
  wire delay_PIPERX0ELECIDLE;
  wire delay_PIPERX0PHYSTATUS;
  wire delay_PIPERX0VALID;
  wire delay_PIPERX1CHANISALIGNED;
  wire delay_PIPERX1ELECIDLE;
  wire delay_PIPERX1PHYSTATUS;
  wire delay_PIPERX1VALID;
  wire delay_PIPERX2CHANISALIGNED;
  wire delay_PIPERX2ELECIDLE;
  wire delay_PIPERX2PHYSTATUS;
  wire delay_PIPERX2VALID;
  wire delay_PIPERX3CHANISALIGNED;
  wire delay_PIPERX3ELECIDLE;
  wire delay_PIPERX3PHYSTATUS;
  wire delay_PIPERX3VALID;
  wire delay_PIPERX4CHANISALIGNED;
  wire delay_PIPERX4ELECIDLE;
  wire delay_PIPERX4PHYSTATUS;
  wire delay_PIPERX4VALID;
  wire delay_PIPERX5CHANISALIGNED;
  wire delay_PIPERX5ELECIDLE;
  wire delay_PIPERX5PHYSTATUS;
  wire delay_PIPERX5VALID;
  wire delay_PIPERX6CHANISALIGNED;
  wire delay_PIPERX6ELECIDLE;
  wire delay_PIPERX6PHYSTATUS;
  wire delay_PIPERX6VALID;
  wire delay_PIPERX7CHANISALIGNED;
  wire delay_PIPERX7ELECIDLE;
  wire delay_PIPERX7PHYSTATUS;
  wire delay_PIPERX7VALID;
  wire delay_PLDIRECTEDLINKAUTON;
  wire delay_PLDIRECTEDLINKSPEED;
  wire delay_PLDIRECTEDLTSSMNEWVLD;
  wire delay_PLDIRECTEDLTSSMSTALL;
  wire delay_PLDOWNSTREAMDEEMPHSOURCE;
  wire delay_PLRSTN;
  wire delay_PLTRANSMITHOTRST;
  wire delay_PLUPSTREAMPREFERDEEMPH;
  wire delay_SYSRSTN;
  wire delay_TL2ASPMSUSPENDCREDITCHECK;
  wire delay_TL2PPMSUSPENDREQ;
  wire delay_TLRSTN;
  wire delay_TRNRDSTRDY;
  wire delay_TRNRFCPRET;
  wire delay_TRNRNPOK;
  wire delay_TRNRNPREQ;
  wire delay_TRNTCFGGNT;
  wire delay_TRNTDLLPSRCRDY;
  wire delay_TRNTECRCGEN;
  wire delay_TRNTEOF;
  wire delay_TRNTERRFWD;
  wire delay_TRNTSOF;
  wire delay_TRNTSRCDSC;
  wire delay_TRNTSRCRDY;
  wire delay_TRNTSTR;
  wire delay_USERCLK2;
  wire delay_USERCLK;


   //drp monitor
   reg drpen_r1 = 1'b0;
   reg drpen_r2 = 1'b0;
   reg drpwe_r1 = 1'b0;
   reg drpwe_r2 = 1'b0;
   
   reg [1:0] sfsm = 2'b01;
    
   localparam FSM_IDLE = 2'b01;  
   localparam FSM_WAIT = 2'b10;
  

   always @(posedge delay_DRPCLK)
     begin
	// pipeline the DRPEN and DRPWE
        drpen_r1 <= delay_DRPEN;
        drpwe_r1 <= delay_DRPWE;
	drpen_r2 <= drpen_r1;
        drpwe_r2 <= drpwe_r1;

	
	// Check -  if DRPEN or DRPWE is more than 1 DCLK
	if ((drpen_r1 == 1'b1) && (drpen_r2 == 1'b1)) 
	  begin
	     $display("DRC Error : DRPEN is high for more than 1 DRPCLK on %m instance");
	     $finish; 
          end
	
	if ((drpwe_r1 == 1'b1) && (drpwe_r2 == 1'b1))
	  begin
             $display("DRC Error : DRPWE is high for more than 1 DRPCLK on %m instance");
             $finish;
          end


	//After the 1st DRPEN pulse, check the DRPEN and DRPRDY.
	case (sfsm)
          FSM_IDLE:   
            begin
               if(delay_DRPEN == 1'b1)
		 sfsm <= FSM_WAIT;  
            end
          
          FSM_WAIT:
            begin
               // After the 1st DRPEN, 4 cases can happen
               // DRPEN DRPRDY NEXT STATE
               // 0     0      FSM_WAIT - wait for DRPRDY
               // 0     1      FSM_IDLE - normal operation
               // 1     0      FSM_WAIT - display error and wait for DRPRDY
               // 1     1      FSM_WAIT - normal operation. Per UG470, DRPEN and DRPRDY can be at the same cycle.
               
               //Add the check for another DPREN pulse
               if(delay_DRPEN === 1'b1 && delay_DRPRDY === 1'b0) 
		 begin
		    $display("DRC Error : DRPEN is enabled before DRPRDY returns on %m instance");  
		    $finish;
		 end

               //Add the check for another DRPWE pulse
               if ((delay_DRPWE === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    $display("DRC Error : DRPWE is enabled before DRPRDY returns on %m instance");
		    $finish;
		 end
                    
               if ((delay_DRPRDY === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    sfsm <= FSM_IDLE;
		 end  
               
               if ((delay_DRPRDY === 1'b1)&& (delay_DRPEN === 1'b1))
		 begin
		    sfsm <= FSM_WAIT;
		 end  
            end
        
          default:                  
            begin
               $display("DRC Error : Default state in DRP FSM.");
               $finish;
            end
	endcase

     end // always @ (posedge delay_DRPCLK)
   //end drp monitor   

   
  assign #(out_delay) CFGAERECRCCHECKEN = delay_CFGAERECRCCHECKEN;
  assign #(out_delay) CFGAERECRCGENEN = delay_CFGAERECRCGENEN;
  assign #(out_delay) CFGAERROOTERRCORRERRRECEIVED = delay_CFGAERROOTERRCORRERRRECEIVED;
  assign #(out_delay) CFGAERROOTERRCORRERRREPORTINGEN = delay_CFGAERROOTERRCORRERRREPORTINGEN;
  assign #(out_delay) CFGAERROOTERRFATALERRRECEIVED = delay_CFGAERROOTERRFATALERRRECEIVED;
  assign #(out_delay) CFGAERROOTERRFATALERRREPORTINGEN = delay_CFGAERROOTERRFATALERRREPORTINGEN;
  assign #(out_delay) CFGAERROOTERRNONFATALERRRECEIVED = delay_CFGAERROOTERRNONFATALERRRECEIVED;
  assign #(out_delay) CFGAERROOTERRNONFATALERRREPORTINGEN = delay_CFGAERROOTERRNONFATALERRREPORTINGEN;
  assign #(out_delay) CFGBRIDGESERREN = delay_CFGBRIDGESERREN;
  assign #(out_delay) CFGCOMMANDBUSMASTERENABLE = delay_CFGCOMMANDBUSMASTERENABLE;
  assign #(out_delay) CFGCOMMANDINTERRUPTDISABLE = delay_CFGCOMMANDINTERRUPTDISABLE;
  assign #(out_delay) CFGCOMMANDIOENABLE = delay_CFGCOMMANDIOENABLE;
  assign #(out_delay) CFGCOMMANDMEMENABLE = delay_CFGCOMMANDMEMENABLE;
  assign #(out_delay) CFGCOMMANDSERREN = delay_CFGCOMMANDSERREN;
  assign #(out_delay) CFGDEVCONTROL2ARIFORWARDEN = delay_CFGDEVCONTROL2ARIFORWARDEN;
  assign #(out_delay) CFGDEVCONTROL2ATOMICEGRESSBLOCK = delay_CFGDEVCONTROL2ATOMICEGRESSBLOCK;
  assign #(out_delay) CFGDEVCONTROL2ATOMICREQUESTEREN = delay_CFGDEVCONTROL2ATOMICREQUESTEREN;
  assign #(out_delay) CFGDEVCONTROL2CPLTIMEOUTDIS = delay_CFGDEVCONTROL2CPLTIMEOUTDIS;
  assign #(out_delay) CFGDEVCONTROL2CPLTIMEOUTVAL = delay_CFGDEVCONTROL2CPLTIMEOUTVAL;
  assign #(out_delay) CFGDEVCONTROL2IDOCPLEN = delay_CFGDEVCONTROL2IDOCPLEN;
  assign #(out_delay) CFGDEVCONTROL2IDOREQEN = delay_CFGDEVCONTROL2IDOREQEN;
  assign #(out_delay) CFGDEVCONTROL2LTREN = delay_CFGDEVCONTROL2LTREN;
  assign #(out_delay) CFGDEVCONTROL2TLPPREFIXBLOCK = delay_CFGDEVCONTROL2TLPPREFIXBLOCK;
  assign #(out_delay) CFGDEVCONTROLAUXPOWEREN = delay_CFGDEVCONTROLAUXPOWEREN;
  assign #(out_delay) CFGDEVCONTROLCORRERRREPORTINGEN = delay_CFGDEVCONTROLCORRERRREPORTINGEN;
  assign #(out_delay) CFGDEVCONTROLENABLERO = delay_CFGDEVCONTROLENABLERO;
  assign #(out_delay) CFGDEVCONTROLEXTTAGEN = delay_CFGDEVCONTROLEXTTAGEN;
  assign #(out_delay) CFGDEVCONTROLFATALERRREPORTINGEN = delay_CFGDEVCONTROLFATALERRREPORTINGEN;
  assign #(out_delay) CFGDEVCONTROLMAXPAYLOAD = delay_CFGDEVCONTROLMAXPAYLOAD;
  assign #(out_delay) CFGDEVCONTROLMAXREADREQ = delay_CFGDEVCONTROLMAXREADREQ;
  assign #(out_delay) CFGDEVCONTROLNONFATALREPORTINGEN = delay_CFGDEVCONTROLNONFATALREPORTINGEN;
  assign #(out_delay) CFGDEVCONTROLNOSNOOPEN = delay_CFGDEVCONTROLNOSNOOPEN;
  assign #(out_delay) CFGDEVCONTROLPHANTOMEN = delay_CFGDEVCONTROLPHANTOMEN;
  assign #(out_delay) CFGDEVCONTROLURERRREPORTINGEN = delay_CFGDEVCONTROLURERRREPORTINGEN;
  assign #(out_delay) CFGDEVSTATUSCORRERRDETECTED = delay_CFGDEVSTATUSCORRERRDETECTED;
  assign #(out_delay) CFGDEVSTATUSFATALERRDETECTED = delay_CFGDEVSTATUSFATALERRDETECTED;
  assign #(out_delay) CFGDEVSTATUSNONFATALERRDETECTED = delay_CFGDEVSTATUSNONFATALERRDETECTED;
  assign #(out_delay) CFGDEVSTATUSURDETECTED = delay_CFGDEVSTATUSURDETECTED;
  assign #(out_delay) CFGERRAERHEADERLOGSETN = delay_CFGERRAERHEADERLOGSETN;
  assign #(out_delay) CFGERRCPLRDYN = delay_CFGERRCPLRDYN;
  assign #(out_delay) CFGINTERRUPTDO = delay_CFGINTERRUPTDO;
  assign #(out_delay) CFGINTERRUPTMMENABLE = delay_CFGINTERRUPTMMENABLE;
  assign #(out_delay) CFGINTERRUPTMSIENABLE = delay_CFGINTERRUPTMSIENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXENABLE = delay_CFGINTERRUPTMSIXENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXFM = delay_CFGINTERRUPTMSIXFM;
  assign #(out_delay) CFGINTERRUPTRDYN = delay_CFGINTERRUPTRDYN;
  assign #(out_delay) CFGLINKCONTROLASPMCONTROL = delay_CFGLINKCONTROLASPMCONTROL;
  assign #(out_delay) CFGLINKCONTROLAUTOBANDWIDTHINTEN = delay_CFGLINKCONTROLAUTOBANDWIDTHINTEN;
  assign #(out_delay) CFGLINKCONTROLBANDWIDTHINTEN = delay_CFGLINKCONTROLBANDWIDTHINTEN;
  assign #(out_delay) CFGLINKCONTROLCLOCKPMEN = delay_CFGLINKCONTROLCLOCKPMEN;
  assign #(out_delay) CFGLINKCONTROLCOMMONCLOCK = delay_CFGLINKCONTROLCOMMONCLOCK;
  assign #(out_delay) CFGLINKCONTROLEXTENDEDSYNC = delay_CFGLINKCONTROLEXTENDEDSYNC;
  assign #(out_delay) CFGLINKCONTROLHWAUTOWIDTHDIS = delay_CFGLINKCONTROLHWAUTOWIDTHDIS;
  assign #(out_delay) CFGLINKCONTROLLINKDISABLE = delay_CFGLINKCONTROLLINKDISABLE;
  assign #(out_delay) CFGLINKCONTROLRCB = delay_CFGLINKCONTROLRCB;
  assign #(out_delay) CFGLINKCONTROLRETRAINLINK = delay_CFGLINKCONTROLRETRAINLINK;
  assign #(out_delay) CFGLINKSTATUSAUTOBANDWIDTHSTATUS = delay_CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
  assign #(out_delay) CFGLINKSTATUSBANDWIDTHSTATUS = delay_CFGLINKSTATUSBANDWIDTHSTATUS;
  assign #(out_delay) CFGLINKSTATUSCURRENTSPEED = delay_CFGLINKSTATUSCURRENTSPEED;
  assign #(out_delay) CFGLINKSTATUSDLLACTIVE = delay_CFGLINKSTATUSDLLACTIVE;
  assign #(out_delay) CFGLINKSTATUSLINKTRAINING = delay_CFGLINKSTATUSLINKTRAINING;
  assign #(out_delay) CFGLINKSTATUSNEGOTIATEDWIDTH = delay_CFGLINKSTATUSNEGOTIATEDWIDTH;
  assign #(out_delay) CFGMGMTDO = delay_CFGMGMTDO;
  assign #(out_delay) CFGMGMTRDWRDONEN = delay_CFGMGMTRDWRDONEN;
  assign #(out_delay) CFGMSGDATA = delay_CFGMSGDATA;
  assign #(out_delay) CFGMSGRECEIVED = delay_CFGMSGRECEIVED;
  assign #(out_delay) CFGMSGRECEIVEDASSERTINTA = delay_CFGMSGRECEIVEDASSERTINTA;
  assign #(out_delay) CFGMSGRECEIVEDASSERTINTB = delay_CFGMSGRECEIVEDASSERTINTB;
  assign #(out_delay) CFGMSGRECEIVEDASSERTINTC = delay_CFGMSGRECEIVEDASSERTINTC;
  assign #(out_delay) CFGMSGRECEIVEDASSERTINTD = delay_CFGMSGRECEIVEDASSERTINTD;
  assign #(out_delay) CFGMSGRECEIVEDDEASSERTINTA = delay_CFGMSGRECEIVEDDEASSERTINTA;
  assign #(out_delay) CFGMSGRECEIVEDDEASSERTINTB = delay_CFGMSGRECEIVEDDEASSERTINTB;
  assign #(out_delay) CFGMSGRECEIVEDDEASSERTINTC = delay_CFGMSGRECEIVEDDEASSERTINTC;
  assign #(out_delay) CFGMSGRECEIVEDDEASSERTINTD = delay_CFGMSGRECEIVEDDEASSERTINTD;
  assign #(out_delay) CFGMSGRECEIVEDERRCOR = delay_CFGMSGRECEIVEDERRCOR;
  assign #(out_delay) CFGMSGRECEIVEDERRFATAL = delay_CFGMSGRECEIVEDERRFATAL;
  assign #(out_delay) CFGMSGRECEIVEDERRNONFATAL = delay_CFGMSGRECEIVEDERRNONFATAL;
  assign #(out_delay) CFGMSGRECEIVEDPMASNAK = delay_CFGMSGRECEIVEDPMASNAK;
  assign #(out_delay) CFGMSGRECEIVEDPMETO = delay_CFGMSGRECEIVEDPMETO;
  assign #(out_delay) CFGMSGRECEIVEDPMETOACK = delay_CFGMSGRECEIVEDPMETOACK;
  assign #(out_delay) CFGMSGRECEIVEDPMPME = delay_CFGMSGRECEIVEDPMPME;
  assign #(out_delay) CFGMSGRECEIVEDSETSLOTPOWERLIMIT = delay_CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
  assign #(out_delay) CFGMSGRECEIVEDUNLOCK = delay_CFGMSGRECEIVEDUNLOCK;
  assign #(out_delay) CFGPCIELINKSTATE = delay_CFGPCIELINKSTATE;
  assign #(out_delay) CFGPMCSRPMEEN = delay_CFGPMCSRPMEEN;
  assign #(out_delay) CFGPMCSRPMESTATUS = delay_CFGPMCSRPMESTATUS;
  assign #(out_delay) CFGPMCSRPOWERSTATE = delay_CFGPMCSRPOWERSTATE;
  assign #(out_delay) CFGPMRCVASREQL1N = delay_CFGPMRCVASREQL1N;
  assign #(out_delay) CFGPMRCVENTERL1N = delay_CFGPMRCVENTERL1N;
  assign #(out_delay) CFGPMRCVENTERL23N = delay_CFGPMRCVENTERL23N;
  assign #(out_delay) CFGPMRCVREQACKN = delay_CFGPMRCVREQACKN;
  assign #(out_delay) CFGROOTCONTROLPMEINTEN = delay_CFGROOTCONTROLPMEINTEN;
  assign #(out_delay) CFGROOTCONTROLSYSERRCORRERREN = delay_CFGROOTCONTROLSYSERRCORRERREN;
  assign #(out_delay) CFGROOTCONTROLSYSERRFATALERREN = delay_CFGROOTCONTROLSYSERRFATALERREN;
  assign #(out_delay) CFGROOTCONTROLSYSERRNONFATALERREN = delay_CFGROOTCONTROLSYSERRNONFATALERREN;
  assign #(out_delay) CFGSLOTCONTROLELECTROMECHILCTLPULSE = delay_CFGSLOTCONTROLELECTROMECHILCTLPULSE;
  assign #(out_delay) CFGTRANSACTION = delay_CFGTRANSACTION;
  assign #(out_delay) CFGTRANSACTIONADDR = delay_CFGTRANSACTIONADDR;
  assign #(out_delay) CFGTRANSACTIONTYPE = delay_CFGTRANSACTIONTYPE;
  assign #(out_delay) CFGVCTCVCMAP = delay_CFGVCTCVCMAP;
  assign #(out_delay) DBGSCLRA = delay_DBGSCLRA;
  assign #(out_delay) DBGSCLRB = delay_DBGSCLRB;
  assign #(out_delay) DBGSCLRC = delay_DBGSCLRC;
  assign #(out_delay) DBGSCLRD = delay_DBGSCLRD;
  assign #(out_delay) DBGSCLRE = delay_DBGSCLRE;
  assign #(out_delay) DBGSCLRF = delay_DBGSCLRF;
  assign #(out_delay) DBGSCLRG = delay_DBGSCLRG;
  assign #(out_delay) DBGSCLRH = delay_DBGSCLRH;
  assign #(out_delay) DBGSCLRI = delay_DBGSCLRI;
  assign #(out_delay) DBGSCLRJ = delay_DBGSCLRJ;
  assign #(out_delay) DBGSCLRK = delay_DBGSCLRK;
  assign #(out_delay) DBGVECA = delay_DBGVECA;
  assign #(out_delay) DBGVECB = delay_DBGVECB;
  assign #(out_delay) DBGVECC = delay_DBGVECC;
  assign #(out_delay) DRPDO = delay_DRPDO;
  assign #(out_delay) DRPRDY = delay_DRPRDY;
  assign #(out_delay) LL2BADDLLPERR = delay_LL2BADDLLPERR;
  assign #(out_delay) LL2BADTLPERR = delay_LL2BADTLPERR;
  assign #(out_delay) LL2LINKSTATUS = delay_LL2LINKSTATUS;
  assign #(out_delay) LL2PROTOCOLERR = delay_LL2PROTOCOLERR;
  assign #(out_delay) LL2RECEIVERERR = delay_LL2RECEIVERERR;
  assign #(out_delay) LL2REPLAYROERR = delay_LL2REPLAYROERR;
  assign #(out_delay) LL2REPLAYTOERR = delay_LL2REPLAYTOERR;
  assign #(out_delay) LL2SUSPENDOK = delay_LL2SUSPENDOK;
  assign #(out_delay) LL2TFCINIT1SEQ = delay_LL2TFCINIT1SEQ;
  assign #(out_delay) LL2TFCINIT2SEQ = delay_LL2TFCINIT2SEQ;
  assign #(out_delay) LL2TXIDLE = delay_LL2TXIDLE;
  assign #(out_delay) LNKCLKEN = delay_LNKCLKEN;
  assign #(out_delay) MIMRXRADDR = delay_MIMRXRADDR;
  assign #(out_delay) MIMRXREN = delay_MIMRXREN;
  assign #(out_delay) MIMRXWADDR = delay_MIMRXWADDR;
  assign #(out_delay) MIMRXWDATA = delay_MIMRXWDATA;
  assign #(out_delay) MIMRXWEN = delay_MIMRXWEN;
  assign #(out_delay) MIMTXRADDR = delay_MIMTXRADDR;
  assign #(out_delay) MIMTXREN = delay_MIMTXREN;
  assign #(out_delay) MIMTXWADDR = delay_MIMTXWADDR;
  assign #(out_delay) MIMTXWDATA = delay_MIMTXWDATA;
  assign #(out_delay) MIMTXWEN = delay_MIMTXWEN;
  assign #(out_delay) PIPERX0POLARITY = delay_PIPERX0POLARITY;
  assign #(out_delay) PIPERX1POLARITY = delay_PIPERX1POLARITY;
  assign #(out_delay) PIPERX2POLARITY = delay_PIPERX2POLARITY;
  assign #(out_delay) PIPERX3POLARITY = delay_PIPERX3POLARITY;
  assign #(out_delay) PIPERX4POLARITY = delay_PIPERX4POLARITY;
  assign #(out_delay) PIPERX5POLARITY = delay_PIPERX5POLARITY;
  assign #(out_delay) PIPERX6POLARITY = delay_PIPERX6POLARITY;
  assign #(out_delay) PIPERX7POLARITY = delay_PIPERX7POLARITY;
  assign #(out_delay) PIPETX0CHARISK = delay_PIPETX0CHARISK;
  assign #(out_delay) PIPETX0COMPLIANCE = delay_PIPETX0COMPLIANCE;
  assign #(out_delay) PIPETX0DATA = delay_PIPETX0DATA;
  assign #(out_delay) PIPETX0ELECIDLE = delay_PIPETX0ELECIDLE;
  assign #(out_delay) PIPETX0POWERDOWN = delay_PIPETX0POWERDOWN;
  assign #(out_delay) PIPETX1CHARISK = delay_PIPETX1CHARISK;
  assign #(out_delay) PIPETX1COMPLIANCE = delay_PIPETX1COMPLIANCE;
  assign #(out_delay) PIPETX1DATA = delay_PIPETX1DATA;
  assign #(out_delay) PIPETX1ELECIDLE = delay_PIPETX1ELECIDLE;
  assign #(out_delay) PIPETX1POWERDOWN = delay_PIPETX1POWERDOWN;
  assign #(out_delay) PIPETX2CHARISK = delay_PIPETX2CHARISK;
  assign #(out_delay) PIPETX2COMPLIANCE = delay_PIPETX2COMPLIANCE;
  assign #(out_delay) PIPETX2DATA = delay_PIPETX2DATA;
  assign #(out_delay) PIPETX2ELECIDLE = delay_PIPETX2ELECIDLE;
  assign #(out_delay) PIPETX2POWERDOWN = delay_PIPETX2POWERDOWN;
  assign #(out_delay) PIPETX3CHARISK = delay_PIPETX3CHARISK;
  assign #(out_delay) PIPETX3COMPLIANCE = delay_PIPETX3COMPLIANCE;
  assign #(out_delay) PIPETX3DATA = delay_PIPETX3DATA;
  assign #(out_delay) PIPETX3ELECIDLE = delay_PIPETX3ELECIDLE;
  assign #(out_delay) PIPETX3POWERDOWN = delay_PIPETX3POWERDOWN;
  assign #(out_delay) PIPETX4CHARISK = delay_PIPETX4CHARISK;
  assign #(out_delay) PIPETX4COMPLIANCE = delay_PIPETX4COMPLIANCE;
  assign #(out_delay) PIPETX4DATA = delay_PIPETX4DATA;
  assign #(out_delay) PIPETX4ELECIDLE = delay_PIPETX4ELECIDLE;
  assign #(out_delay) PIPETX4POWERDOWN = delay_PIPETX4POWERDOWN;
  assign #(out_delay) PIPETX5CHARISK = delay_PIPETX5CHARISK;
  assign #(out_delay) PIPETX5COMPLIANCE = delay_PIPETX5COMPLIANCE;
  assign #(out_delay) PIPETX5DATA = delay_PIPETX5DATA;
  assign #(out_delay) PIPETX5ELECIDLE = delay_PIPETX5ELECIDLE;
  assign #(out_delay) PIPETX5POWERDOWN = delay_PIPETX5POWERDOWN;
  assign #(out_delay) PIPETX6CHARISK = delay_PIPETX6CHARISK;
  assign #(out_delay) PIPETX6COMPLIANCE = delay_PIPETX6COMPLIANCE;
  assign #(out_delay) PIPETX6DATA = delay_PIPETX6DATA;
  assign #(out_delay) PIPETX6ELECIDLE = delay_PIPETX6ELECIDLE;
  assign #(out_delay) PIPETX6POWERDOWN = delay_PIPETX6POWERDOWN;
  assign #(out_delay) PIPETX7CHARISK = delay_PIPETX7CHARISK;
  assign #(out_delay) PIPETX7COMPLIANCE = delay_PIPETX7COMPLIANCE;
  assign #(out_delay) PIPETX7DATA = delay_PIPETX7DATA;
  assign #(out_delay) PIPETX7ELECIDLE = delay_PIPETX7ELECIDLE;
  assign #(out_delay) PIPETX7POWERDOWN = delay_PIPETX7POWERDOWN;
  assign #(out_delay) PIPETXDEEMPH = delay_PIPETXDEEMPH;
  assign #(out_delay) PIPETXMARGIN = delay_PIPETXMARGIN;
  assign #(out_delay) PIPETXRATE = delay_PIPETXRATE;
  assign #(out_delay) PIPETXRCVRDET = delay_PIPETXRCVRDET;
  assign #(out_delay) PIPETXRESET = delay_PIPETXRESET;
  assign #(out_delay) PL2L0REQ = delay_PL2L0REQ;
  assign #(out_delay) PL2LINKUP = delay_PL2LINKUP;
  assign #(out_delay) PL2RECEIVERERR = delay_PL2RECEIVERERR;
  assign #(out_delay) PL2RECOVERY = delay_PL2RECOVERY;
  assign #(out_delay) PL2RXELECIDLE = delay_PL2RXELECIDLE;
  assign #(out_delay) PL2RXPMSTATE = delay_PL2RXPMSTATE;
  assign #(out_delay) PL2SUSPENDOK = delay_PL2SUSPENDOK;
  assign #(out_delay) PLDBGVEC = delay_PLDBGVEC;
  assign #(out_delay) PLDIRECTEDCHANGEDONE = delay_PLDIRECTEDCHANGEDONE;
  assign #(out_delay) PLINITIALLINKWIDTH = delay_PLINITIALLINKWIDTH;
  assign #(out_delay) PLLANEREVERSALMODE = delay_PLLANEREVERSALMODE;
  assign #(out_delay) PLLINKGEN2CAP = delay_PLLINKGEN2CAP;
  assign #(out_delay) PLLINKPARTNERGEN2SUPPORTED = delay_PLLINKPARTNERGEN2SUPPORTED;
  assign #(out_delay) PLLINKUPCFGCAP = delay_PLLINKUPCFGCAP;
  assign #(out_delay) PLLTSSMSTATE = delay_PLLTSSMSTATE;
  assign #(out_delay) PLPHYLNKUPN = delay_PLPHYLNKUPN;
  assign #(out_delay) PLRECEIVEDHOTRST = delay_PLRECEIVEDHOTRST;
  assign #(out_delay) PLRXPMSTATE = delay_PLRXPMSTATE;
  assign #(out_delay) PLSELLNKRATE = delay_PLSELLNKRATE;
  assign #(out_delay) PLSELLNKWIDTH = delay_PLSELLNKWIDTH;
  assign #(out_delay) PLTXPMSTATE = delay_PLTXPMSTATE;
  assign #(out_delay) RECEIVEDFUNCLVLRSTN = delay_RECEIVEDFUNCLVLRSTN;
  assign #(out_delay) TL2ASPMSUSPENDCREDITCHECKOK = delay_TL2ASPMSUSPENDCREDITCHECKOK;
  assign #(out_delay) TL2ASPMSUSPENDREQ = delay_TL2ASPMSUSPENDREQ;
  assign #(out_delay) TL2ERRFCPE = delay_TL2ERRFCPE;
  assign #(out_delay) TL2ERRHDR = delay_TL2ERRHDR;
  assign #(out_delay) TL2ERRMALFORMED = delay_TL2ERRMALFORMED;
  assign #(out_delay) TL2ERRRXOVERFLOW = delay_TL2ERRRXOVERFLOW;
  assign #(out_delay) TL2PPMSUSPENDOK = delay_TL2PPMSUSPENDOK;
  assign #(out_delay) TRNFCCPLD = delay_TRNFCCPLD;
  assign #(out_delay) TRNFCCPLH = delay_TRNFCCPLH;
  assign #(out_delay) TRNFCNPD = delay_TRNFCNPD;
  assign #(out_delay) TRNFCNPH = delay_TRNFCNPH;
  assign #(out_delay) TRNFCPD = delay_TRNFCPD;
  assign #(out_delay) TRNFCPH = delay_TRNFCPH;
  assign #(out_delay) TRNLNKUP = delay_TRNLNKUP;
  assign #(out_delay) TRNRBARHIT = delay_TRNRBARHIT;
  assign #(out_delay) TRNRD = delay_TRNRD;
  assign #(out_delay) TRNRDLLPDATA = delay_TRNRDLLPDATA;
  assign #(out_delay) TRNRDLLPSRCRDY = delay_TRNRDLLPSRCRDY;
  assign #(out_delay) TRNRECRCERR = delay_TRNRECRCERR;
  assign #(out_delay) TRNREOF = delay_TRNREOF;
  assign #(out_delay) TRNRERRFWD = delay_TRNRERRFWD;
  assign #(out_delay) TRNRREM = delay_TRNRREM;
  assign #(out_delay) TRNRSOF = delay_TRNRSOF;
  assign #(out_delay) TRNRSRCDSC = delay_TRNRSRCDSC;
  assign #(out_delay) TRNRSRCRDY = delay_TRNRSRCRDY;
  assign #(out_delay) TRNTBUFAV = delay_TRNTBUFAV;
  assign #(out_delay) TRNTCFGREQ = delay_TRNTCFGREQ;
  assign #(out_delay) TRNTDLLPDSTRDY = delay_TRNTDLLPDSTRDY;
  assign #(out_delay) TRNTDSTRDY = delay_TRNTDSTRDY;
  assign #(out_delay) TRNTERRDROP = delay_TRNTERRDROP;
  assign #(out_delay) USERRSTN = delay_USERRSTN;
  
`ifndef XIL_TIMING // unisim
  assign #(INCLK_DELAY) delay_DRPCLK = DRPCLK;
  assign #(INCLK_DELAY) delay_PIPECLK = PIPECLK;
  assign #(INCLK_DELAY) delay_USERCLK = USERCLK;
  assign #(INCLK_DELAY) delay_USERCLK2 = USERCLK2;

  assign #(in_delay) delay_CFGAERINTERRUPTMSGNUM = CFGAERINTERRUPTMSGNUM;
  assign #(in_delay) delay_CFGDEVID = CFGDEVID;
  assign #(in_delay) delay_CFGDSBUSNUMBER = CFGDSBUSNUMBER;
  assign #(in_delay) delay_CFGDSDEVICENUMBER = CFGDSDEVICENUMBER;
  assign #(in_delay) delay_CFGDSFUNCTIONNUMBER = CFGDSFUNCTIONNUMBER;
  assign #(in_delay) delay_CFGDSN = CFGDSN;
  assign #(in_delay) delay_CFGERRACSN = CFGERRACSN;
  assign #(in_delay) delay_CFGERRAERHEADERLOG = CFGERRAERHEADERLOG;
  assign #(in_delay) delay_CFGERRATOMICEGRESSBLOCKEDN = CFGERRATOMICEGRESSBLOCKEDN;
  assign #(in_delay) delay_CFGERRCORN = CFGERRCORN;
  assign #(in_delay) delay_CFGERRCPLABORTN = CFGERRCPLABORTN;
  assign #(in_delay) delay_CFGERRCPLTIMEOUTN = CFGERRCPLTIMEOUTN;
  assign #(in_delay) delay_CFGERRCPLUNEXPECTN = CFGERRCPLUNEXPECTN;
  assign #(in_delay) delay_CFGERRECRCN = CFGERRECRCN;
  assign #(in_delay) delay_CFGERRINTERNALCORN = CFGERRINTERNALCORN;
  assign #(in_delay) delay_CFGERRINTERNALUNCORN = CFGERRINTERNALUNCORN;
  assign #(in_delay) delay_CFGERRLOCKEDN = CFGERRLOCKEDN;
  assign #(in_delay) delay_CFGERRMALFORMEDN = CFGERRMALFORMEDN;
  assign #(in_delay) delay_CFGERRMCBLOCKEDN = CFGERRMCBLOCKEDN;
  assign #(in_delay) delay_CFGERRNORECOVERYN = CFGERRNORECOVERYN;
  assign #(in_delay) delay_CFGERRPOISONEDN = CFGERRPOISONEDN;
  assign #(in_delay) delay_CFGERRPOSTEDN = CFGERRPOSTEDN;
  assign #(in_delay) delay_CFGERRTLPCPLHEADER = CFGERRTLPCPLHEADER;
  assign #(in_delay) delay_CFGERRURN = CFGERRURN;
  assign #(in_delay) delay_CFGFORCECOMMONCLOCKOFF = CFGFORCECOMMONCLOCKOFF;
  assign #(in_delay) delay_CFGFORCEEXTENDEDSYNCON = CFGFORCEEXTENDEDSYNCON;
  assign #(in_delay) delay_CFGFORCEMPS = CFGFORCEMPS;
  assign #(in_delay) delay_CFGINTERRUPTASSERTN = CFGINTERRUPTASSERTN;
  assign #(in_delay) delay_CFGINTERRUPTDI = CFGINTERRUPTDI;
  assign #(in_delay) delay_CFGINTERRUPTN = CFGINTERRUPTN;
  assign #(in_delay) delay_CFGINTERRUPTSTATN = CFGINTERRUPTSTATN;
  assign #(in_delay) delay_CFGMGMTBYTEENN = CFGMGMTBYTEENN;
  assign #(in_delay) delay_CFGMGMTDI = CFGMGMTDI;
  assign #(in_delay) delay_CFGMGMTDWADDR = CFGMGMTDWADDR;
  assign #(in_delay) delay_CFGMGMTRDENN = CFGMGMTRDENN;
  assign #(in_delay) delay_CFGMGMTWRENN = CFGMGMTWRENN;
  assign #(in_delay) delay_CFGMGMTWRREADONLYN = CFGMGMTWRREADONLYN;
  assign #(in_delay) delay_CFGMGMTWRRW1CASRWN = CFGMGMTWRRW1CASRWN;
  assign #(in_delay) delay_CFGPCIECAPINTERRUPTMSGNUM = CFGPCIECAPINTERRUPTMSGNUM;
  assign #(in_delay) delay_CFGPMFORCESTATE = CFGPMFORCESTATE;
  assign #(in_delay) delay_CFGPMFORCESTATEENN = CFGPMFORCESTATEENN;
  assign #(in_delay) delay_CFGPMHALTASPML0SN = CFGPMHALTASPML0SN;
  assign #(in_delay) delay_CFGPMHALTASPML1N = CFGPMHALTASPML1N;
  assign #(in_delay) delay_CFGPMSENDPMETON = CFGPMSENDPMETON;
  assign #(in_delay) delay_CFGPMTURNOFFOKN = CFGPMTURNOFFOKN;
  assign #(in_delay) delay_CFGPMWAKEN = CFGPMWAKEN;
  assign #(in_delay) delay_CFGPORTNUMBER = CFGPORTNUMBER;
  assign #(in_delay) delay_CFGREVID = CFGREVID;
  assign #(in_delay) delay_CFGSUBSYSID = CFGSUBSYSID;
  assign #(in_delay) delay_CFGSUBSYSVENDID = CFGSUBSYSVENDID;
  assign #(in_delay) delay_CFGTRNPENDINGN = CFGTRNPENDINGN;
  assign #(in_delay) delay_CFGVENDID = CFGVENDID;
  assign #(in_delay) delay_CMRSTN = CMRSTN;
  assign #(in_delay) delay_CMSTICKYRSTN = CMSTICKYRSTN;
  assign #(in_delay) delay_DBGMODE = DBGMODE;
  assign #(in_delay) delay_DBGSUBMODE = DBGSUBMODE;
  assign #(in_delay) delay_DLRSTN = DLRSTN;
  assign #(in_delay) delay_DRPADDR = DRPADDR;
  assign #(in_delay) delay_DRPDI = DRPDI;
  assign #(in_delay) delay_DRPEN = DRPEN;
  assign #(in_delay) delay_DRPWE = DRPWE;
  assign #(in_delay) delay_FUNCLVLRSTN = FUNCLVLRSTN;
  assign #(in_delay) delay_LL2SENDASREQL1 = LL2SENDASREQL1;
  assign #(in_delay) delay_LL2SENDENTERL1 = LL2SENDENTERL1;
  assign #(in_delay) delay_LL2SENDENTERL23 = LL2SENDENTERL23;
  assign #(in_delay) delay_LL2SENDPMACK = LL2SENDPMACK;
  assign #(in_delay) delay_LL2SUSPENDNOW = LL2SUSPENDNOW;
  assign #(in_delay) delay_LL2TLPRCV = LL2TLPRCV;
  assign #(in_delay) delay_MIMRXRDATA = MIMRXRDATA;
  assign #(in_delay) delay_MIMTXRDATA = MIMTXRDATA;
  assign #(in_delay) delay_PIPERX0CHANISALIGNED = PIPERX0CHANISALIGNED;
  assign #(in_delay) delay_PIPERX0CHARISK = PIPERX0CHARISK;
  assign #(in_delay) delay_PIPERX0DATA = PIPERX0DATA;
  assign #(in_delay) delay_PIPERX0ELECIDLE = PIPERX0ELECIDLE;
  assign #(in_delay) delay_PIPERX0PHYSTATUS = PIPERX0PHYSTATUS;
  assign #(in_delay) delay_PIPERX0STATUS = PIPERX0STATUS;
  assign #(in_delay) delay_PIPERX0VALID = PIPERX0VALID;
  assign #(in_delay) delay_PIPERX1CHANISALIGNED = PIPERX1CHANISALIGNED;
  assign #(in_delay) delay_PIPERX1CHARISK = PIPERX1CHARISK;
  assign #(in_delay) delay_PIPERX1DATA = PIPERX1DATA;
  assign #(in_delay) delay_PIPERX1ELECIDLE = PIPERX1ELECIDLE;
  assign #(in_delay) delay_PIPERX1PHYSTATUS = PIPERX1PHYSTATUS;
  assign #(in_delay) delay_PIPERX1STATUS = PIPERX1STATUS;
  assign #(in_delay) delay_PIPERX1VALID = PIPERX1VALID;
  assign #(in_delay) delay_PIPERX2CHANISALIGNED = PIPERX2CHANISALIGNED;
  assign #(in_delay) delay_PIPERX2CHARISK = PIPERX2CHARISK;
  assign #(in_delay) delay_PIPERX2DATA = PIPERX2DATA;
  assign #(in_delay) delay_PIPERX2ELECIDLE = PIPERX2ELECIDLE;
  assign #(in_delay) delay_PIPERX2PHYSTATUS = PIPERX2PHYSTATUS;
  assign #(in_delay) delay_PIPERX2STATUS = PIPERX2STATUS;
  assign #(in_delay) delay_PIPERX2VALID = PIPERX2VALID;
  assign #(in_delay) delay_PIPERX3CHANISALIGNED = PIPERX3CHANISALIGNED;
  assign #(in_delay) delay_PIPERX3CHARISK = PIPERX3CHARISK;
  assign #(in_delay) delay_PIPERX3DATA = PIPERX3DATA;
  assign #(in_delay) delay_PIPERX3ELECIDLE = PIPERX3ELECIDLE;
  assign #(in_delay) delay_PIPERX3PHYSTATUS = PIPERX3PHYSTATUS;
  assign #(in_delay) delay_PIPERX3STATUS = PIPERX3STATUS;
  assign #(in_delay) delay_PIPERX3VALID = PIPERX3VALID;
  assign #(in_delay) delay_PIPERX4CHANISALIGNED = PIPERX4CHANISALIGNED;
  assign #(in_delay) delay_PIPERX4CHARISK = PIPERX4CHARISK;
  assign #(in_delay) delay_PIPERX4DATA = PIPERX4DATA;
  assign #(in_delay) delay_PIPERX4ELECIDLE = PIPERX4ELECIDLE;
  assign #(in_delay) delay_PIPERX4PHYSTATUS = PIPERX4PHYSTATUS;
  assign #(in_delay) delay_PIPERX4STATUS = PIPERX4STATUS;
  assign #(in_delay) delay_PIPERX4VALID = PIPERX4VALID;
  assign #(in_delay) delay_PIPERX5CHANISALIGNED = PIPERX5CHANISALIGNED;
  assign #(in_delay) delay_PIPERX5CHARISK = PIPERX5CHARISK;
  assign #(in_delay) delay_PIPERX5DATA = PIPERX5DATA;
  assign #(in_delay) delay_PIPERX5ELECIDLE = PIPERX5ELECIDLE;
  assign #(in_delay) delay_PIPERX5PHYSTATUS = PIPERX5PHYSTATUS;
  assign #(in_delay) delay_PIPERX5STATUS = PIPERX5STATUS;
  assign #(in_delay) delay_PIPERX5VALID = PIPERX5VALID;
  assign #(in_delay) delay_PIPERX6CHANISALIGNED = PIPERX6CHANISALIGNED;
  assign #(in_delay) delay_PIPERX6CHARISK = PIPERX6CHARISK;
  assign #(in_delay) delay_PIPERX6DATA = PIPERX6DATA;
  assign #(in_delay) delay_PIPERX6ELECIDLE = PIPERX6ELECIDLE;
  assign #(in_delay) delay_PIPERX6PHYSTATUS = PIPERX6PHYSTATUS;
  assign #(in_delay) delay_PIPERX6STATUS = PIPERX6STATUS;
  assign #(in_delay) delay_PIPERX6VALID = PIPERX6VALID;
  assign #(in_delay) delay_PIPERX7CHANISALIGNED = PIPERX7CHANISALIGNED;
  assign #(in_delay) delay_PIPERX7CHARISK = PIPERX7CHARISK;
  assign #(in_delay) delay_PIPERX7DATA = PIPERX7DATA;
  assign #(in_delay) delay_PIPERX7ELECIDLE = PIPERX7ELECIDLE;
  assign #(in_delay) delay_PIPERX7PHYSTATUS = PIPERX7PHYSTATUS;
  assign #(in_delay) delay_PIPERX7STATUS = PIPERX7STATUS;
  assign #(in_delay) delay_PIPERX7VALID = PIPERX7VALID;
  assign #(in_delay) delay_PL2DIRECTEDLSTATE = PL2DIRECTEDLSTATE;
  assign #(in_delay) delay_PLDBGMODE = PLDBGMODE;
  assign #(in_delay) delay_PLDIRECTEDLINKAUTON = PLDIRECTEDLINKAUTON;
  assign #(in_delay) delay_PLDIRECTEDLINKCHANGE = PLDIRECTEDLINKCHANGE;
  assign #(in_delay) delay_PLDIRECTEDLINKSPEED = PLDIRECTEDLINKSPEED;
  assign #(in_delay) delay_PLDIRECTEDLINKWIDTH = PLDIRECTEDLINKWIDTH;
  assign #(in_delay) delay_PLDIRECTEDLTSSMNEW = PLDIRECTEDLTSSMNEW;
  assign #(in_delay) delay_PLDIRECTEDLTSSMNEWVLD = PLDIRECTEDLTSSMNEWVLD;
  assign #(in_delay) delay_PLDIRECTEDLTSSMSTALL = PLDIRECTEDLTSSMSTALL;
  assign #(in_delay) delay_PLDOWNSTREAMDEEMPHSOURCE = PLDOWNSTREAMDEEMPHSOURCE;
  assign #(in_delay) delay_PLRSTN = PLRSTN;
  assign #(in_delay) delay_PLTRANSMITHOTRST = PLTRANSMITHOTRST;
  assign #(in_delay) delay_PLUPSTREAMPREFERDEEMPH = PLUPSTREAMPREFERDEEMPH;
  assign #(in_delay) delay_SYSRSTN = SYSRSTN;
  assign #(in_delay) delay_TL2ASPMSUSPENDCREDITCHECK = TL2ASPMSUSPENDCREDITCHECK;
  assign #(in_delay) delay_TL2PPMSUSPENDREQ = TL2PPMSUSPENDREQ;
  assign #(in_delay) delay_TLRSTN = TLRSTN;
  assign #(in_delay) delay_TRNFCSEL = TRNFCSEL;
  assign #(in_delay) delay_TRNRDSTRDY = TRNRDSTRDY;
  assign #(in_delay) delay_TRNRFCPRET = TRNRFCPRET;
  assign #(in_delay) delay_TRNRNPOK = TRNRNPOK;
  assign #(in_delay) delay_TRNRNPREQ = TRNRNPREQ;
  assign #(in_delay) delay_TRNTCFGGNT = TRNTCFGGNT;
  assign #(in_delay) delay_TRNTD = TRNTD;
  assign #(in_delay) delay_TRNTDLLPDATA = TRNTDLLPDATA;
  assign #(in_delay) delay_TRNTDLLPSRCRDY = TRNTDLLPSRCRDY;
  assign #(in_delay) delay_TRNTECRCGEN = TRNTECRCGEN;
  assign #(in_delay) delay_TRNTEOF = TRNTEOF;
  assign #(in_delay) delay_TRNTERRFWD = TRNTERRFWD;
  assign #(in_delay) delay_TRNTREM = TRNTREM;
  assign #(in_delay) delay_TRNTSOF = TRNTSOF;
  assign #(in_delay) delay_TRNTSRCDSC = TRNTSRCDSC;
  assign #(in_delay) delay_TRNTSRCRDY = TRNTSRCRDY;
  assign #(in_delay) delay_TRNTSTR = TRNTSTR;
`endif //  `ifndef XIL_TIMING

`ifdef XIL_TIMING //Simprim
  assign delay_SYSRSTN = SYSRSTN;
`endif

  B_PCIE_2_1 #(
    .AER_BASE_PTR (AER_BASE_PTR),
    .AER_CAP_ECRC_CHECK_CAPABLE (AER_CAP_ECRC_CHECK_CAPABLE),
    .AER_CAP_ECRC_GEN_CAPABLE (AER_CAP_ECRC_GEN_CAPABLE),
    .AER_CAP_ID (AER_CAP_ID),
    .AER_CAP_MULTIHEADER (AER_CAP_MULTIHEADER),
    .AER_CAP_NEXTPTR (AER_CAP_NEXTPTR),
    .AER_CAP_ON (AER_CAP_ON),
    .AER_CAP_OPTIONAL_ERR_SUPPORT (AER_CAP_OPTIONAL_ERR_SUPPORT),
    .AER_CAP_PERMIT_ROOTERR_UPDATE (AER_CAP_PERMIT_ROOTERR_UPDATE),
    .AER_CAP_VERSION (AER_CAP_VERSION),
    .ALLOW_X8_GEN2 (ALLOW_X8_GEN2),
    .BAR0 (BAR0),
    .BAR1 (BAR1),
    .BAR2 (BAR2),
    .BAR3 (BAR3),
    .BAR4 (BAR4),
    .BAR5 (BAR5),
    .CAPABILITIES_PTR (CAPABILITIES_PTR),
    .CARDBUS_CIS_POINTER (CARDBUS_CIS_POINTER),
    .CFG_ECRC_ERR_CPLSTAT (CFG_ECRC_ERR_CPLSTAT),
    .CLASS_CODE (CLASS_CODE),
    .CMD_INTX_IMPLEMENTED (CMD_INTX_IMPLEMENTED),
    .CPL_TIMEOUT_DISABLE_SUPPORTED (CPL_TIMEOUT_DISABLE_SUPPORTED),
    .CPL_TIMEOUT_RANGES_SUPPORTED (CPL_TIMEOUT_RANGES_SUPPORTED),
    .CRM_MODULE_RSTS (CRM_MODULE_RSTS),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED (DEV_CAP2_ARI_FORWARDING_SUPPORTED),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED (DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED (DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED (DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED (DEV_CAP2_CAS128_COMPLETER_SUPPORTED),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED (DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED (DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED (DEV_CAP2_LTR_MECHANISM_SUPPORTED),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES (DEV_CAP2_MAX_ENDEND_TLP_PREFIXES),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING (DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED (DEV_CAP2_TPH_COMPLETER_SUPPORTED),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE (DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE (DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE),
    .DEV_CAP_ENDPOINT_L0S_LATENCY (DEV_CAP_ENDPOINT_L0S_LATENCY),
    .DEV_CAP_ENDPOINT_L1_LATENCY (DEV_CAP_ENDPOINT_L1_LATENCY),
    .DEV_CAP_EXT_TAG_SUPPORTED (DEV_CAP_EXT_TAG_SUPPORTED),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE (DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED (DEV_CAP_MAX_PAYLOAD_SUPPORTED),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT (DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT),
    .DEV_CAP_ROLE_BASED_ERROR (DEV_CAP_ROLE_BASED_ERROR),
    .DEV_CAP_RSVD_14_12 (DEV_CAP_RSVD_14_12),
    .DEV_CAP_RSVD_17_16 (DEV_CAP_RSVD_17_16),
    .DEV_CAP_RSVD_31_29 (DEV_CAP_RSVD_31_29),
    .DEV_CONTROL_AUX_POWER_SUPPORTED (DEV_CONTROL_AUX_POWER_SUPPORTED),
    .DEV_CONTROL_EXT_TAG_DEFAULT (DEV_CONTROL_EXT_TAG_DEFAULT),
    .DISABLE_ASPM_L1_TIMER (DISABLE_ASPM_L1_TIMER),
    .DISABLE_BAR_FILTERING (DISABLE_BAR_FILTERING),
    .DISABLE_ERR_MSG (DISABLE_ERR_MSG),
    .DISABLE_ID_CHECK (DISABLE_ID_CHECK),
    .DISABLE_LANE_REVERSAL (DISABLE_LANE_REVERSAL),
    .DISABLE_LOCKED_FILTER (DISABLE_LOCKED_FILTER),
    .DISABLE_PPM_FILTER (DISABLE_PPM_FILTER),
    .DISABLE_RX_POISONED_RESP (DISABLE_RX_POISONED_RESP),
    .DISABLE_RX_TC_FILTER (DISABLE_RX_TC_FILTER),
    .DISABLE_SCRAMBLING (DISABLE_SCRAMBLING),
    .DNSTREAM_LINK_NUM (DNSTREAM_LINK_NUM),
    .DSN_BASE_PTR (DSN_BASE_PTR),
    .DSN_CAP_ID (DSN_CAP_ID),
    .DSN_CAP_NEXTPTR (DSN_CAP_NEXTPTR),
    .DSN_CAP_ON (DSN_CAP_ON),
    .DSN_CAP_VERSION (DSN_CAP_VERSION),
    .ENABLE_MSG_ROUTE (ENABLE_MSG_ROUTE),
    .ENABLE_RX_TD_ECRC_TRIM (ENABLE_RX_TD_ECRC_TRIM),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED (ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED),
    .ENTER_RVRY_EI_L0 (ENTER_RVRY_EI_L0),
    .EXIT_LOOPBACK_ON_EI (EXIT_LOOPBACK_ON_EI),
    .EXPANSION_ROM (EXPANSION_ROM),
    .EXT_CFG_CAP_PTR (EXT_CFG_CAP_PTR),
    .EXT_CFG_XP_CAP_PTR (EXT_CFG_XP_CAP_PTR),
    .HEADER_TYPE (HEADER_TYPE),
    .INFER_EI (INFER_EI),
    .INTERRUPT_PIN (INTERRUPT_PIN),
    .INTERRUPT_STAT_AUTO (INTERRUPT_STAT_AUTO),
    .IS_SWITCH (IS_SWITCH),
    .LAST_CONFIG_DWORD (LAST_CONFIG_DWORD),
    .LINK_CAP_ASPM_OPTIONALITY (LINK_CAP_ASPM_OPTIONALITY),
    .LINK_CAP_ASPM_SUPPORT (LINK_CAP_ASPM_SUPPORT),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT (LINK_CAP_CLOCK_POWER_MANAGEMENT),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP (LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 (LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 (LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1 (LINK_CAP_L0S_EXIT_LATENCY_GEN1),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2 (LINK_CAP_L0S_EXIT_LATENCY_GEN2),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 (LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 (LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1 (LINK_CAP_L1_EXIT_LATENCY_GEN1),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2 (LINK_CAP_L1_EXIT_LATENCY_GEN2),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP (LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP),
    .LINK_CAP_MAX_LINK_SPEED (LINK_CAP_MAX_LINK_SPEED),
    .LINK_CAP_MAX_LINK_WIDTH (LINK_CAP_MAX_LINK_WIDTH),
    .LINK_CAP_RSVD_23 (LINK_CAP_RSVD_23),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE (LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE),
    .LINK_CONTROL_RCB (LINK_CONTROL_RCB),
    .LINK_CTRL2_DEEMPHASIS (LINK_CTRL2_DEEMPHASIS),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE (LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE),
    .LINK_CTRL2_TARGET_LINK_SPEED (LINK_CTRL2_TARGET_LINK_SPEED),
    .LINK_STATUS_SLOT_CLOCK_CONFIG (LINK_STATUS_SLOT_CLOCK_CONFIG),
    .LL_ACK_TIMEOUT (LL_ACK_TIMEOUT),
    .LL_ACK_TIMEOUT_EN (LL_ACK_TIMEOUT_EN),
    .LL_ACK_TIMEOUT_FUNC (LL_ACK_TIMEOUT_FUNC),
    .LL_REPLAY_TIMEOUT (LL_REPLAY_TIMEOUT),
    .LL_REPLAY_TIMEOUT_EN (LL_REPLAY_TIMEOUT_EN),
    .LL_REPLAY_TIMEOUT_FUNC (LL_REPLAY_TIMEOUT_FUNC),
    .LTSSM_MAX_LINK_WIDTH (LTSSM_MAX_LINK_WIDTH),
    .MPS_FORCE (MPS_FORCE),
    .MSIX_BASE_PTR (MSIX_BASE_PTR),
    .MSIX_CAP_ID (MSIX_CAP_ID),
    .MSIX_CAP_NEXTPTR (MSIX_CAP_NEXTPTR),
    .MSIX_CAP_ON (MSIX_CAP_ON),
    .MSIX_CAP_PBA_BIR (MSIX_CAP_PBA_BIR),
    .MSIX_CAP_PBA_OFFSET (MSIX_CAP_PBA_OFFSET),
    .MSIX_CAP_TABLE_BIR (MSIX_CAP_TABLE_BIR),
    .MSIX_CAP_TABLE_OFFSET (MSIX_CAP_TABLE_OFFSET),
    .MSIX_CAP_TABLE_SIZE (MSIX_CAP_TABLE_SIZE),
    .MSI_BASE_PTR (MSI_BASE_PTR),
    .MSI_CAP_64_BIT_ADDR_CAPABLE (MSI_CAP_64_BIT_ADDR_CAPABLE),
    .MSI_CAP_ID (MSI_CAP_ID),
    .MSI_CAP_MULTIMSGCAP (MSI_CAP_MULTIMSGCAP),
    .MSI_CAP_MULTIMSG_EXTENSION (MSI_CAP_MULTIMSG_EXTENSION),
    .MSI_CAP_NEXTPTR (MSI_CAP_NEXTPTR),
    .MSI_CAP_ON (MSI_CAP_ON),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE (MSI_CAP_PER_VECTOR_MASKING_CAPABLE),
    .N_FTS_COMCLK_GEN1 (N_FTS_COMCLK_GEN1),
    .N_FTS_COMCLK_GEN2 (N_FTS_COMCLK_GEN2),
    .N_FTS_GEN1 (N_FTS_GEN1),
    .N_FTS_GEN2 (N_FTS_GEN2),
    .PCIE_BASE_PTR (PCIE_BASE_PTR),
    .PCIE_CAP_CAPABILITY_ID (PCIE_CAP_CAPABILITY_ID),
    .PCIE_CAP_CAPABILITY_VERSION (PCIE_CAP_CAPABILITY_VERSION),
    .PCIE_CAP_DEVICE_PORT_TYPE (PCIE_CAP_DEVICE_PORT_TYPE),
    .PCIE_CAP_NEXTPTR (PCIE_CAP_NEXTPTR),
    .PCIE_CAP_ON (PCIE_CAP_ON),
    .PCIE_CAP_RSVD_15_14 (PCIE_CAP_RSVD_15_14),
    .PCIE_CAP_SLOT_IMPLEMENTED (PCIE_CAP_SLOT_IMPLEMENTED),
    .PCIE_REVISION (PCIE_REVISION),
    .PL_AUTO_CONFIG (PL_AUTO_CONFIG),
    .PL_FAST_TRAIN (PL_FAST_TRAIN),
    .PM_ASPML0S_TIMEOUT (PM_ASPML0S_TIMEOUT),
    .PM_ASPML0S_TIMEOUT_EN (PM_ASPML0S_TIMEOUT_EN),
    .PM_ASPML0S_TIMEOUT_FUNC (PM_ASPML0S_TIMEOUT_FUNC),
    .PM_ASPM_FASTEXIT (PM_ASPM_FASTEXIT),
    .PM_BASE_PTR (PM_BASE_PTR),
    .PM_CAP_AUXCURRENT (PM_CAP_AUXCURRENT),
    .PM_CAP_D1SUPPORT (PM_CAP_D1SUPPORT),
    .PM_CAP_D2SUPPORT (PM_CAP_D2SUPPORT),
    .PM_CAP_DSI (PM_CAP_DSI),
    .PM_CAP_ID (PM_CAP_ID),
    .PM_CAP_NEXTPTR (PM_CAP_NEXTPTR),
    .PM_CAP_ON (PM_CAP_ON),
    .PM_CAP_PMESUPPORT (PM_CAP_PMESUPPORT),
    .PM_CAP_PME_CLOCK (PM_CAP_PME_CLOCK),
    .PM_CAP_RSVD_04 (PM_CAP_RSVD_04),
    .PM_CAP_VERSION (PM_CAP_VERSION),
    .PM_CSR_B2B3 (PM_CSR_B2B3),
    .PM_CSR_BPCCEN (PM_CSR_BPCCEN),
    .PM_CSR_NOSOFTRST (PM_CSR_NOSOFTRST),
    .PM_DATA0 (PM_DATA0),
    .PM_DATA1 (PM_DATA1),
    .PM_DATA2 (PM_DATA2),
    .PM_DATA3 (PM_DATA3),
    .PM_DATA4 (PM_DATA4),
    .PM_DATA5 (PM_DATA5),
    .PM_DATA6 (PM_DATA6),
    .PM_DATA7 (PM_DATA7),
    .PM_DATA_SCALE0 (PM_DATA_SCALE0),
    .PM_DATA_SCALE1 (PM_DATA_SCALE1),
    .PM_DATA_SCALE2 (PM_DATA_SCALE2),
    .PM_DATA_SCALE3 (PM_DATA_SCALE3),
    .PM_DATA_SCALE4 (PM_DATA_SCALE4),
    .PM_DATA_SCALE5 (PM_DATA_SCALE5),
    .PM_DATA_SCALE6 (PM_DATA_SCALE6),
    .PM_DATA_SCALE7 (PM_DATA_SCALE7),
    .PM_MF (PM_MF),
    .RBAR_BASE_PTR (RBAR_BASE_PTR),
    .RBAR_CAP_CONTROL_ENCODEDBAR0 (RBAR_CAP_CONTROL_ENCODEDBAR0),
    .RBAR_CAP_CONTROL_ENCODEDBAR1 (RBAR_CAP_CONTROL_ENCODEDBAR1),
    .RBAR_CAP_CONTROL_ENCODEDBAR2 (RBAR_CAP_CONTROL_ENCODEDBAR2),
    .RBAR_CAP_CONTROL_ENCODEDBAR3 (RBAR_CAP_CONTROL_ENCODEDBAR3),
    .RBAR_CAP_CONTROL_ENCODEDBAR4 (RBAR_CAP_CONTROL_ENCODEDBAR4),
    .RBAR_CAP_CONTROL_ENCODEDBAR5 (RBAR_CAP_CONTROL_ENCODEDBAR5),
    .RBAR_CAP_ID (RBAR_CAP_ID),
    .RBAR_CAP_INDEX0 (RBAR_CAP_INDEX0),
    .RBAR_CAP_INDEX1 (RBAR_CAP_INDEX1),
    .RBAR_CAP_INDEX2 (RBAR_CAP_INDEX2),
    .RBAR_CAP_INDEX3 (RBAR_CAP_INDEX3),
    .RBAR_CAP_INDEX4 (RBAR_CAP_INDEX4),
    .RBAR_CAP_INDEX5 (RBAR_CAP_INDEX5),
    .RBAR_CAP_NEXTPTR (RBAR_CAP_NEXTPTR),
    .RBAR_CAP_ON (RBAR_CAP_ON),
    .RBAR_CAP_SUP0 (RBAR_CAP_SUP0),
    .RBAR_CAP_SUP1 (RBAR_CAP_SUP1),
    .RBAR_CAP_SUP2 (RBAR_CAP_SUP2),
    .RBAR_CAP_SUP3 (RBAR_CAP_SUP3),
    .RBAR_CAP_SUP4 (RBAR_CAP_SUP4),
    .RBAR_CAP_SUP5 (RBAR_CAP_SUP5),
    .RBAR_CAP_VERSION (RBAR_CAP_VERSION),
    .RBAR_NUM (RBAR_NUM),
    .RECRC_CHK (RECRC_CHK),
    .RECRC_CHK_TRIM (RECRC_CHK_TRIM),
    .ROOT_CAP_CRS_SW_VISIBILITY (ROOT_CAP_CRS_SW_VISIBILITY),
    .RP_AUTO_SPD (RP_AUTO_SPD),
    .RP_AUTO_SPD_LOOPCNT (RP_AUTO_SPD_LOOPCNT),
    .SELECT_DLL_IF (SELECT_DLL_IF),
    .SIM_VERSION (SIM_VERSION),
    .SLOT_CAP_ATT_BUTTON_PRESENT (SLOT_CAP_ATT_BUTTON_PRESENT),
    .SLOT_CAP_ATT_INDICATOR_PRESENT (SLOT_CAP_ATT_INDICATOR_PRESENT),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT (SLOT_CAP_ELEC_INTERLOCK_PRESENT),
    .SLOT_CAP_HOTPLUG_CAPABLE (SLOT_CAP_HOTPLUG_CAPABLE),
    .SLOT_CAP_HOTPLUG_SURPRISE (SLOT_CAP_HOTPLUG_SURPRISE),
    .SLOT_CAP_MRL_SENSOR_PRESENT (SLOT_CAP_MRL_SENSOR_PRESENT),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT (SLOT_CAP_NO_CMD_COMPLETED_SUPPORT),
    .SLOT_CAP_PHYSICAL_SLOT_NUM (SLOT_CAP_PHYSICAL_SLOT_NUM),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT (SLOT_CAP_POWER_CONTROLLER_PRESENT),
    .SLOT_CAP_POWER_INDICATOR_PRESENT (SLOT_CAP_POWER_INDICATOR_PRESENT),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE (SLOT_CAP_SLOT_POWER_LIMIT_SCALE),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE (SLOT_CAP_SLOT_POWER_LIMIT_VALUE),
    .SPARE_BIT0 (SPARE_BIT0),
    .SPARE_BIT1 (SPARE_BIT1),
    .SPARE_BIT2 (SPARE_BIT2),
    .SPARE_BIT3 (SPARE_BIT3),
    .SPARE_BIT4 (SPARE_BIT4),
    .SPARE_BIT5 (SPARE_BIT5),
    .SPARE_BIT6 (SPARE_BIT6),
    .SPARE_BIT7 (SPARE_BIT7),
    .SPARE_BIT8 (SPARE_BIT8),
    .SPARE_BYTE0 (SPARE_BYTE0),
    .SPARE_BYTE1 (SPARE_BYTE1),
    .SPARE_BYTE2 (SPARE_BYTE2),
    .SPARE_BYTE3 (SPARE_BYTE3),
    .SPARE_WORD0 (SPARE_WORD0),
    .SPARE_WORD1 (SPARE_WORD1),
    .SPARE_WORD2 (SPARE_WORD2),
    .SPARE_WORD3 (SPARE_WORD3),
    .SSL_MESSAGE_AUTO (SSL_MESSAGE_AUTO),
    .TECRC_EP_INV (TECRC_EP_INV),
    .TL_RBYPASS (TL_RBYPASS),
    .TL_RX_RAM_RADDR_LATENCY (TL_RX_RAM_RADDR_LATENCY),
    .TL_RX_RAM_RDATA_LATENCY (TL_RX_RAM_RDATA_LATENCY),
    .TL_RX_RAM_WRITE_LATENCY (TL_RX_RAM_WRITE_LATENCY),
    .TL_TFC_DISABLE (TL_TFC_DISABLE),
    .TL_TX_CHECKS_DISABLE (TL_TX_CHECKS_DISABLE),
    .TL_TX_RAM_RADDR_LATENCY (TL_TX_RAM_RADDR_LATENCY),
    .TL_TX_RAM_RDATA_LATENCY (TL_TX_RAM_RDATA_LATENCY),
    .TL_TX_RAM_WRITE_LATENCY (TL_TX_RAM_WRITE_LATENCY),
    .TRN_DW (TRN_DW),
    .TRN_NP_FC (TRN_NP_FC),
    .UPCONFIG_CAPABLE (UPCONFIG_CAPABLE),
    .UPSTREAM_FACING (UPSTREAM_FACING),
    .UR_ATOMIC (UR_ATOMIC),
    .UR_CFG1 (UR_CFG1),
    .UR_INV_REQ (UR_INV_REQ),
    .UR_PRS_RESPONSE (UR_PRS_RESPONSE),
    .USER_CLK2_DIV2 (USER_CLK2_DIV2),
    .USER_CLK_FREQ (USER_CLK_FREQ),
    .USE_RID_PINS (USE_RID_PINS),
    .VC0_CPL_INFINITE (VC0_CPL_INFINITE),
    .VC0_RX_RAM_LIMIT (VC0_RX_RAM_LIMIT),
    .VC0_TOTAL_CREDITS_CD (VC0_TOTAL_CREDITS_CD),
    .VC0_TOTAL_CREDITS_CH (VC0_TOTAL_CREDITS_CH),
    .VC0_TOTAL_CREDITS_NPD (VC0_TOTAL_CREDITS_NPD),
    .VC0_TOTAL_CREDITS_NPH (VC0_TOTAL_CREDITS_NPH),
    .VC0_TOTAL_CREDITS_PD (VC0_TOTAL_CREDITS_PD),
    .VC0_TOTAL_CREDITS_PH (VC0_TOTAL_CREDITS_PH),
    .VC0_TX_LASTPACKET (VC0_TX_LASTPACKET),
    .VC_BASE_PTR (VC_BASE_PTR),
    .VC_CAP_ID (VC_CAP_ID),
    .VC_CAP_NEXTPTR (VC_CAP_NEXTPTR),
    .VC_CAP_ON (VC_CAP_ON),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS (VC_CAP_REJECT_SNOOP_TRANSACTIONS),
    .VC_CAP_VERSION (VC_CAP_VERSION),
    .VSEC_BASE_PTR (VSEC_BASE_PTR),
    .VSEC_CAP_HDR_ID (VSEC_CAP_HDR_ID),
    .VSEC_CAP_HDR_LENGTH (VSEC_CAP_HDR_LENGTH),
    .VSEC_CAP_HDR_REVISION (VSEC_CAP_HDR_REVISION),
    .VSEC_CAP_ID (VSEC_CAP_ID),
    .VSEC_CAP_IS_LINK_VISIBLE (VSEC_CAP_IS_LINK_VISIBLE),
    .VSEC_CAP_NEXTPTR (VSEC_CAP_NEXTPTR),
    .VSEC_CAP_ON (VSEC_CAP_ON),
    .VSEC_CAP_VERSION (VSEC_CAP_VERSION))

    B_PCIE_2_1_INST (
    .CFGAERECRCCHECKEN (delay_CFGAERECRCCHECKEN),
    .CFGAERECRCGENEN (delay_CFGAERECRCGENEN),
    .CFGAERROOTERRCORRERRRECEIVED (delay_CFGAERROOTERRCORRERRRECEIVED),
    .CFGAERROOTERRCORRERRREPORTINGEN (delay_CFGAERROOTERRCORRERRREPORTINGEN),
    .CFGAERROOTERRFATALERRRECEIVED (delay_CFGAERROOTERRFATALERRRECEIVED),
    .CFGAERROOTERRFATALERRREPORTINGEN (delay_CFGAERROOTERRFATALERRREPORTINGEN),
    .CFGAERROOTERRNONFATALERRRECEIVED (delay_CFGAERROOTERRNONFATALERRRECEIVED),
    .CFGAERROOTERRNONFATALERRREPORTINGEN (delay_CFGAERROOTERRNONFATALERRREPORTINGEN),
    .CFGBRIDGESERREN (delay_CFGBRIDGESERREN),
    .CFGCOMMANDBUSMASTERENABLE (delay_CFGCOMMANDBUSMASTERENABLE),
    .CFGCOMMANDINTERRUPTDISABLE (delay_CFGCOMMANDINTERRUPTDISABLE),
    .CFGCOMMANDIOENABLE (delay_CFGCOMMANDIOENABLE),
    .CFGCOMMANDMEMENABLE (delay_CFGCOMMANDMEMENABLE),
    .CFGCOMMANDSERREN (delay_CFGCOMMANDSERREN),
    .CFGDEVCONTROL2ARIFORWARDEN (delay_CFGDEVCONTROL2ARIFORWARDEN),
    .CFGDEVCONTROL2ATOMICEGRESSBLOCK (delay_CFGDEVCONTROL2ATOMICEGRESSBLOCK),
    .CFGDEVCONTROL2ATOMICREQUESTEREN (delay_CFGDEVCONTROL2ATOMICREQUESTEREN),
    .CFGDEVCONTROL2CPLTIMEOUTDIS (delay_CFGDEVCONTROL2CPLTIMEOUTDIS),
    .CFGDEVCONTROL2CPLTIMEOUTVAL (delay_CFGDEVCONTROL2CPLTIMEOUTVAL),
    .CFGDEVCONTROL2IDOCPLEN (delay_CFGDEVCONTROL2IDOCPLEN),
    .CFGDEVCONTROL2IDOREQEN (delay_CFGDEVCONTROL2IDOREQEN),
    .CFGDEVCONTROL2LTREN (delay_CFGDEVCONTROL2LTREN),
    .CFGDEVCONTROL2TLPPREFIXBLOCK (delay_CFGDEVCONTROL2TLPPREFIXBLOCK),
    .CFGDEVCONTROLAUXPOWEREN (delay_CFGDEVCONTROLAUXPOWEREN),
    .CFGDEVCONTROLCORRERRREPORTINGEN (delay_CFGDEVCONTROLCORRERRREPORTINGEN),
    .CFGDEVCONTROLENABLERO (delay_CFGDEVCONTROLENABLERO),
    .CFGDEVCONTROLEXTTAGEN (delay_CFGDEVCONTROLEXTTAGEN),
    .CFGDEVCONTROLFATALERRREPORTINGEN (delay_CFGDEVCONTROLFATALERRREPORTINGEN),
    .CFGDEVCONTROLMAXPAYLOAD (delay_CFGDEVCONTROLMAXPAYLOAD),
    .CFGDEVCONTROLMAXREADREQ (delay_CFGDEVCONTROLMAXREADREQ),
    .CFGDEVCONTROLNONFATALREPORTINGEN (delay_CFGDEVCONTROLNONFATALREPORTINGEN),
    .CFGDEVCONTROLNOSNOOPEN (delay_CFGDEVCONTROLNOSNOOPEN),
    .CFGDEVCONTROLPHANTOMEN (delay_CFGDEVCONTROLPHANTOMEN),
    .CFGDEVCONTROLURERRREPORTINGEN (delay_CFGDEVCONTROLURERRREPORTINGEN),
    .CFGDEVSTATUSCORRERRDETECTED (delay_CFGDEVSTATUSCORRERRDETECTED),
    .CFGDEVSTATUSFATALERRDETECTED (delay_CFGDEVSTATUSFATALERRDETECTED),
    .CFGDEVSTATUSNONFATALERRDETECTED (delay_CFGDEVSTATUSNONFATALERRDETECTED),
    .CFGDEVSTATUSURDETECTED (delay_CFGDEVSTATUSURDETECTED),
    .CFGERRAERHEADERLOGSETN (delay_CFGERRAERHEADERLOGSETN),
    .CFGERRCPLRDYN (delay_CFGERRCPLRDYN),
    .CFGINTERRUPTDO (delay_CFGINTERRUPTDO),
    .CFGINTERRUPTMMENABLE (delay_CFGINTERRUPTMMENABLE),
    .CFGINTERRUPTMSIENABLE (delay_CFGINTERRUPTMSIENABLE),
    .CFGINTERRUPTMSIXENABLE (delay_CFGINTERRUPTMSIXENABLE),
    .CFGINTERRUPTMSIXFM (delay_CFGINTERRUPTMSIXFM),
    .CFGINTERRUPTRDYN (delay_CFGINTERRUPTRDYN),
    .CFGLINKCONTROLASPMCONTROL (delay_CFGLINKCONTROLASPMCONTROL),
    .CFGLINKCONTROLAUTOBANDWIDTHINTEN (delay_CFGLINKCONTROLAUTOBANDWIDTHINTEN),
    .CFGLINKCONTROLBANDWIDTHINTEN (delay_CFGLINKCONTROLBANDWIDTHINTEN),
    .CFGLINKCONTROLCLOCKPMEN (delay_CFGLINKCONTROLCLOCKPMEN),
    .CFGLINKCONTROLCOMMONCLOCK (delay_CFGLINKCONTROLCOMMONCLOCK),
    .CFGLINKCONTROLEXTENDEDSYNC (delay_CFGLINKCONTROLEXTENDEDSYNC),
    .CFGLINKCONTROLHWAUTOWIDTHDIS (delay_CFGLINKCONTROLHWAUTOWIDTHDIS),
    .CFGLINKCONTROLLINKDISABLE (delay_CFGLINKCONTROLLINKDISABLE),
    .CFGLINKCONTROLRCB (delay_CFGLINKCONTROLRCB),
    .CFGLINKCONTROLRETRAINLINK (delay_CFGLINKCONTROLRETRAINLINK),
    .CFGLINKSTATUSAUTOBANDWIDTHSTATUS (delay_CFGLINKSTATUSAUTOBANDWIDTHSTATUS),
    .CFGLINKSTATUSBANDWIDTHSTATUS (delay_CFGLINKSTATUSBANDWIDTHSTATUS),
    .CFGLINKSTATUSCURRENTSPEED (delay_CFGLINKSTATUSCURRENTSPEED),
    .CFGLINKSTATUSDLLACTIVE (delay_CFGLINKSTATUSDLLACTIVE),
    .CFGLINKSTATUSLINKTRAINING (delay_CFGLINKSTATUSLINKTRAINING),
    .CFGLINKSTATUSNEGOTIATEDWIDTH (delay_CFGLINKSTATUSNEGOTIATEDWIDTH),
    .CFGMGMTDO (delay_CFGMGMTDO),
    .CFGMGMTRDWRDONEN (delay_CFGMGMTRDWRDONEN),
    .CFGMSGDATA (delay_CFGMSGDATA),
    .CFGMSGRECEIVED (delay_CFGMSGRECEIVED),
    .CFGMSGRECEIVEDASSERTINTA (delay_CFGMSGRECEIVEDASSERTINTA),
    .CFGMSGRECEIVEDASSERTINTB (delay_CFGMSGRECEIVEDASSERTINTB),
    .CFGMSGRECEIVEDASSERTINTC (delay_CFGMSGRECEIVEDASSERTINTC),
    .CFGMSGRECEIVEDASSERTINTD (delay_CFGMSGRECEIVEDASSERTINTD),
    .CFGMSGRECEIVEDDEASSERTINTA (delay_CFGMSGRECEIVEDDEASSERTINTA),
    .CFGMSGRECEIVEDDEASSERTINTB (delay_CFGMSGRECEIVEDDEASSERTINTB),
    .CFGMSGRECEIVEDDEASSERTINTC (delay_CFGMSGRECEIVEDDEASSERTINTC),
    .CFGMSGRECEIVEDDEASSERTINTD (delay_CFGMSGRECEIVEDDEASSERTINTD),
    .CFGMSGRECEIVEDERRCOR (delay_CFGMSGRECEIVEDERRCOR),
    .CFGMSGRECEIVEDERRFATAL (delay_CFGMSGRECEIVEDERRFATAL),
    .CFGMSGRECEIVEDERRNONFATAL (delay_CFGMSGRECEIVEDERRNONFATAL),
    .CFGMSGRECEIVEDPMASNAK (delay_CFGMSGRECEIVEDPMASNAK),
    .CFGMSGRECEIVEDPMETO (delay_CFGMSGRECEIVEDPMETO),
    .CFGMSGRECEIVEDPMETOACK (delay_CFGMSGRECEIVEDPMETOACK),
    .CFGMSGRECEIVEDPMPME (delay_CFGMSGRECEIVEDPMPME),
    .CFGMSGRECEIVEDSETSLOTPOWERLIMIT (delay_CFGMSGRECEIVEDSETSLOTPOWERLIMIT),
    .CFGMSGRECEIVEDUNLOCK (delay_CFGMSGRECEIVEDUNLOCK),
    .CFGPCIELINKSTATE (delay_CFGPCIELINKSTATE),
    .CFGPMCSRPMEEN (delay_CFGPMCSRPMEEN),
    .CFGPMCSRPMESTATUS (delay_CFGPMCSRPMESTATUS),
    .CFGPMCSRPOWERSTATE (delay_CFGPMCSRPOWERSTATE),
    .CFGPMRCVASREQL1N (delay_CFGPMRCVASREQL1N),
    .CFGPMRCVENTERL1N (delay_CFGPMRCVENTERL1N),
    .CFGPMRCVENTERL23N (delay_CFGPMRCVENTERL23N),
    .CFGPMRCVREQACKN (delay_CFGPMRCVREQACKN),
    .CFGROOTCONTROLPMEINTEN (delay_CFGROOTCONTROLPMEINTEN),
    .CFGROOTCONTROLSYSERRCORRERREN (delay_CFGROOTCONTROLSYSERRCORRERREN),
    .CFGROOTCONTROLSYSERRFATALERREN (delay_CFGROOTCONTROLSYSERRFATALERREN),
    .CFGROOTCONTROLSYSERRNONFATALERREN (delay_CFGROOTCONTROLSYSERRNONFATALERREN),
    .CFGSLOTCONTROLELECTROMECHILCTLPULSE (delay_CFGSLOTCONTROLELECTROMECHILCTLPULSE),
    .CFGTRANSACTION (delay_CFGTRANSACTION),
    .CFGTRANSACTIONADDR (delay_CFGTRANSACTIONADDR),
    .CFGTRANSACTIONTYPE (delay_CFGTRANSACTIONTYPE),
    .CFGVCTCVCMAP (delay_CFGVCTCVCMAP),
    .DBGSCLRA (delay_DBGSCLRA),
    .DBGSCLRB (delay_DBGSCLRB),
    .DBGSCLRC (delay_DBGSCLRC),
    .DBGSCLRD (delay_DBGSCLRD),
    .DBGSCLRE (delay_DBGSCLRE),
    .DBGSCLRF (delay_DBGSCLRF),
    .DBGSCLRG (delay_DBGSCLRG),
    .DBGSCLRH (delay_DBGSCLRH),
    .DBGSCLRI (delay_DBGSCLRI),
    .DBGSCLRJ (delay_DBGSCLRJ),
    .DBGSCLRK (delay_DBGSCLRK),
    .DBGVECA (delay_DBGVECA),
    .DBGVECB (delay_DBGVECB),
    .DBGVECC (delay_DBGVECC),
    .DRPDO (delay_DRPDO),
    .DRPRDY (delay_DRPRDY),
    .LL2BADDLLPERR (delay_LL2BADDLLPERR),
    .LL2BADTLPERR (delay_LL2BADTLPERR),
    .LL2LINKSTATUS (delay_LL2LINKSTATUS),
    .LL2PROTOCOLERR (delay_LL2PROTOCOLERR),
    .LL2RECEIVERERR (delay_LL2RECEIVERERR),
    .LL2REPLAYROERR (delay_LL2REPLAYROERR),
    .LL2REPLAYTOERR (delay_LL2REPLAYTOERR),
    .LL2SUSPENDOK (delay_LL2SUSPENDOK),
    .LL2TFCINIT1SEQ (delay_LL2TFCINIT1SEQ),
    .LL2TFCINIT2SEQ (delay_LL2TFCINIT2SEQ),
    .LL2TXIDLE (delay_LL2TXIDLE),
    .LNKCLKEN (delay_LNKCLKEN),
    .MIMRXRADDR (delay_MIMRXRADDR),
    .MIMRXREN (delay_MIMRXREN),
    .MIMRXWADDR (delay_MIMRXWADDR),
    .MIMRXWDATA (delay_MIMRXWDATA),
    .MIMRXWEN (delay_MIMRXWEN),
    .MIMTXRADDR (delay_MIMTXRADDR),
    .MIMTXREN (delay_MIMTXREN),
    .MIMTXWADDR (delay_MIMTXWADDR),
    .MIMTXWDATA (delay_MIMTXWDATA),
    .MIMTXWEN (delay_MIMTXWEN),
    .PIPERX0POLARITY (delay_PIPERX0POLARITY),
    .PIPERX1POLARITY (delay_PIPERX1POLARITY),
    .PIPERX2POLARITY (delay_PIPERX2POLARITY),
    .PIPERX3POLARITY (delay_PIPERX3POLARITY),
    .PIPERX4POLARITY (delay_PIPERX4POLARITY),
    .PIPERX5POLARITY (delay_PIPERX5POLARITY),
    .PIPERX6POLARITY (delay_PIPERX6POLARITY),
    .PIPERX7POLARITY (delay_PIPERX7POLARITY),
    .PIPETX0CHARISK (delay_PIPETX0CHARISK),
    .PIPETX0COMPLIANCE (delay_PIPETX0COMPLIANCE),
    .PIPETX0DATA (delay_PIPETX0DATA),
    .PIPETX0ELECIDLE (delay_PIPETX0ELECIDLE),
    .PIPETX0POWERDOWN (delay_PIPETX0POWERDOWN),
    .PIPETX1CHARISK (delay_PIPETX1CHARISK),
    .PIPETX1COMPLIANCE (delay_PIPETX1COMPLIANCE),
    .PIPETX1DATA (delay_PIPETX1DATA),
    .PIPETX1ELECIDLE (delay_PIPETX1ELECIDLE),
    .PIPETX1POWERDOWN (delay_PIPETX1POWERDOWN),
    .PIPETX2CHARISK (delay_PIPETX2CHARISK),
    .PIPETX2COMPLIANCE (delay_PIPETX2COMPLIANCE),
    .PIPETX2DATA (delay_PIPETX2DATA),
    .PIPETX2ELECIDLE (delay_PIPETX2ELECIDLE),
    .PIPETX2POWERDOWN (delay_PIPETX2POWERDOWN),
    .PIPETX3CHARISK (delay_PIPETX3CHARISK),
    .PIPETX3COMPLIANCE (delay_PIPETX3COMPLIANCE),
    .PIPETX3DATA (delay_PIPETX3DATA),
    .PIPETX3ELECIDLE (delay_PIPETX3ELECIDLE),
    .PIPETX3POWERDOWN (delay_PIPETX3POWERDOWN),
    .PIPETX4CHARISK (delay_PIPETX4CHARISK),
    .PIPETX4COMPLIANCE (delay_PIPETX4COMPLIANCE),
    .PIPETX4DATA (delay_PIPETX4DATA),
    .PIPETX4ELECIDLE (delay_PIPETX4ELECIDLE),
    .PIPETX4POWERDOWN (delay_PIPETX4POWERDOWN),
    .PIPETX5CHARISK (delay_PIPETX5CHARISK),
    .PIPETX5COMPLIANCE (delay_PIPETX5COMPLIANCE),
    .PIPETX5DATA (delay_PIPETX5DATA),
    .PIPETX5ELECIDLE (delay_PIPETX5ELECIDLE),
    .PIPETX5POWERDOWN (delay_PIPETX5POWERDOWN),
    .PIPETX6CHARISK (delay_PIPETX6CHARISK),
    .PIPETX6COMPLIANCE (delay_PIPETX6COMPLIANCE),
    .PIPETX6DATA (delay_PIPETX6DATA),
    .PIPETX6ELECIDLE (delay_PIPETX6ELECIDLE),
    .PIPETX6POWERDOWN (delay_PIPETX6POWERDOWN),
    .PIPETX7CHARISK (delay_PIPETX7CHARISK),
    .PIPETX7COMPLIANCE (delay_PIPETX7COMPLIANCE),
    .PIPETX7DATA (delay_PIPETX7DATA),
    .PIPETX7ELECIDLE (delay_PIPETX7ELECIDLE),
    .PIPETX7POWERDOWN (delay_PIPETX7POWERDOWN),
    .PIPETXDEEMPH (delay_PIPETXDEEMPH),
    .PIPETXMARGIN (delay_PIPETXMARGIN),
    .PIPETXRATE (delay_PIPETXRATE),
    .PIPETXRCVRDET (delay_PIPETXRCVRDET),
    .PIPETXRESET (delay_PIPETXRESET),
    .PL2L0REQ (delay_PL2L0REQ),
    .PL2LINKUP (delay_PL2LINKUP),
    .PL2RECEIVERERR (delay_PL2RECEIVERERR),
    .PL2RECOVERY (delay_PL2RECOVERY),
    .PL2RXELECIDLE (delay_PL2RXELECIDLE),
    .PL2RXPMSTATE (delay_PL2RXPMSTATE),
    .PL2SUSPENDOK (delay_PL2SUSPENDOK),
    .PLDBGVEC (delay_PLDBGVEC),
    .PLDIRECTEDCHANGEDONE (delay_PLDIRECTEDCHANGEDONE),
    .PLINITIALLINKWIDTH (delay_PLINITIALLINKWIDTH),
    .PLLANEREVERSALMODE (delay_PLLANEREVERSALMODE),
    .PLLINKGEN2CAP (delay_PLLINKGEN2CAP),
    .PLLINKPARTNERGEN2SUPPORTED (delay_PLLINKPARTNERGEN2SUPPORTED),
    .PLLINKUPCFGCAP (delay_PLLINKUPCFGCAP),
    .PLLTSSMSTATE (delay_PLLTSSMSTATE),
    .PLPHYLNKUPN (delay_PLPHYLNKUPN),
    .PLRECEIVEDHOTRST (delay_PLRECEIVEDHOTRST),
    .PLRXPMSTATE (delay_PLRXPMSTATE),
    .PLSELLNKRATE (delay_PLSELLNKRATE),
    .PLSELLNKWIDTH (delay_PLSELLNKWIDTH),
    .PLTXPMSTATE (delay_PLTXPMSTATE),
    .RECEIVEDFUNCLVLRSTN (delay_RECEIVEDFUNCLVLRSTN),
    .TL2ASPMSUSPENDCREDITCHECKOK (delay_TL2ASPMSUSPENDCREDITCHECKOK),
    .TL2ASPMSUSPENDREQ (delay_TL2ASPMSUSPENDREQ),
    .TL2ERRFCPE (delay_TL2ERRFCPE),
    .TL2ERRHDR (delay_TL2ERRHDR),
    .TL2ERRMALFORMED (delay_TL2ERRMALFORMED),
    .TL2ERRRXOVERFLOW (delay_TL2ERRRXOVERFLOW),
    .TL2PPMSUSPENDOK (delay_TL2PPMSUSPENDOK),
    .TRNFCCPLD (delay_TRNFCCPLD),
    .TRNFCCPLH (delay_TRNFCCPLH),
    .TRNFCNPD (delay_TRNFCNPD),
    .TRNFCNPH (delay_TRNFCNPH),
    .TRNFCPD (delay_TRNFCPD),
    .TRNFCPH (delay_TRNFCPH),
    .TRNLNKUP (delay_TRNLNKUP),
    .TRNRBARHIT (delay_TRNRBARHIT),
    .TRNRD (delay_TRNRD),
    .TRNRDLLPDATA (delay_TRNRDLLPDATA),
    .TRNRDLLPSRCRDY (delay_TRNRDLLPSRCRDY),
    .TRNRECRCERR (delay_TRNRECRCERR),
    .TRNREOF (delay_TRNREOF),
    .TRNRERRFWD (delay_TRNRERRFWD),
    .TRNRREM (delay_TRNRREM),
    .TRNRSOF (delay_TRNRSOF),
    .TRNRSRCDSC (delay_TRNRSRCDSC),
    .TRNRSRCRDY (delay_TRNRSRCRDY),
    .TRNTBUFAV (delay_TRNTBUFAV),
    .TRNTCFGREQ (delay_TRNTCFGREQ),
    .TRNTDLLPDSTRDY (delay_TRNTDLLPDSTRDY),
    .TRNTDSTRDY (delay_TRNTDSTRDY),
    .TRNTERRDROP (delay_TRNTERRDROP),
    .USERRSTN (delay_USERRSTN),
    .CFGAERINTERRUPTMSGNUM (delay_CFGAERINTERRUPTMSGNUM),
    .CFGDEVID (delay_CFGDEVID),
    .CFGDSBUSNUMBER (delay_CFGDSBUSNUMBER),
    .CFGDSDEVICENUMBER (delay_CFGDSDEVICENUMBER),
    .CFGDSFUNCTIONNUMBER (delay_CFGDSFUNCTIONNUMBER),
    .CFGDSN (delay_CFGDSN),
    .CFGERRACSN (delay_CFGERRACSN),
    .CFGERRAERHEADERLOG (delay_CFGERRAERHEADERLOG),
    .CFGERRATOMICEGRESSBLOCKEDN (delay_CFGERRATOMICEGRESSBLOCKEDN),
    .CFGERRCORN (delay_CFGERRCORN),
    .CFGERRCPLABORTN (delay_CFGERRCPLABORTN),
    .CFGERRCPLTIMEOUTN (delay_CFGERRCPLTIMEOUTN),
    .CFGERRCPLUNEXPECTN (delay_CFGERRCPLUNEXPECTN),
    .CFGERRECRCN (delay_CFGERRECRCN),
    .CFGERRINTERNALCORN (delay_CFGERRINTERNALCORN),
    .CFGERRINTERNALUNCORN (delay_CFGERRINTERNALUNCORN),
    .CFGERRLOCKEDN (delay_CFGERRLOCKEDN),
    .CFGERRMALFORMEDN (delay_CFGERRMALFORMEDN),
    .CFGERRMCBLOCKEDN (delay_CFGERRMCBLOCKEDN),
    .CFGERRNORECOVERYN (delay_CFGERRNORECOVERYN),
    .CFGERRPOISONEDN (delay_CFGERRPOISONEDN),
    .CFGERRPOSTEDN (delay_CFGERRPOSTEDN),
    .CFGERRTLPCPLHEADER (delay_CFGERRTLPCPLHEADER),
    .CFGERRURN (delay_CFGERRURN),
    .CFGFORCECOMMONCLOCKOFF (delay_CFGFORCECOMMONCLOCKOFF),
    .CFGFORCEEXTENDEDSYNCON (delay_CFGFORCEEXTENDEDSYNCON),
    .CFGFORCEMPS (delay_CFGFORCEMPS),
    .CFGINTERRUPTASSERTN (delay_CFGINTERRUPTASSERTN),
    .CFGINTERRUPTDI (delay_CFGINTERRUPTDI),
    .CFGINTERRUPTN (delay_CFGINTERRUPTN),
    .CFGINTERRUPTSTATN (delay_CFGINTERRUPTSTATN),
    .CFGMGMTBYTEENN (delay_CFGMGMTBYTEENN),
    .CFGMGMTDI (delay_CFGMGMTDI),
    .CFGMGMTDWADDR (delay_CFGMGMTDWADDR),
    .CFGMGMTRDENN (delay_CFGMGMTRDENN),
    .CFGMGMTWRENN (delay_CFGMGMTWRENN),
    .CFGMGMTWRREADONLYN (delay_CFGMGMTWRREADONLYN),
    .CFGMGMTWRRW1CASRWN (delay_CFGMGMTWRRW1CASRWN),
    .CFGPCIECAPINTERRUPTMSGNUM (delay_CFGPCIECAPINTERRUPTMSGNUM),
    .CFGPMFORCESTATE (delay_CFGPMFORCESTATE),
    .CFGPMFORCESTATEENN (delay_CFGPMFORCESTATEENN),
    .CFGPMHALTASPML0SN (delay_CFGPMHALTASPML0SN),
    .CFGPMHALTASPML1N (delay_CFGPMHALTASPML1N),
    .CFGPMSENDPMETON (delay_CFGPMSENDPMETON),
    .CFGPMTURNOFFOKN (delay_CFGPMTURNOFFOKN),
    .CFGPMWAKEN (delay_CFGPMWAKEN),
    .CFGPORTNUMBER (delay_CFGPORTNUMBER),
    .CFGREVID (delay_CFGREVID),
    .CFGSUBSYSID (delay_CFGSUBSYSID),
    .CFGSUBSYSVENDID (delay_CFGSUBSYSVENDID),
    .CFGTRNPENDINGN (delay_CFGTRNPENDINGN),
    .CFGVENDID (delay_CFGVENDID),
    .CMRSTN (delay_CMRSTN),
    .CMSTICKYRSTN (delay_CMSTICKYRSTN),
    .DBGMODE (delay_DBGMODE),
    .DBGSUBMODE (delay_DBGSUBMODE),
    .DLRSTN (delay_DLRSTN),
    .DRPADDR (delay_DRPADDR),
    .DRPCLK (delay_DRPCLK),
    .DRPDI (delay_DRPDI),
    .DRPEN (delay_DRPEN),
    .DRPWE (delay_DRPWE),
    .FUNCLVLRSTN (delay_FUNCLVLRSTN),
    .LL2SENDASREQL1 (delay_LL2SENDASREQL1),
    .LL2SENDENTERL1 (delay_LL2SENDENTERL1),
    .LL2SENDENTERL23 (delay_LL2SENDENTERL23),
    .LL2SENDPMACK (delay_LL2SENDPMACK),
    .LL2SUSPENDNOW (delay_LL2SUSPENDNOW),
    .LL2TLPRCV (delay_LL2TLPRCV),
    .MIMRXRDATA (delay_MIMRXRDATA),
    .MIMTXRDATA (delay_MIMTXRDATA),
    .PIPECLK (delay_PIPECLK),
    .PIPERX0CHANISALIGNED (delay_PIPERX0CHANISALIGNED),
    .PIPERX0CHARISK (delay_PIPERX0CHARISK),
    .PIPERX0DATA (delay_PIPERX0DATA),
    .PIPERX0ELECIDLE (delay_PIPERX0ELECIDLE),
    .PIPERX0PHYSTATUS (delay_PIPERX0PHYSTATUS),
    .PIPERX0STATUS (delay_PIPERX0STATUS),
    .PIPERX0VALID (delay_PIPERX0VALID),
    .PIPERX1CHANISALIGNED (delay_PIPERX1CHANISALIGNED),
    .PIPERX1CHARISK (delay_PIPERX1CHARISK),
    .PIPERX1DATA (delay_PIPERX1DATA),
    .PIPERX1ELECIDLE (delay_PIPERX1ELECIDLE),
    .PIPERX1PHYSTATUS (delay_PIPERX1PHYSTATUS),
    .PIPERX1STATUS (delay_PIPERX1STATUS),
    .PIPERX1VALID (delay_PIPERX1VALID),
    .PIPERX2CHANISALIGNED (delay_PIPERX2CHANISALIGNED),
    .PIPERX2CHARISK (delay_PIPERX2CHARISK),
    .PIPERX2DATA (delay_PIPERX2DATA),
    .PIPERX2ELECIDLE (delay_PIPERX2ELECIDLE),
    .PIPERX2PHYSTATUS (delay_PIPERX2PHYSTATUS),
    .PIPERX2STATUS (delay_PIPERX2STATUS),
    .PIPERX2VALID (delay_PIPERX2VALID),
    .PIPERX3CHANISALIGNED (delay_PIPERX3CHANISALIGNED),
    .PIPERX3CHARISK (delay_PIPERX3CHARISK),
    .PIPERX3DATA (delay_PIPERX3DATA),
    .PIPERX3ELECIDLE (delay_PIPERX3ELECIDLE),
    .PIPERX3PHYSTATUS (delay_PIPERX3PHYSTATUS),
    .PIPERX3STATUS (delay_PIPERX3STATUS),
    .PIPERX3VALID (delay_PIPERX3VALID),
    .PIPERX4CHANISALIGNED (delay_PIPERX4CHANISALIGNED),
    .PIPERX4CHARISK (delay_PIPERX4CHARISK),
    .PIPERX4DATA (delay_PIPERX4DATA),
    .PIPERX4ELECIDLE (delay_PIPERX4ELECIDLE),
    .PIPERX4PHYSTATUS (delay_PIPERX4PHYSTATUS),
    .PIPERX4STATUS (delay_PIPERX4STATUS),
    .PIPERX4VALID (delay_PIPERX4VALID),
    .PIPERX5CHANISALIGNED (delay_PIPERX5CHANISALIGNED),
    .PIPERX5CHARISK (delay_PIPERX5CHARISK),
    .PIPERX5DATA (delay_PIPERX5DATA),
    .PIPERX5ELECIDLE (delay_PIPERX5ELECIDLE),
    .PIPERX5PHYSTATUS (delay_PIPERX5PHYSTATUS),
    .PIPERX5STATUS (delay_PIPERX5STATUS),
    .PIPERX5VALID (delay_PIPERX5VALID),
    .PIPERX6CHANISALIGNED (delay_PIPERX6CHANISALIGNED),
    .PIPERX6CHARISK (delay_PIPERX6CHARISK),
    .PIPERX6DATA (delay_PIPERX6DATA),
    .PIPERX6ELECIDLE (delay_PIPERX6ELECIDLE),
    .PIPERX6PHYSTATUS (delay_PIPERX6PHYSTATUS),
    .PIPERX6STATUS (delay_PIPERX6STATUS),
    .PIPERX6VALID (delay_PIPERX6VALID),
    .PIPERX7CHANISALIGNED (delay_PIPERX7CHANISALIGNED),
    .PIPERX7CHARISK (delay_PIPERX7CHARISK),
    .PIPERX7DATA (delay_PIPERX7DATA),
    .PIPERX7ELECIDLE (delay_PIPERX7ELECIDLE),
    .PIPERX7PHYSTATUS (delay_PIPERX7PHYSTATUS),
    .PIPERX7STATUS (delay_PIPERX7STATUS),
    .PIPERX7VALID (delay_PIPERX7VALID),
    .PL2DIRECTEDLSTATE (delay_PL2DIRECTEDLSTATE),
    .PLDBGMODE (delay_PLDBGMODE),
    .PLDIRECTEDLINKAUTON (delay_PLDIRECTEDLINKAUTON),
    .PLDIRECTEDLINKCHANGE (delay_PLDIRECTEDLINKCHANGE),
    .PLDIRECTEDLINKSPEED (delay_PLDIRECTEDLINKSPEED),
    .PLDIRECTEDLINKWIDTH (delay_PLDIRECTEDLINKWIDTH),
    .PLDIRECTEDLTSSMNEW (delay_PLDIRECTEDLTSSMNEW),
    .PLDIRECTEDLTSSMNEWVLD (delay_PLDIRECTEDLTSSMNEWVLD),
    .PLDIRECTEDLTSSMSTALL (delay_PLDIRECTEDLTSSMSTALL),
    .PLDOWNSTREAMDEEMPHSOURCE (delay_PLDOWNSTREAMDEEMPHSOURCE),
    .PLRSTN (delay_PLRSTN),
    .PLTRANSMITHOTRST (delay_PLTRANSMITHOTRST),
    .PLUPSTREAMPREFERDEEMPH (delay_PLUPSTREAMPREFERDEEMPH),
    .SYSRSTN (delay_SYSRSTN),
    .TL2ASPMSUSPENDCREDITCHECK (delay_TL2ASPMSUSPENDCREDITCHECK),
    .TL2PPMSUSPENDREQ (delay_TL2PPMSUSPENDREQ),
    .TLRSTN (delay_TLRSTN),
    .TRNFCSEL (delay_TRNFCSEL),
    .TRNRDSTRDY (delay_TRNRDSTRDY),
    .TRNRFCPRET (delay_TRNRFCPRET),
    .TRNRNPOK (delay_TRNRNPOK),
    .TRNRNPREQ (delay_TRNRNPREQ),
    .TRNTCFGGNT (delay_TRNTCFGGNT),
    .TRNTD (delay_TRNTD),
    .TRNTDLLPDATA (delay_TRNTDLLPDATA),
    .TRNTDLLPSRCRDY (delay_TRNTDLLPSRCRDY),
    .TRNTECRCGEN (delay_TRNTECRCGEN),
    .TRNTEOF (delay_TRNTEOF),
    .TRNTERRFWD (delay_TRNTERRFWD),
    .TRNTREM (delay_TRNTREM),
    .TRNTSOF (delay_TRNTSOF),
    .TRNTSRCDSC (delay_TRNTSRCDSC),
    .TRNTSRCRDY (delay_TRNTSRCRDY),
    .TRNTSTR (delay_TRNTSTR),
    .USERCLK (delay_USERCLK),
    .USERCLK2 (delay_USERCLK2)
//    .GSR (GSR)
  );

  specify
`ifdef XIL_TIMING // Simprim
    $period (posedge DRPCLK, 0:0:0, notifier);
    $period (posedge PIPECLK, 0:0:0, notifier);
    $period (posedge USERCLK, 0:0:0, notifier);
    $period (posedge USERCLK2, 0:0:0, notifier);
    $setuphold (posedge DRPCLK, negedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, negedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, negedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, negedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, negedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, negedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, negedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, negedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, negedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, negedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, negedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, negedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, negedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, negedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, negedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, negedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, negedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, negedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, negedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge DRPCLK, posedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, posedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, posedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, posedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, posedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, posedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, posedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, posedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, posedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, posedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, posedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, posedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, posedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, posedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, posedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, posedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, posedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, posedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, posedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge PIPECLK, negedge PIPERX0CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX1CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX2CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX3CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX4CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX5CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX6CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6VALID);
    $setuphold (posedge PIPECLK, negedge PIPERX7CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHANISALIGNED);
    $setuphold (posedge PIPECLK, negedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge PIPECLK, negedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7VALID);
    $setuphold (posedge PIPECLK, negedge PLDBGMODE[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[0]);
    $setuphold (posedge PIPECLK, negedge PLDBGMODE[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[1]);
    $setuphold (posedge PIPECLK, negedge PLDBGMODE[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[2]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKAUTON, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKAUTON);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKCHANGE[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKCHANGE[0]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKCHANGE[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKCHANGE[1]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKSPEED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKSPEED);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKWIDTH[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKWIDTH[0]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLINKWIDTH[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKWIDTH[1]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEWVLD, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEWVLD);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[0]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[1]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[2]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[3]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[4]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMNEW[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[5]);
    $setuphold (posedge PIPECLK, negedge PLDIRECTEDLTSSMSTALL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMSTALL);
    $setuphold (posedge PIPECLK, negedge PLDOWNSTREAMDEEMPHSOURCE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDOWNSTREAMDEEMPHSOURCE);
    $setuphold (posedge PIPECLK, negedge PLRSTN, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLRSTN);
    $setuphold (posedge PIPECLK, negedge PLTRANSMITHOTRST, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLTRANSMITHOTRST);
    $setuphold (posedge PIPECLK, negedge PLUPSTREAMPREFERDEEMPH, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLUPSTREAMPREFERDEEMPH);
    $setuphold (posedge PIPECLK, posedge PIPERX0CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX1CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX2CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX3CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX4CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX5CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX6CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6VALID);
    $setuphold (posedge PIPECLK, posedge PIPERX7CHANISALIGNED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHANISALIGNED);
    $setuphold (posedge PIPECLK, posedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge PIPECLK, posedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7VALID);
    $setuphold (posedge PIPECLK, posedge PLDBGMODE[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[0]);
    $setuphold (posedge PIPECLK, posedge PLDBGMODE[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[1]);
    $setuphold (posedge PIPECLK, posedge PLDBGMODE[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDBGMODE[2]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKAUTON, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKAUTON);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKCHANGE[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKCHANGE[0]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKCHANGE[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKCHANGE[1]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKSPEED, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKSPEED);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKWIDTH[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKWIDTH[0]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLINKWIDTH[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLINKWIDTH[1]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEWVLD, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEWVLD);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[0]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[1]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[2]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[3]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[4]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMNEW[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMNEW[5]);
    $setuphold (posedge PIPECLK, posedge PLDIRECTEDLTSSMSTALL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDIRECTEDLTSSMSTALL);
    $setuphold (posedge PIPECLK, posedge PLDOWNSTREAMDEEMPHSOURCE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDOWNSTREAMDEEMPHSOURCE);
    $setuphold (posedge PIPECLK, posedge PLRSTN, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLRSTN);
    $setuphold (posedge PIPECLK, posedge PLTRANSMITHOTRST, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLTRANSMITHOTRST);
    $setuphold (posedge PIPECLK, posedge PLUPSTREAMPREFERDEEMPH, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLUPSTREAMPREFERDEEMPH);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[0]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[10]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[11]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[12]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[13]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[14]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[15]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[16]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[17]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[18]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[19]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[1]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[20]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[21]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[22]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[23]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[24]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[25]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[26]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[27]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[28]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[29]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[2]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[30]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[31]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[32]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[33]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[34]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[35]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[36]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[37]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[38]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[39]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[3]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[40]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[41]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[42]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[43]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[44]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[45]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[46]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[47]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[48]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[49]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[4]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[50]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[51]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[52]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[53]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[54]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[55]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[56]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[57]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[58]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[59]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[5]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[60]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[61]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[62]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[63]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[64]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[65]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[66]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[67]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[6]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[7]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[8]);
    $setuphold (posedge USERCLK, negedge MIMRXRDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[9]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[0]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[10]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[11]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[12]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[13]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[14]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[15]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[16]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[17]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[18]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[19]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[1]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[20]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[21]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[22]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[23]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[24]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[25]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[26]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[27]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[28]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[29]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[2]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[30]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[31]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[32]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[33]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[34]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[35]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[36]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[37]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[38]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[39]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[3]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[40]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[41]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[42]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[43]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[44]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[45]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[46]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[47]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[48]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[49]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[4]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[50]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[51]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[52]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[53]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[54]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[55]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[56]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[57]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[58]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[59]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[5]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[60]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[61]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[62]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[63]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[64]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[65]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[66]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[67]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[68]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[6]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[7]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[8]);
    $setuphold (posedge USERCLK, negedge MIMTXRDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[9]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[0]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[10]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[11]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[12]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[13]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[14]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[15]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[16]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[17]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[18]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[19]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[1]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[20]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[21]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[22]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[23]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[24]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[25]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[26]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[27]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[28]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[29]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[2]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[30]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[31]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[32]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[33]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[34]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[35]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[36]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[37]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[38]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[39]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[3]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[40]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[41]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[42]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[43]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[44]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[45]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[46]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[47]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[48]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[49]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[4]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[50]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[51]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[52]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[53]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[54]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[55]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[56]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[57]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[58]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[59]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[5]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[60]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[61]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[62]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[63]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[64]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[65]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[66]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[67]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[6]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[7]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[8]);
    $setuphold (posedge USERCLK, posedge MIMRXRDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMRXRDATA[9]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[0]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[10]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[11]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[12]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[13]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[14]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[15]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[16]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[17]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[18]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[19]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[1]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[20]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[21]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[22]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[23]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[24]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[25]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[26]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[27]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[28]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[29]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[2]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[30]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[31]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[32]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[33]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[34]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[35]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[36]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[37]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[38]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[39]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[3]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[40]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[41]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[42]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[43]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[44]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[45]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[46]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[47]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[48]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[49]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[4]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[50]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[51]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[52]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[53]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[54]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[55]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[56]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[57]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[58]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[59]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[5]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[60]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[61]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[62]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[63]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[64]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[65]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[66]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[67]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[68]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[6]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[7]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[8]);
    $setuphold (posedge USERCLK, posedge MIMTXRDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MIMTXRDATA[9]);
    $setuphold (posedge USERCLK2, negedge CFGAERINTERRUPTMSGNUM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[0]);
    $setuphold (posedge USERCLK2, negedge CFGAERINTERRUPTMSGNUM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[1]);
    $setuphold (posedge USERCLK2, negedge CFGAERINTERRUPTMSGNUM[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[2]);
    $setuphold (posedge USERCLK2, negedge CFGAERINTERRUPTMSGNUM[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[3]);
    $setuphold (posedge USERCLK2, negedge CFGAERINTERRUPTMSGNUM[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[4]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK2, negedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK2, negedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK2, negedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK2, negedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK2, negedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK2, negedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK2, negedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK2, negedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK2, negedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK2, negedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK2, negedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK2, negedge CFGERRACSN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRACSN);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[0]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[100]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[101]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[102]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[103]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[104]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[105]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[106]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[107]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[108]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[109]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[10]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[110]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[111]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[112]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[113]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[114]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[115]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[116]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[117]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[118]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[119]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[11]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[120]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[121]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[122]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[123]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[124]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[125]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[126]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[127]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[12]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[13]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[14]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[15]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[16]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[17]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[18]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[19]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[1]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[20]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[21]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[22]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[23]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[24]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[25]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[26]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[27]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[28]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[29]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[2]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[30]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[31]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[32]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[33]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[34]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[35]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[36]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[37]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[38]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[39]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[3]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[40]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[41]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[42]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[43]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[44]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[45]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[46]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[47]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[48]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[49]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[4]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[50]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[51]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[52]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[53]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[54]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[55]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[56]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[57]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[58]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[59]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[5]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[60]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[61]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[62]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[63]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[64]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[65]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[66]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[67]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[68]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[69]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[6]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[70]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[71]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[72]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[73]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[74]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[75]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[76]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[77]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[78]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[79]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[7]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[80]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[81]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[82]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[83]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[84]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[85]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[86]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[87]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[88]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[89]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[8]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[90]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[91]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[92]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[93]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[94]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[95]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[96]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[97]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[98]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[99]);
    $setuphold (posedge USERCLK2, negedge CFGERRAERHEADERLOG[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[9]);
    $setuphold (posedge USERCLK2, negedge CFGERRATOMICEGRESSBLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRATOMICEGRESSBLOCKEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCORN);
    $setuphold (posedge USERCLK2, negedge CFGERRCPLABORTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLABORTN);
    $setuphold (posedge USERCLK2, negedge CFGERRCPLTIMEOUTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLTIMEOUTN);
    $setuphold (posedge USERCLK2, negedge CFGERRCPLUNEXPECTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLUNEXPECTN);
    $setuphold (posedge USERCLK2, negedge CFGERRECRCN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRECRCN);
    $setuphold (posedge USERCLK2, negedge CFGERRINTERNALCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRINTERNALCORN);
    $setuphold (posedge USERCLK2, negedge CFGERRINTERNALUNCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRINTERNALUNCORN);
    $setuphold (posedge USERCLK2, negedge CFGERRLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRLOCKEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRMALFORMEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRMALFORMEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRMCBLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRMCBLOCKEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRNORECOVERYN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRNORECOVERYN);
    $setuphold (posedge USERCLK2, negedge CFGERRPOISONEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRPOISONEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRPOSTEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRPOSTEDN);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[0]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[10]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[11]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[12]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[13]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[14]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[15]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[16]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[17]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[18]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[19]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[1]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[20]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[21]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[22]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[23]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[24]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[25]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[26]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[27]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[28]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[29]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[2]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[30]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[31]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[32]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[33]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[34]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[35]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[36]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[37]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[38]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[39]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[3]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[40]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[41]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[42]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[43]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[44]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[45]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[46]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[47]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[4]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[5]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[6]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[7]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[8]);
    $setuphold (posedge USERCLK2, negedge CFGERRTLPCPLHEADER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[9]);
    $setuphold (posedge USERCLK2, negedge CFGERRURN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRURN);
    $setuphold (posedge USERCLK2, negedge CFGFORCECOMMONCLOCKOFF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCECOMMONCLOCKOFF);
    $setuphold (posedge USERCLK2, negedge CFGFORCEEXTENDEDSYNCON, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEEXTENDEDSYNCON);
    $setuphold (posedge USERCLK2, negedge CFGFORCEMPS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[0]);
    $setuphold (posedge USERCLK2, negedge CFGFORCEMPS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[1]);
    $setuphold (posedge USERCLK2, negedge CFGFORCEMPS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[2]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTASSERTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTASSERTN);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[0]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[1]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[2]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[3]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[4]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[5]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[6]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTDI[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[7]);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTN);
    $setuphold (posedge USERCLK2, negedge CFGINTERRUPTSTATN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTSTATN);
    $setuphold (posedge USERCLK2, negedge CFGMGMTBYTEENN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[0]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTBYTEENN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[1]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTBYTEENN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[2]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTBYTEENN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[3]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[0]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[10]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[11]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[12]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[13]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[14]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[15]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[16]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[17]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[18]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[19]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[1]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[20]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[21]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[22]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[23]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[24]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[25]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[26]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[27]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[28]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[29]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[2]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[30]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[31]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[3]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[4]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[5]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[6]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[7]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[8]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDI[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[9]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[0]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[1]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[2]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[3]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[4]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[5]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[6]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[7]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[8]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTDWADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[9]);
    $setuphold (posedge USERCLK2, negedge CFGMGMTRDENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTRDENN);
    $setuphold (posedge USERCLK2, negedge CFGMGMTWRENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRENN);
    $setuphold (posedge USERCLK2, negedge CFGMGMTWRREADONLYN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRREADONLYN);
    $setuphold (posedge USERCLK2, negedge CFGMGMTWRRW1CASRWN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRRW1CASRWN);
    $setuphold (posedge USERCLK2, negedge CFGPCIECAPINTERRUPTMSGNUM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[0]);
    $setuphold (posedge USERCLK2, negedge CFGPCIECAPINTERRUPTMSGNUM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[1]);
    $setuphold (posedge USERCLK2, negedge CFGPCIECAPINTERRUPTMSGNUM[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[2]);
    $setuphold (posedge USERCLK2, negedge CFGPCIECAPINTERRUPTMSGNUM[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[3]);
    $setuphold (posedge USERCLK2, negedge CFGPCIECAPINTERRUPTMSGNUM[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[4]);
    $setuphold (posedge USERCLK2, negedge CFGPMFORCESTATEENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATEENN);
    $setuphold (posedge USERCLK2, negedge CFGPMFORCESTATE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATE[0]);
    $setuphold (posedge USERCLK2, negedge CFGPMFORCESTATE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATE[1]);
    $setuphold (posedge USERCLK2, negedge CFGPMHALTASPML0SN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMHALTASPML0SN);
    $setuphold (posedge USERCLK2, negedge CFGPMHALTASPML1N, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMHALTASPML1N);
    $setuphold (posedge USERCLK2, negedge CFGPMSENDPMETON, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMSENDPMETON);
    $setuphold (posedge USERCLK2, negedge CFGPMTURNOFFOKN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMTURNOFFOKN);
    $setuphold (posedge USERCLK2, negedge CFGPMWAKEN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMWAKEN);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[0]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[1]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[2]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[3]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[4]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[5]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[6]);
    $setuphold (posedge USERCLK2, negedge CFGPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[7]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK2, negedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK2, negedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK2, negedge CFGTRNPENDINGN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGTRNPENDINGN);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK2, negedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK2, negedge CMRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CMRSTN);
    $setuphold (posedge USERCLK2, negedge CMSTICKYRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CMSTICKYRSTN);
    $setuphold (posedge USERCLK2, negedge DBGMODE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGMODE[0]);
    $setuphold (posedge USERCLK2, negedge DBGMODE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGMODE[1]);
    $setuphold (posedge USERCLK2, negedge DBGSUBMODE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGSUBMODE);
    $setuphold (posedge USERCLK2, negedge DLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DLRSTN);
    $setuphold (posedge USERCLK2, negedge FUNCLVLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_FUNCLVLRSTN);
    $setuphold (posedge USERCLK2, negedge LL2SENDASREQL1, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDASREQL1);
    $setuphold (posedge USERCLK2, negedge LL2SENDENTERL1, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDENTERL1);
    $setuphold (posedge USERCLK2, negedge LL2SENDENTERL23, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDENTERL23);
    $setuphold (posedge USERCLK2, negedge LL2SENDPMACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDPMACK);
    $setuphold (posedge USERCLK2, negedge LL2SUSPENDNOW, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SUSPENDNOW);
    $setuphold (posedge USERCLK2, negedge LL2TLPRCV, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2TLPRCV);
    $setuphold (posedge USERCLK2, negedge PL2DIRECTEDLSTATE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[0]);
    $setuphold (posedge USERCLK2, negedge PL2DIRECTEDLSTATE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[1]);
    $setuphold (posedge USERCLK2, negedge PL2DIRECTEDLSTATE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[2]);
    $setuphold (posedge USERCLK2, negedge PL2DIRECTEDLSTATE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[3]);
    $setuphold (posedge USERCLK2, negedge PL2DIRECTEDLSTATE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[4]);
    $setuphold (posedge USERCLK2, negedge TL2ASPMSUSPENDCREDITCHECK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TL2ASPMSUSPENDCREDITCHECK);
    $setuphold (posedge USERCLK2, negedge TL2PPMSUSPENDREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TL2PPMSUSPENDREQ);
    $setuphold (posedge USERCLK2, negedge TLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TLRSTN);
    $setuphold (posedge USERCLK2, negedge TRNFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[0]);
    $setuphold (posedge USERCLK2, negedge TRNFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[1]);
    $setuphold (posedge USERCLK2, negedge TRNFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[2]);
    $setuphold (posedge USERCLK2, negedge TRNRDSTRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRDSTRDY);
    $setuphold (posedge USERCLK2, negedge TRNRFCPRET, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRFCPRET);
    $setuphold (posedge USERCLK2, negedge TRNRNPOK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRNPOK);
    $setuphold (posedge USERCLK2, negedge TRNRNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRNPREQ);
    $setuphold (posedge USERCLK2, negedge TRNTCFGGNT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTCFGGNT);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[0]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[10]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[11]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[12]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[13]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[14]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[15]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[16]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[17]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[18]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[19]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[1]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[20]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[21]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[22]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[23]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[24]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[25]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[26]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[27]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[28]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[29]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[2]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[30]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[31]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[3]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[4]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[5]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[6]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[7]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[8]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[9]);
    $setuphold (posedge USERCLK2, negedge TRNTDLLPSRCRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPSRCRDY);
    $setuphold (posedge USERCLK2, negedge TRNTD[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[0]);
    $setuphold (posedge USERCLK2, negedge TRNTD[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[100]);
    $setuphold (posedge USERCLK2, negedge TRNTD[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[101]);
    $setuphold (posedge USERCLK2, negedge TRNTD[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[102]);
    $setuphold (posedge USERCLK2, negedge TRNTD[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[103]);
    $setuphold (posedge USERCLK2, negedge TRNTD[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[104]);
    $setuphold (posedge USERCLK2, negedge TRNTD[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[105]);
    $setuphold (posedge USERCLK2, negedge TRNTD[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[106]);
    $setuphold (posedge USERCLK2, negedge TRNTD[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[107]);
    $setuphold (posedge USERCLK2, negedge TRNTD[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[108]);
    $setuphold (posedge USERCLK2, negedge TRNTD[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[109]);
    $setuphold (posedge USERCLK2, negedge TRNTD[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[10]);
    $setuphold (posedge USERCLK2, negedge TRNTD[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[110]);
    $setuphold (posedge USERCLK2, negedge TRNTD[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[111]);
    $setuphold (posedge USERCLK2, negedge TRNTD[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[112]);
    $setuphold (posedge USERCLK2, negedge TRNTD[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[113]);
    $setuphold (posedge USERCLK2, negedge TRNTD[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[114]);
    $setuphold (posedge USERCLK2, negedge TRNTD[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[115]);
    $setuphold (posedge USERCLK2, negedge TRNTD[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[116]);
    $setuphold (posedge USERCLK2, negedge TRNTD[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[117]);
    $setuphold (posedge USERCLK2, negedge TRNTD[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[118]);
    $setuphold (posedge USERCLK2, negedge TRNTD[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[119]);
    $setuphold (posedge USERCLK2, negedge TRNTD[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[11]);
    $setuphold (posedge USERCLK2, negedge TRNTD[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[120]);
    $setuphold (posedge USERCLK2, negedge TRNTD[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[121]);
    $setuphold (posedge USERCLK2, negedge TRNTD[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[122]);
    $setuphold (posedge USERCLK2, negedge TRNTD[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[123]);
    $setuphold (posedge USERCLK2, negedge TRNTD[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[124]);
    $setuphold (posedge USERCLK2, negedge TRNTD[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[125]);
    $setuphold (posedge USERCLK2, negedge TRNTD[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[126]);
    $setuphold (posedge USERCLK2, negedge TRNTD[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[127]);
    $setuphold (posedge USERCLK2, negedge TRNTD[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[12]);
    $setuphold (posedge USERCLK2, negedge TRNTD[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[13]);
    $setuphold (posedge USERCLK2, negedge TRNTD[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[14]);
    $setuphold (posedge USERCLK2, negedge TRNTD[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[15]);
    $setuphold (posedge USERCLK2, negedge TRNTD[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[16]);
    $setuphold (posedge USERCLK2, negedge TRNTD[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[17]);
    $setuphold (posedge USERCLK2, negedge TRNTD[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[18]);
    $setuphold (posedge USERCLK2, negedge TRNTD[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[19]);
    $setuphold (posedge USERCLK2, negedge TRNTD[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[1]);
    $setuphold (posedge USERCLK2, negedge TRNTD[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[20]);
    $setuphold (posedge USERCLK2, negedge TRNTD[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[21]);
    $setuphold (posedge USERCLK2, negedge TRNTD[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[22]);
    $setuphold (posedge USERCLK2, negedge TRNTD[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[23]);
    $setuphold (posedge USERCLK2, negedge TRNTD[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[24]);
    $setuphold (posedge USERCLK2, negedge TRNTD[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[25]);
    $setuphold (posedge USERCLK2, negedge TRNTD[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[26]);
    $setuphold (posedge USERCLK2, negedge TRNTD[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[27]);
    $setuphold (posedge USERCLK2, negedge TRNTD[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[28]);
    $setuphold (posedge USERCLK2, negedge TRNTD[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[29]);
    $setuphold (posedge USERCLK2, negedge TRNTD[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[2]);
    $setuphold (posedge USERCLK2, negedge TRNTD[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[30]);
    $setuphold (posedge USERCLK2, negedge TRNTD[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[31]);
    $setuphold (posedge USERCLK2, negedge TRNTD[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[32]);
    $setuphold (posedge USERCLK2, negedge TRNTD[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[33]);
    $setuphold (posedge USERCLK2, negedge TRNTD[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[34]);
    $setuphold (posedge USERCLK2, negedge TRNTD[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[35]);
    $setuphold (posedge USERCLK2, negedge TRNTD[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[36]);
    $setuphold (posedge USERCLK2, negedge TRNTD[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[37]);
    $setuphold (posedge USERCLK2, negedge TRNTD[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[38]);
    $setuphold (posedge USERCLK2, negedge TRNTD[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[39]);
    $setuphold (posedge USERCLK2, negedge TRNTD[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[3]);
    $setuphold (posedge USERCLK2, negedge TRNTD[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[40]);
    $setuphold (posedge USERCLK2, negedge TRNTD[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[41]);
    $setuphold (posedge USERCLK2, negedge TRNTD[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[42]);
    $setuphold (posedge USERCLK2, negedge TRNTD[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[43]);
    $setuphold (posedge USERCLK2, negedge TRNTD[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[44]);
    $setuphold (posedge USERCLK2, negedge TRNTD[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[45]);
    $setuphold (posedge USERCLK2, negedge TRNTD[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[46]);
    $setuphold (posedge USERCLK2, negedge TRNTD[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[47]);
    $setuphold (posedge USERCLK2, negedge TRNTD[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[48]);
    $setuphold (posedge USERCLK2, negedge TRNTD[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[49]);
    $setuphold (posedge USERCLK2, negedge TRNTD[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[4]);
    $setuphold (posedge USERCLK2, negedge TRNTD[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[50]);
    $setuphold (posedge USERCLK2, negedge TRNTD[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[51]);
    $setuphold (posedge USERCLK2, negedge TRNTD[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[52]);
    $setuphold (posedge USERCLK2, negedge TRNTD[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[53]);
    $setuphold (posedge USERCLK2, negedge TRNTD[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[54]);
    $setuphold (posedge USERCLK2, negedge TRNTD[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[55]);
    $setuphold (posedge USERCLK2, negedge TRNTD[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[56]);
    $setuphold (posedge USERCLK2, negedge TRNTD[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[57]);
    $setuphold (posedge USERCLK2, negedge TRNTD[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[58]);
    $setuphold (posedge USERCLK2, negedge TRNTD[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[59]);
    $setuphold (posedge USERCLK2, negedge TRNTD[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[5]);
    $setuphold (posedge USERCLK2, negedge TRNTD[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[60]);
    $setuphold (posedge USERCLK2, negedge TRNTD[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[61]);
    $setuphold (posedge USERCLK2, negedge TRNTD[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[62]);
    $setuphold (posedge USERCLK2, negedge TRNTD[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[63]);
    $setuphold (posedge USERCLK2, negedge TRNTD[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[64]);
    $setuphold (posedge USERCLK2, negedge TRNTD[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[65]);
    $setuphold (posedge USERCLK2, negedge TRNTD[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[66]);
    $setuphold (posedge USERCLK2, negedge TRNTD[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[67]);
    $setuphold (posedge USERCLK2, negedge TRNTD[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[68]);
    $setuphold (posedge USERCLK2, negedge TRNTD[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[69]);
    $setuphold (posedge USERCLK2, negedge TRNTD[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[6]);
    $setuphold (posedge USERCLK2, negedge TRNTD[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[70]);
    $setuphold (posedge USERCLK2, negedge TRNTD[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[71]);
    $setuphold (posedge USERCLK2, negedge TRNTD[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[72]);
    $setuphold (posedge USERCLK2, negedge TRNTD[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[73]);
    $setuphold (posedge USERCLK2, negedge TRNTD[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[74]);
    $setuphold (posedge USERCLK2, negedge TRNTD[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[75]);
    $setuphold (posedge USERCLK2, negedge TRNTD[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[76]);
    $setuphold (posedge USERCLK2, negedge TRNTD[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[77]);
    $setuphold (posedge USERCLK2, negedge TRNTD[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[78]);
    $setuphold (posedge USERCLK2, negedge TRNTD[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[79]);
    $setuphold (posedge USERCLK2, negedge TRNTD[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[7]);
    $setuphold (posedge USERCLK2, negedge TRNTD[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[80]);
    $setuphold (posedge USERCLK2, negedge TRNTD[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[81]);
    $setuphold (posedge USERCLK2, negedge TRNTD[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[82]);
    $setuphold (posedge USERCLK2, negedge TRNTD[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[83]);
    $setuphold (posedge USERCLK2, negedge TRNTD[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[84]);
    $setuphold (posedge USERCLK2, negedge TRNTD[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[85]);
    $setuphold (posedge USERCLK2, negedge TRNTD[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[86]);
    $setuphold (posedge USERCLK2, negedge TRNTD[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[87]);
    $setuphold (posedge USERCLK2, negedge TRNTD[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[88]);
    $setuphold (posedge USERCLK2, negedge TRNTD[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[89]);
    $setuphold (posedge USERCLK2, negedge TRNTD[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[8]);
    $setuphold (posedge USERCLK2, negedge TRNTD[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[90]);
    $setuphold (posedge USERCLK2, negedge TRNTD[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[91]);
    $setuphold (posedge USERCLK2, negedge TRNTD[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[92]);
    $setuphold (posedge USERCLK2, negedge TRNTD[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[93]);
    $setuphold (posedge USERCLK2, negedge TRNTD[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[94]);
    $setuphold (posedge USERCLK2, negedge TRNTD[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[95]);
    $setuphold (posedge USERCLK2, negedge TRNTD[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[96]);
    $setuphold (posedge USERCLK2, negedge TRNTD[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[97]);
    $setuphold (posedge USERCLK2, negedge TRNTD[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[98]);
    $setuphold (posedge USERCLK2, negedge TRNTD[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[99]);
    $setuphold (posedge USERCLK2, negedge TRNTD[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[9]);
    $setuphold (posedge USERCLK2, negedge TRNTECRCGEN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTECRCGEN);
    $setuphold (posedge USERCLK2, negedge TRNTEOF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTEOF);
    $setuphold (posedge USERCLK2, negedge TRNTERRFWD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTERRFWD);
    $setuphold (posedge USERCLK2, negedge TRNTREM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTREM[0]);
    $setuphold (posedge USERCLK2, negedge TRNTREM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTREM[1]);
    $setuphold (posedge USERCLK2, negedge TRNTSOF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSOF);
    $setuphold (posedge USERCLK2, negedge TRNTSRCDSC, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSRCDSC);
    $setuphold (posedge USERCLK2, negedge TRNTSRCRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSRCRDY);
    $setuphold (posedge USERCLK2, negedge TRNTSTR, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSTR);
    $setuphold (posedge USERCLK2, posedge CFGAERINTERRUPTMSGNUM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[0]);
    $setuphold (posedge USERCLK2, posedge CFGAERINTERRUPTMSGNUM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[1]);
    $setuphold (posedge USERCLK2, posedge CFGAERINTERRUPTMSGNUM[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[2]);
    $setuphold (posedge USERCLK2, posedge CFGAERINTERRUPTMSGNUM[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[3]);
    $setuphold (posedge USERCLK2, posedge CFGAERINTERRUPTMSGNUM[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGAERINTERRUPTMSGNUM[4]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK2, posedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK2, posedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK2, posedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK2, posedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK2, posedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK2, posedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK2, posedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK2, posedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK2, posedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK2, posedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK2, posedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK2, posedge CFGERRACSN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRACSN);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[0]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[100]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[101]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[102]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[103]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[104]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[105]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[106]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[107]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[108]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[109]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[10]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[110]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[111]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[112]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[113]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[114]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[115]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[116]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[117]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[118]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[119]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[11]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[120]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[121]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[122]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[123]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[124]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[125]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[126]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[127]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[12]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[13]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[14]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[15]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[16]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[17]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[18]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[19]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[1]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[20]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[21]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[22]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[23]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[24]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[25]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[26]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[27]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[28]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[29]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[2]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[30]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[31]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[32]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[33]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[34]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[35]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[36]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[37]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[38]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[39]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[3]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[40]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[41]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[42]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[43]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[44]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[45]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[46]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[47]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[48]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[49]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[4]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[50]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[51]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[52]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[53]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[54]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[55]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[56]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[57]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[58]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[59]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[5]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[60]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[61]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[62]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[63]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[64]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[65]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[66]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[67]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[68]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[69]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[6]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[70]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[71]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[72]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[73]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[74]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[75]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[76]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[77]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[78]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[79]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[7]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[80]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[81]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[82]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[83]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[84]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[85]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[86]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[87]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[88]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[89]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[8]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[90]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[91]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[92]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[93]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[94]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[95]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[96]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[97]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[98]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[99]);
    $setuphold (posedge USERCLK2, posedge CFGERRAERHEADERLOG[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRAERHEADERLOG[9]);
    $setuphold (posedge USERCLK2, posedge CFGERRATOMICEGRESSBLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRATOMICEGRESSBLOCKEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCORN);
    $setuphold (posedge USERCLK2, posedge CFGERRCPLABORTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLABORTN);
    $setuphold (posedge USERCLK2, posedge CFGERRCPLTIMEOUTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLTIMEOUTN);
    $setuphold (posedge USERCLK2, posedge CFGERRCPLUNEXPECTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRCPLUNEXPECTN);
    $setuphold (posedge USERCLK2, posedge CFGERRECRCN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRECRCN);
    $setuphold (posedge USERCLK2, posedge CFGERRINTERNALCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRINTERNALCORN);
    $setuphold (posedge USERCLK2, posedge CFGERRINTERNALUNCORN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRINTERNALUNCORN);
    $setuphold (posedge USERCLK2, posedge CFGERRLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRLOCKEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRMALFORMEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRMALFORMEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRMCBLOCKEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRMCBLOCKEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRNORECOVERYN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRNORECOVERYN);
    $setuphold (posedge USERCLK2, posedge CFGERRPOISONEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRPOISONEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRPOSTEDN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRPOSTEDN);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[0]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[10]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[11]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[12]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[13]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[14]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[15]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[16]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[17]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[18]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[19]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[1]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[20]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[21]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[22]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[23]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[24]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[25]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[26]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[27]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[28]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[29]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[2]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[30]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[31]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[32]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[33]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[34]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[35]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[36]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[37]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[38]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[39]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[3]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[40]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[41]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[42]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[43]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[44]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[45]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[46]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[47]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[4]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[5]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[6]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[7]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[8]);
    $setuphold (posedge USERCLK2, posedge CFGERRTLPCPLHEADER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRTLPCPLHEADER[9]);
    $setuphold (posedge USERCLK2, posedge CFGERRURN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGERRURN);
    $setuphold (posedge USERCLK2, posedge CFGFORCECOMMONCLOCKOFF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCECOMMONCLOCKOFF);
    $setuphold (posedge USERCLK2, posedge CFGFORCEEXTENDEDSYNCON, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEEXTENDEDSYNCON);
    $setuphold (posedge USERCLK2, posedge CFGFORCEMPS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[0]);
    $setuphold (posedge USERCLK2, posedge CFGFORCEMPS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[1]);
    $setuphold (posedge USERCLK2, posedge CFGFORCEMPS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGFORCEMPS[2]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTASSERTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTASSERTN);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[0]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[1]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[2]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[3]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[4]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[5]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[6]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTDI[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTDI[7]);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTN);
    $setuphold (posedge USERCLK2, posedge CFGINTERRUPTSTATN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGINTERRUPTSTATN);
    $setuphold (posedge USERCLK2, posedge CFGMGMTBYTEENN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[0]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTBYTEENN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[1]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTBYTEENN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[2]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTBYTEENN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTBYTEENN[3]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[0]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[10]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[11]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[12]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[13]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[14]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[15]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[16]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[17]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[18]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[19]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[1]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[20]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[21]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[22]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[23]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[24]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[25]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[26]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[27]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[28]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[29]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[2]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[30]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[31]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[3]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[4]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[5]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[6]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[7]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[8]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDI[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDI[9]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[0]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[1]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[2]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[3]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[4]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[5]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[6]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[7]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[8]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTDWADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTDWADDR[9]);
    $setuphold (posedge USERCLK2, posedge CFGMGMTRDENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTRDENN);
    $setuphold (posedge USERCLK2, posedge CFGMGMTWRENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRENN);
    $setuphold (posedge USERCLK2, posedge CFGMGMTWRREADONLYN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRREADONLYN);
    $setuphold (posedge USERCLK2, posedge CFGMGMTWRRW1CASRWN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGMGMTWRRW1CASRWN);
    $setuphold (posedge USERCLK2, posedge CFGPCIECAPINTERRUPTMSGNUM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[0]);
    $setuphold (posedge USERCLK2, posedge CFGPCIECAPINTERRUPTMSGNUM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[1]);
    $setuphold (posedge USERCLK2, posedge CFGPCIECAPINTERRUPTMSGNUM[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[2]);
    $setuphold (posedge USERCLK2, posedge CFGPCIECAPINTERRUPTMSGNUM[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[3]);
    $setuphold (posedge USERCLK2, posedge CFGPCIECAPINTERRUPTMSGNUM[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPCIECAPINTERRUPTMSGNUM[4]);
    $setuphold (posedge USERCLK2, posedge CFGPMFORCESTATEENN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATEENN);
    $setuphold (posedge USERCLK2, posedge CFGPMFORCESTATE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATE[0]);
    $setuphold (posedge USERCLK2, posedge CFGPMFORCESTATE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMFORCESTATE[1]);
    $setuphold (posedge USERCLK2, posedge CFGPMHALTASPML0SN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMHALTASPML0SN);
    $setuphold (posedge USERCLK2, posedge CFGPMHALTASPML1N, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMHALTASPML1N);
    $setuphold (posedge USERCLK2, posedge CFGPMSENDPMETON, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMSENDPMETON);
    $setuphold (posedge USERCLK2, posedge CFGPMTURNOFFOKN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMTURNOFFOKN);
    $setuphold (posedge USERCLK2, posedge CFGPMWAKEN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPMWAKEN);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[0]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[1]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[2]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[3]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[4]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[5]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[6]);
    $setuphold (posedge USERCLK2, posedge CFGPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGPORTNUMBER[7]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK2, posedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK2, posedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK2, posedge CFGTRNPENDINGN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGTRNPENDINGN);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK2, posedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK2, posedge CMRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CMRSTN);
    $setuphold (posedge USERCLK2, posedge CMSTICKYRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_CMSTICKYRSTN);
    $setuphold (posedge USERCLK2, posedge DBGMODE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGMODE[0]);
    $setuphold (posedge USERCLK2, posedge DBGMODE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGMODE[1]);
    $setuphold (posedge USERCLK2, posedge DBGSUBMODE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DBGSUBMODE);
    $setuphold (posedge USERCLK2, posedge DLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_DLRSTN);
    $setuphold (posedge USERCLK2, posedge FUNCLVLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_FUNCLVLRSTN);
    $setuphold (posedge USERCLK2, posedge LL2SENDASREQL1, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDASREQL1);
    $setuphold (posedge USERCLK2, posedge LL2SENDENTERL1, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDENTERL1);
    $setuphold (posedge USERCLK2, posedge LL2SENDENTERL23, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDENTERL23);
    $setuphold (posedge USERCLK2, posedge LL2SENDPMACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SENDPMACK);
    $setuphold (posedge USERCLK2, posedge LL2SUSPENDNOW, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2SUSPENDNOW);
    $setuphold (posedge USERCLK2, posedge LL2TLPRCV, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_LL2TLPRCV);
    $setuphold (posedge USERCLK2, posedge PL2DIRECTEDLSTATE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[0]);
    $setuphold (posedge USERCLK2, posedge PL2DIRECTEDLSTATE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[1]);
    $setuphold (posedge USERCLK2, posedge PL2DIRECTEDLSTATE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[2]);
    $setuphold (posedge USERCLK2, posedge PL2DIRECTEDLSTATE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[3]);
    $setuphold (posedge USERCLK2, posedge PL2DIRECTEDLSTATE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_PL2DIRECTEDLSTATE[4]);
    $setuphold (posedge USERCLK2, posedge TL2ASPMSUSPENDCREDITCHECK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TL2ASPMSUSPENDCREDITCHECK);
    $setuphold (posedge USERCLK2, posedge TL2PPMSUSPENDREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TL2PPMSUSPENDREQ);
    $setuphold (posedge USERCLK2, posedge TLRSTN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TLRSTN);
    $setuphold (posedge USERCLK2, posedge TRNFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[0]);
    $setuphold (posedge USERCLK2, posedge TRNFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[1]);
    $setuphold (posedge USERCLK2, posedge TRNFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNFCSEL[2]);
    $setuphold (posedge USERCLK2, posedge TRNRDSTRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRDSTRDY);
    $setuphold (posedge USERCLK2, posedge TRNRFCPRET, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRFCPRET);
    $setuphold (posedge USERCLK2, posedge TRNRNPOK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRNPOK);
    $setuphold (posedge USERCLK2, posedge TRNRNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNRNPREQ);
    $setuphold (posedge USERCLK2, posedge TRNTCFGGNT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTCFGGNT);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[0]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[10]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[11]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[12]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[13]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[14]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[15]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[16]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[17]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[18]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[19]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[1]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[20]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[21]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[22]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[23]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[24]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[25]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[26]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[27]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[28]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[29]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[2]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[30]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[31]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[3]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[4]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[5]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[6]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[7]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[8]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPDATA[9]);
    $setuphold (posedge USERCLK2, posedge TRNTDLLPSRCRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTDLLPSRCRDY);
    $setuphold (posedge USERCLK2, posedge TRNTD[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[0]);
    $setuphold (posedge USERCLK2, posedge TRNTD[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[100]);
    $setuphold (posedge USERCLK2, posedge TRNTD[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[101]);
    $setuphold (posedge USERCLK2, posedge TRNTD[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[102]);
    $setuphold (posedge USERCLK2, posedge TRNTD[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[103]);
    $setuphold (posedge USERCLK2, posedge TRNTD[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[104]);
    $setuphold (posedge USERCLK2, posedge TRNTD[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[105]);
    $setuphold (posedge USERCLK2, posedge TRNTD[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[106]);
    $setuphold (posedge USERCLK2, posedge TRNTD[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[107]);
    $setuphold (posedge USERCLK2, posedge TRNTD[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[108]);
    $setuphold (posedge USERCLK2, posedge TRNTD[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[109]);
    $setuphold (posedge USERCLK2, posedge TRNTD[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[10]);
    $setuphold (posedge USERCLK2, posedge TRNTD[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[110]);
    $setuphold (posedge USERCLK2, posedge TRNTD[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[111]);
    $setuphold (posedge USERCLK2, posedge TRNTD[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[112]);
    $setuphold (posedge USERCLK2, posedge TRNTD[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[113]);
    $setuphold (posedge USERCLK2, posedge TRNTD[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[114]);
    $setuphold (posedge USERCLK2, posedge TRNTD[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[115]);
    $setuphold (posedge USERCLK2, posedge TRNTD[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[116]);
    $setuphold (posedge USERCLK2, posedge TRNTD[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[117]);
    $setuphold (posedge USERCLK2, posedge TRNTD[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[118]);
    $setuphold (posedge USERCLK2, posedge TRNTD[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[119]);
    $setuphold (posedge USERCLK2, posedge TRNTD[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[11]);
    $setuphold (posedge USERCLK2, posedge TRNTD[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[120]);
    $setuphold (posedge USERCLK2, posedge TRNTD[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[121]);
    $setuphold (posedge USERCLK2, posedge TRNTD[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[122]);
    $setuphold (posedge USERCLK2, posedge TRNTD[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[123]);
    $setuphold (posedge USERCLK2, posedge TRNTD[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[124]);
    $setuphold (posedge USERCLK2, posedge TRNTD[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[125]);
    $setuphold (posedge USERCLK2, posedge TRNTD[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[126]);
    $setuphold (posedge USERCLK2, posedge TRNTD[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[127]);
    $setuphold (posedge USERCLK2, posedge TRNTD[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[12]);
    $setuphold (posedge USERCLK2, posedge TRNTD[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[13]);
    $setuphold (posedge USERCLK2, posedge TRNTD[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[14]);
    $setuphold (posedge USERCLK2, posedge TRNTD[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[15]);
    $setuphold (posedge USERCLK2, posedge TRNTD[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[16]);
    $setuphold (posedge USERCLK2, posedge TRNTD[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[17]);
    $setuphold (posedge USERCLK2, posedge TRNTD[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[18]);
    $setuphold (posedge USERCLK2, posedge TRNTD[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[19]);
    $setuphold (posedge USERCLK2, posedge TRNTD[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[1]);
    $setuphold (posedge USERCLK2, posedge TRNTD[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[20]);
    $setuphold (posedge USERCLK2, posedge TRNTD[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[21]);
    $setuphold (posedge USERCLK2, posedge TRNTD[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[22]);
    $setuphold (posedge USERCLK2, posedge TRNTD[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[23]);
    $setuphold (posedge USERCLK2, posedge TRNTD[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[24]);
    $setuphold (posedge USERCLK2, posedge TRNTD[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[25]);
    $setuphold (posedge USERCLK2, posedge TRNTD[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[26]);
    $setuphold (posedge USERCLK2, posedge TRNTD[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[27]);
    $setuphold (posedge USERCLK2, posedge TRNTD[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[28]);
    $setuphold (posedge USERCLK2, posedge TRNTD[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[29]);
    $setuphold (posedge USERCLK2, posedge TRNTD[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[2]);
    $setuphold (posedge USERCLK2, posedge TRNTD[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[30]);
    $setuphold (posedge USERCLK2, posedge TRNTD[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[31]);
    $setuphold (posedge USERCLK2, posedge TRNTD[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[32]);
    $setuphold (posedge USERCLK2, posedge TRNTD[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[33]);
    $setuphold (posedge USERCLK2, posedge TRNTD[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[34]);
    $setuphold (posedge USERCLK2, posedge TRNTD[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[35]);
    $setuphold (posedge USERCLK2, posedge TRNTD[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[36]);
    $setuphold (posedge USERCLK2, posedge TRNTD[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[37]);
    $setuphold (posedge USERCLK2, posedge TRNTD[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[38]);
    $setuphold (posedge USERCLK2, posedge TRNTD[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[39]);
    $setuphold (posedge USERCLK2, posedge TRNTD[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[3]);
    $setuphold (posedge USERCLK2, posedge TRNTD[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[40]);
    $setuphold (posedge USERCLK2, posedge TRNTD[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[41]);
    $setuphold (posedge USERCLK2, posedge TRNTD[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[42]);
    $setuphold (posedge USERCLK2, posedge TRNTD[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[43]);
    $setuphold (posedge USERCLK2, posedge TRNTD[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[44]);
    $setuphold (posedge USERCLK2, posedge TRNTD[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[45]);
    $setuphold (posedge USERCLK2, posedge TRNTD[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[46]);
    $setuphold (posedge USERCLK2, posedge TRNTD[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[47]);
    $setuphold (posedge USERCLK2, posedge TRNTD[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[48]);
    $setuphold (posedge USERCLK2, posedge TRNTD[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[49]);
    $setuphold (posedge USERCLK2, posedge TRNTD[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[4]);
    $setuphold (posedge USERCLK2, posedge TRNTD[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[50]);
    $setuphold (posedge USERCLK2, posedge TRNTD[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[51]);
    $setuphold (posedge USERCLK2, posedge TRNTD[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[52]);
    $setuphold (posedge USERCLK2, posedge TRNTD[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[53]);
    $setuphold (posedge USERCLK2, posedge TRNTD[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[54]);
    $setuphold (posedge USERCLK2, posedge TRNTD[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[55]);
    $setuphold (posedge USERCLK2, posedge TRNTD[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[56]);
    $setuphold (posedge USERCLK2, posedge TRNTD[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[57]);
    $setuphold (posedge USERCLK2, posedge TRNTD[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[58]);
    $setuphold (posedge USERCLK2, posedge TRNTD[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[59]);
    $setuphold (posedge USERCLK2, posedge TRNTD[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[5]);
    $setuphold (posedge USERCLK2, posedge TRNTD[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[60]);
    $setuphold (posedge USERCLK2, posedge TRNTD[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[61]);
    $setuphold (posedge USERCLK2, posedge TRNTD[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[62]);
    $setuphold (posedge USERCLK2, posedge TRNTD[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[63]);
    $setuphold (posedge USERCLK2, posedge TRNTD[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[64]);
    $setuphold (posedge USERCLK2, posedge TRNTD[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[65]);
    $setuphold (posedge USERCLK2, posedge TRNTD[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[66]);
    $setuphold (posedge USERCLK2, posedge TRNTD[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[67]);
    $setuphold (posedge USERCLK2, posedge TRNTD[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[68]);
    $setuphold (posedge USERCLK2, posedge TRNTD[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[69]);
    $setuphold (posedge USERCLK2, posedge TRNTD[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[6]);
    $setuphold (posedge USERCLK2, posedge TRNTD[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[70]);
    $setuphold (posedge USERCLK2, posedge TRNTD[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[71]);
    $setuphold (posedge USERCLK2, posedge TRNTD[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[72]);
    $setuphold (posedge USERCLK2, posedge TRNTD[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[73]);
    $setuphold (posedge USERCLK2, posedge TRNTD[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[74]);
    $setuphold (posedge USERCLK2, posedge TRNTD[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[75]);
    $setuphold (posedge USERCLK2, posedge TRNTD[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[76]);
    $setuphold (posedge USERCLK2, posedge TRNTD[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[77]);
    $setuphold (posedge USERCLK2, posedge TRNTD[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[78]);
    $setuphold (posedge USERCLK2, posedge TRNTD[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[79]);
    $setuphold (posedge USERCLK2, posedge TRNTD[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[7]);
    $setuphold (posedge USERCLK2, posedge TRNTD[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[80]);
    $setuphold (posedge USERCLK2, posedge TRNTD[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[81]);
    $setuphold (posedge USERCLK2, posedge TRNTD[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[82]);
    $setuphold (posedge USERCLK2, posedge TRNTD[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[83]);
    $setuphold (posedge USERCLK2, posedge TRNTD[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[84]);
    $setuphold (posedge USERCLK2, posedge TRNTD[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[85]);
    $setuphold (posedge USERCLK2, posedge TRNTD[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[86]);
    $setuphold (posedge USERCLK2, posedge TRNTD[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[87]);
    $setuphold (posedge USERCLK2, posedge TRNTD[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[88]);
    $setuphold (posedge USERCLK2, posedge TRNTD[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[89]);
    $setuphold (posedge USERCLK2, posedge TRNTD[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[8]);
    $setuphold (posedge USERCLK2, posedge TRNTD[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[90]);
    $setuphold (posedge USERCLK2, posedge TRNTD[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[91]);
    $setuphold (posedge USERCLK2, posedge TRNTD[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[92]);
    $setuphold (posedge USERCLK2, posedge TRNTD[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[93]);
    $setuphold (posedge USERCLK2, posedge TRNTD[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[94]);
    $setuphold (posedge USERCLK2, posedge TRNTD[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[95]);
    $setuphold (posedge USERCLK2, posedge TRNTD[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[96]);
    $setuphold (posedge USERCLK2, posedge TRNTD[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[97]);
    $setuphold (posedge USERCLK2, posedge TRNTD[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[98]);
    $setuphold (posedge USERCLK2, posedge TRNTD[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[99]);
    $setuphold (posedge USERCLK2, posedge TRNTD[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTD[9]);
    $setuphold (posedge USERCLK2, posedge TRNTECRCGEN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTECRCGEN);
    $setuphold (posedge USERCLK2, posedge TRNTEOF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTEOF);
    $setuphold (posedge USERCLK2, posedge TRNTERRFWD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTERRFWD);
    $setuphold (posedge USERCLK2, posedge TRNTREM[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTREM[0]);
    $setuphold (posedge USERCLK2, posedge TRNTREM[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTREM[1]);
    $setuphold (posedge USERCLK2, posedge TRNTSOF, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSOF);
    $setuphold (posedge USERCLK2, posedge TRNTSRCDSC, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSRCDSC);
    $setuphold (posedge USERCLK2, posedge TRNTSRCRDY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSRCRDY);
    $setuphold (posedge USERCLK2, posedge TRNTSTR, 0:0:0, 0:0:0, notifier,,, delay_USERCLK2, delay_TRNTSTR);
`endif

    ( DRPCLK *> DRPDO[0]) = (0, 0);
    ( DRPCLK *> DRPDO[10]) = (0, 0);
    ( DRPCLK *> DRPDO[11]) = (0, 0);
    ( DRPCLK *> DRPDO[12]) = (0, 0);
    ( DRPCLK *> DRPDO[13]) = (0, 0);
    ( DRPCLK *> DRPDO[14]) = (0, 0);
    ( DRPCLK *> DRPDO[15]) = (0, 0);
    ( DRPCLK *> DRPDO[1]) = (0, 0);
    ( DRPCLK *> DRPDO[2]) = (0, 0);
    ( DRPCLK *> DRPDO[3]) = (0, 0);
    ( DRPCLK *> DRPDO[4]) = (0, 0);
    ( DRPCLK *> DRPDO[5]) = (0, 0);
    ( DRPCLK *> DRPDO[6]) = (0, 0);
    ( DRPCLK *> DRPDO[7]) = (0, 0);
    ( DRPCLK *> DRPDO[8]) = (0, 0);
    ( DRPCLK *> DRPDO[9]) = (0, 0);
    ( DRPCLK *> DRPRDY) = (0, 0);
    ( PIPECLK *> PIPERX0POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX1POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX2POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX3POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX4POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX5POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX6POLARITY) = (0, 0);
    ( PIPECLK *> PIPERX7POLARITY) = (0, 0);
    ( PIPECLK *> PIPETX0CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX0CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX0COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX0DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX0ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX0POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX0POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX1CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX1CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX1COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX1DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX1ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX1POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX1POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX2CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX2CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX2COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX2DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX2ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX2POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX2POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX3CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX3CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX3COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX3DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX3ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX3POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX3POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX4CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX4CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX4COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX4DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX4ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX4POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX4POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX5CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX5CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX5COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX5DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX5ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX5POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX5POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX6CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX6CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX6COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX6DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX6ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX6POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX6POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETX7CHARISK[0]) = (0, 0);
    ( PIPECLK *> PIPETX7CHARISK[1]) = (0, 0);
    ( PIPECLK *> PIPETX7COMPLIANCE) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[0]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[10]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[11]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[12]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[13]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[14]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[15]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[1]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[2]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[3]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[4]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[5]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[6]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[7]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[8]) = (0, 0);
    ( PIPECLK *> PIPETX7DATA[9]) = (0, 0);
    ( PIPECLK *> PIPETX7ELECIDLE) = (0, 0);
    ( PIPECLK *> PIPETX7POWERDOWN[0]) = (0, 0);
    ( PIPECLK *> PIPETX7POWERDOWN[1]) = (0, 0);
    ( PIPECLK *> PIPETXDEEMPH) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[0]) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[1]) = (0, 0);
    ( PIPECLK *> PIPETXMARGIN[2]) = (0, 0);
    ( PIPECLK *> PIPETXRATE) = (0, 0);
    ( PIPECLK *> PIPETXRCVRDET) = (0, 0);
    ( PIPECLK *> PIPETXRESET) = (0, 0);
    ( PIPECLK *> PLDBGVEC[0]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[10]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[11]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[1]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[2]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[3]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[4]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[5]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[6]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[7]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[8]) = (0, 0);
    ( PIPECLK *> PLDBGVEC[9]) = (0, 0);
    ( PIPECLK *> PLDIRECTEDCHANGEDONE) = (0, 0);
    ( PIPECLK *> PLINITIALLINKWIDTH[0]) = (0, 0);
    ( PIPECLK *> PLINITIALLINKWIDTH[1]) = (0, 0);
    ( PIPECLK *> PLINITIALLINKWIDTH[2]) = (0, 0);
    ( PIPECLK *> PLLANEREVERSALMODE[0]) = (0, 0);
    ( PIPECLK *> PLLANEREVERSALMODE[1]) = (0, 0);
    ( PIPECLK *> PLLINKGEN2CAP) = (0, 0);
    ( PIPECLK *> PLLINKPARTNERGEN2SUPPORTED) = (0, 0);
    ( PIPECLK *> PLLINKUPCFGCAP) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[0]) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[1]) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[2]) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[3]) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[4]) = (0, 0);
    ( PIPECLK *> PLLTSSMSTATE[5]) = (0, 0);
    ( PIPECLK *> PLPHYLNKUPN) = (0, 0);
    ( PIPECLK *> PLRECEIVEDHOTRST) = (0, 0);
    ( PIPECLK *> PLRXPMSTATE[0]) = (0, 0);
    ( PIPECLK *> PLRXPMSTATE[1]) = (0, 0);
    ( PIPECLK *> PLSELLNKRATE) = (0, 0);
    ( PIPECLK *> PLSELLNKWIDTH[0]) = (0, 0);
    ( PIPECLK *> PLSELLNKWIDTH[1]) = (0, 0);
    ( PIPECLK *> PLTXPMSTATE[0]) = (0, 0);
    ( PIPECLK *> PLTXPMSTATE[1]) = (0, 0);
    ( PIPECLK *> PLTXPMSTATE[2]) = (0, 0);
    ( USERCLK *> LNKCLKEN) = (0, 0);
    ( USERCLK *> MIMRXRADDR[0]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[10]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[11]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[12]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[1]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[2]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[3]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[4]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[5]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[6]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[7]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[8]) = (0, 0);
    ( USERCLK *> MIMRXRADDR[9]) = (0, 0);
    ( USERCLK *> MIMRXREN) = (0, 0);
    ( USERCLK *> MIMRXWADDR[0]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[10]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[11]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[12]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[1]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[2]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[3]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[4]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[5]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[6]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[7]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[8]) = (0, 0);
    ( USERCLK *> MIMRXWADDR[9]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[0]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[10]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[11]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[12]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[13]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[14]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[15]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[16]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[17]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[18]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[19]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[1]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[20]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[21]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[22]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[23]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[24]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[25]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[26]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[27]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[28]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[29]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[2]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[30]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[31]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[32]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[33]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[34]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[35]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[36]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[37]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[38]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[39]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[3]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[40]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[41]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[42]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[43]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[44]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[45]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[46]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[47]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[48]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[49]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[4]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[50]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[51]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[52]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[53]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[54]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[55]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[56]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[57]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[58]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[59]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[5]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[60]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[61]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[62]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[63]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[64]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[65]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[66]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[67]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[6]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[7]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[8]) = (0, 0);
    ( USERCLK *> MIMRXWDATA[9]) = (0, 0);
    ( USERCLK *> MIMRXWEN) = (0, 0);
    ( USERCLK *> MIMTXRADDR[0]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[10]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[11]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[12]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[1]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[2]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[3]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[4]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[5]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[6]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[7]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[8]) = (0, 0);
    ( USERCLK *> MIMTXRADDR[9]) = (0, 0);
    ( USERCLK *> MIMTXREN) = (0, 0);
    ( USERCLK *> MIMTXWADDR[0]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[10]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[11]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[12]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[1]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[2]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[3]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[4]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[5]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[6]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[7]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[8]) = (0, 0);
    ( USERCLK *> MIMTXWADDR[9]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[0]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[10]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[11]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[12]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[13]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[14]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[15]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[16]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[17]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[18]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[19]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[1]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[20]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[21]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[22]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[23]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[24]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[25]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[26]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[27]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[28]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[29]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[2]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[30]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[31]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[32]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[33]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[34]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[35]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[36]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[37]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[38]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[39]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[3]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[40]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[41]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[42]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[43]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[44]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[45]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[46]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[47]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[48]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[49]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[4]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[50]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[51]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[52]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[53]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[54]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[55]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[56]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[57]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[58]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[59]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[5]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[60]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[61]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[62]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[63]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[64]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[65]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[66]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[67]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[68]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[6]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[7]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[8]) = (0, 0);
    ( USERCLK *> MIMTXWDATA[9]) = (0, 0);
    ( USERCLK *> MIMTXWEN) = (0, 0);
    ( USERCLK2 *> CFGAERECRCCHECKEN) = (0, 0);
    ( USERCLK2 *> CFGAERECRCGENEN) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRCORRERRRECEIVED) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRCORRERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRFATALERRRECEIVED) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRFATALERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRNONFATALERRRECEIVED) = (0, 0);
    ( USERCLK2 *> CFGAERROOTERRNONFATALERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGBRIDGESERREN) = (0, 0);
    ( USERCLK2 *> CFGCOMMANDBUSMASTERENABLE) = (0, 0);
    ( USERCLK2 *> CFGCOMMANDINTERRUPTDISABLE) = (0, 0);
    ( USERCLK2 *> CFGCOMMANDIOENABLE) = (0, 0);
    ( USERCLK2 *> CFGCOMMANDMEMENABLE) = (0, 0);
    ( USERCLK2 *> CFGCOMMANDSERREN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2ARIFORWARDEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2ATOMICEGRESSBLOCK) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2ATOMICREQUESTEREN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2CPLTIMEOUTDIS) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2CPLTIMEOUTVAL[0]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2CPLTIMEOUTVAL[1]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2CPLTIMEOUTVAL[2]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2CPLTIMEOUTVAL[3]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2IDOCPLEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2IDOREQEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2LTREN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROL2TLPPREFIXBLOCK) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLAUXPOWEREN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLCORRERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLENABLERO) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLEXTTAGEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLFATALERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXPAYLOAD[0]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXPAYLOAD[1]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXPAYLOAD[2]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXREADREQ[0]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXREADREQ[1]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLMAXREADREQ[2]) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLNONFATALREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLNOSNOOPEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLPHANTOMEN) = (0, 0);
    ( USERCLK2 *> CFGDEVCONTROLURERRREPORTINGEN) = (0, 0);
    ( USERCLK2 *> CFGDEVSTATUSCORRERRDETECTED) = (0, 0);
    ( USERCLK2 *> CFGDEVSTATUSFATALERRDETECTED) = (0, 0);
    ( USERCLK2 *> CFGDEVSTATUSNONFATALERRDETECTED) = (0, 0);
    ( USERCLK2 *> CFGDEVSTATUSURDETECTED) = (0, 0);
    ( USERCLK2 *> CFGERRAERHEADERLOGSETN) = (0, 0);
    ( USERCLK2 *> CFGERRCPLRDYN) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[0]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[1]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[2]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[3]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[4]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[5]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[6]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTDO[7]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMMENABLE[0]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMMENABLE[1]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMMENABLE[2]) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMSIENABLE) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMSIXENABLE) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTMSIXFM) = (0, 0);
    ( USERCLK2 *> CFGINTERRUPTRDYN) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLASPMCONTROL[0]) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLASPMCONTROL[1]) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLAUTOBANDWIDTHINTEN) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLBANDWIDTHINTEN) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLCLOCKPMEN) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLCOMMONCLOCK) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLEXTENDEDSYNC) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLHWAUTOWIDTHDIS) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLLINKDISABLE) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLRCB) = (0, 0);
    ( USERCLK2 *> CFGLINKCONTROLRETRAINLINK) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSAUTOBANDWIDTHSTATUS) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSBANDWIDTHSTATUS) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSCURRENTSPEED[0]) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSCURRENTSPEED[1]) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSDLLACTIVE) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSLINKTRAINING) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSNEGOTIATEDWIDTH[0]) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSNEGOTIATEDWIDTH[1]) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSNEGOTIATEDWIDTH[2]) = (0, 0);
    ( USERCLK2 *> CFGLINKSTATUSNEGOTIATEDWIDTH[3]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[0]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[10]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[11]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[12]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[13]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[14]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[15]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[16]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[17]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[18]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[19]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[1]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[20]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[21]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[22]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[23]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[24]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[25]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[26]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[27]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[28]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[29]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[2]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[30]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[31]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[3]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[4]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[5]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[6]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[7]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[8]) = (0, 0);
    ( USERCLK2 *> CFGMGMTDO[9]) = (0, 0);
    ( USERCLK2 *> CFGMGMTRDWRDONEN) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[0]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[10]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[11]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[12]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[13]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[14]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[15]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[1]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[2]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[3]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[4]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[5]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[6]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[7]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[8]) = (0, 0);
    ( USERCLK2 *> CFGMSGDATA[9]) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVED) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDASSERTINTA) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDASSERTINTB) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDASSERTINTC) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDASSERTINTD) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDDEASSERTINTA) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDDEASSERTINTB) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDDEASSERTINTC) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDDEASSERTINTD) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDERRCOR) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDERRFATAL) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDERRNONFATAL) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDPMASNAK) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDPMETO) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDPMETOACK) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDPMPME) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDSETSLOTPOWERLIMIT) = (0, 0);
    ( USERCLK2 *> CFGMSGRECEIVEDUNLOCK) = (0, 0);
    ( USERCLK2 *> CFGPCIELINKSTATE[0]) = (0, 0);
    ( USERCLK2 *> CFGPCIELINKSTATE[1]) = (0, 0);
    ( USERCLK2 *> CFGPCIELINKSTATE[2]) = (0, 0);
    ( USERCLK2 *> CFGPMCSRPMEEN) = (0, 0);
    ( USERCLK2 *> CFGPMCSRPMESTATUS) = (0, 0);
    ( USERCLK2 *> CFGPMCSRPOWERSTATE[0]) = (0, 0);
    ( USERCLK2 *> CFGPMCSRPOWERSTATE[1]) = (0, 0);
    ( USERCLK2 *> CFGPMRCVASREQL1N) = (0, 0);
    ( USERCLK2 *> CFGPMRCVENTERL1N) = (0, 0);
    ( USERCLK2 *> CFGPMRCVENTERL23N) = (0, 0);
    ( USERCLK2 *> CFGPMRCVREQACKN) = (0, 0);
    ( USERCLK2 *> CFGROOTCONTROLPMEINTEN) = (0, 0);
    ( USERCLK2 *> CFGROOTCONTROLSYSERRCORRERREN) = (0, 0);
    ( USERCLK2 *> CFGROOTCONTROLSYSERRFATALERREN) = (0, 0);
    ( USERCLK2 *> CFGROOTCONTROLSYSERRNONFATALERREN) = (0, 0);
    ( USERCLK2 *> CFGSLOTCONTROLELECTROMECHILCTLPULSE) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTION) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[0]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[1]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[2]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[3]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[4]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[5]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONADDR[6]) = (0, 0);
    ( USERCLK2 *> CFGTRANSACTIONTYPE) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[0]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[1]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[2]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[3]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[4]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[5]) = (0, 0);
    ( USERCLK2 *> CFGVCTCVCMAP[6]) = (0, 0);
    ( USERCLK2 *> DBGSCLRA) = (0, 0);
    ( USERCLK2 *> DBGSCLRB) = (0, 0);
    ( USERCLK2 *> DBGSCLRC) = (0, 0);
    ( USERCLK2 *> DBGSCLRD) = (0, 0);
    ( USERCLK2 *> DBGSCLRE) = (0, 0);
    ( USERCLK2 *> DBGSCLRF) = (0, 0);
    ( USERCLK2 *> DBGSCLRG) = (0, 0);
    ( USERCLK2 *> DBGSCLRH) = (0, 0);
    ( USERCLK2 *> DBGSCLRI) = (0, 0);
    ( USERCLK2 *> DBGSCLRJ) = (0, 0);
    ( USERCLK2 *> DBGSCLRK) = (0, 0);
    ( USERCLK2 *> DBGVECA[0]) = (0, 0);
    ( USERCLK2 *> DBGVECA[10]) = (0, 0);
    ( USERCLK2 *> DBGVECA[11]) = (0, 0);
    ( USERCLK2 *> DBGVECA[12]) = (0, 0);
    ( USERCLK2 *> DBGVECA[13]) = (0, 0);
    ( USERCLK2 *> DBGVECA[14]) = (0, 0);
    ( USERCLK2 *> DBGVECA[15]) = (0, 0);
    ( USERCLK2 *> DBGVECA[16]) = (0, 0);
    ( USERCLK2 *> DBGVECA[17]) = (0, 0);
    ( USERCLK2 *> DBGVECA[18]) = (0, 0);
    ( USERCLK2 *> DBGVECA[19]) = (0, 0);
    ( USERCLK2 *> DBGVECA[1]) = (0, 0);
    ( USERCLK2 *> DBGVECA[20]) = (0, 0);
    ( USERCLK2 *> DBGVECA[21]) = (0, 0);
    ( USERCLK2 *> DBGVECA[22]) = (0, 0);
    ( USERCLK2 *> DBGVECA[23]) = (0, 0);
    ( USERCLK2 *> DBGVECA[24]) = (0, 0);
    ( USERCLK2 *> DBGVECA[25]) = (0, 0);
    ( USERCLK2 *> DBGVECA[26]) = (0, 0);
    ( USERCLK2 *> DBGVECA[27]) = (0, 0);
    ( USERCLK2 *> DBGVECA[28]) = (0, 0);
    ( USERCLK2 *> DBGVECA[29]) = (0, 0);
    ( USERCLK2 *> DBGVECA[2]) = (0, 0);
    ( USERCLK2 *> DBGVECA[30]) = (0, 0);
    ( USERCLK2 *> DBGVECA[31]) = (0, 0);
    ( USERCLK2 *> DBGVECA[32]) = (0, 0);
    ( USERCLK2 *> DBGVECA[33]) = (0, 0);
    ( USERCLK2 *> DBGVECA[34]) = (0, 0);
    ( USERCLK2 *> DBGVECA[35]) = (0, 0);
    ( USERCLK2 *> DBGVECA[36]) = (0, 0);
    ( USERCLK2 *> DBGVECA[37]) = (0, 0);
    ( USERCLK2 *> DBGVECA[38]) = (0, 0);
    ( USERCLK2 *> DBGVECA[39]) = (0, 0);
    ( USERCLK2 *> DBGVECA[3]) = (0, 0);
    ( USERCLK2 *> DBGVECA[40]) = (0, 0);
    ( USERCLK2 *> DBGVECA[41]) = (0, 0);
    ( USERCLK2 *> DBGVECA[42]) = (0, 0);
    ( USERCLK2 *> DBGVECA[43]) = (0, 0);
    ( USERCLK2 *> DBGVECA[44]) = (0, 0);
    ( USERCLK2 *> DBGVECA[45]) = (0, 0);
    ( USERCLK2 *> DBGVECA[46]) = (0, 0);
    ( USERCLK2 *> DBGVECA[47]) = (0, 0);
    ( USERCLK2 *> DBGVECA[48]) = (0, 0);
    ( USERCLK2 *> DBGVECA[49]) = (0, 0);
    ( USERCLK2 *> DBGVECA[4]) = (0, 0);
    ( USERCLK2 *> DBGVECA[50]) = (0, 0);
    ( USERCLK2 *> DBGVECA[51]) = (0, 0);
    ( USERCLK2 *> DBGVECA[52]) = (0, 0);
    ( USERCLK2 *> DBGVECA[53]) = (0, 0);
    ( USERCLK2 *> DBGVECA[54]) = (0, 0);
    ( USERCLK2 *> DBGVECA[55]) = (0, 0);
    ( USERCLK2 *> DBGVECA[56]) = (0, 0);
    ( USERCLK2 *> DBGVECA[57]) = (0, 0);
    ( USERCLK2 *> DBGVECA[58]) = (0, 0);
    ( USERCLK2 *> DBGVECA[59]) = (0, 0);
    ( USERCLK2 *> DBGVECA[5]) = (0, 0);
    ( USERCLK2 *> DBGVECA[60]) = (0, 0);
    ( USERCLK2 *> DBGVECA[61]) = (0, 0);
    ( USERCLK2 *> DBGVECA[62]) = (0, 0);
    ( USERCLK2 *> DBGVECA[63]) = (0, 0);
    ( USERCLK2 *> DBGVECA[6]) = (0, 0);
    ( USERCLK2 *> DBGVECA[7]) = (0, 0);
    ( USERCLK2 *> DBGVECA[8]) = (0, 0);
    ( USERCLK2 *> DBGVECA[9]) = (0, 0);
    ( USERCLK2 *> DBGVECB[0]) = (0, 0);
    ( USERCLK2 *> DBGVECB[10]) = (0, 0);
    ( USERCLK2 *> DBGVECB[11]) = (0, 0);
    ( USERCLK2 *> DBGVECB[12]) = (0, 0);
    ( USERCLK2 *> DBGVECB[13]) = (0, 0);
    ( USERCLK2 *> DBGVECB[14]) = (0, 0);
    ( USERCLK2 *> DBGVECB[15]) = (0, 0);
    ( USERCLK2 *> DBGVECB[16]) = (0, 0);
    ( USERCLK2 *> DBGVECB[17]) = (0, 0);
    ( USERCLK2 *> DBGVECB[18]) = (0, 0);
    ( USERCLK2 *> DBGVECB[19]) = (0, 0);
    ( USERCLK2 *> DBGVECB[1]) = (0, 0);
    ( USERCLK2 *> DBGVECB[20]) = (0, 0);
    ( USERCLK2 *> DBGVECB[21]) = (0, 0);
    ( USERCLK2 *> DBGVECB[22]) = (0, 0);
    ( USERCLK2 *> DBGVECB[23]) = (0, 0);
    ( USERCLK2 *> DBGVECB[24]) = (0, 0);
    ( USERCLK2 *> DBGVECB[25]) = (0, 0);
    ( USERCLK2 *> DBGVECB[26]) = (0, 0);
    ( USERCLK2 *> DBGVECB[27]) = (0, 0);
    ( USERCLK2 *> DBGVECB[28]) = (0, 0);
    ( USERCLK2 *> DBGVECB[29]) = (0, 0);
    ( USERCLK2 *> DBGVECB[2]) = (0, 0);
    ( USERCLK2 *> DBGVECB[30]) = (0, 0);
    ( USERCLK2 *> DBGVECB[31]) = (0, 0);
    ( USERCLK2 *> DBGVECB[32]) = (0, 0);
    ( USERCLK2 *> DBGVECB[33]) = (0, 0);
    ( USERCLK2 *> DBGVECB[34]) = (0, 0);
    ( USERCLK2 *> DBGVECB[35]) = (0, 0);
    ( USERCLK2 *> DBGVECB[36]) = (0, 0);
    ( USERCLK2 *> DBGVECB[37]) = (0, 0);
    ( USERCLK2 *> DBGVECB[38]) = (0, 0);
    ( USERCLK2 *> DBGVECB[39]) = (0, 0);
    ( USERCLK2 *> DBGVECB[3]) = (0, 0);
    ( USERCLK2 *> DBGVECB[40]) = (0, 0);
    ( USERCLK2 *> DBGVECB[41]) = (0, 0);
    ( USERCLK2 *> DBGVECB[42]) = (0, 0);
    ( USERCLK2 *> DBGVECB[43]) = (0, 0);
    ( USERCLK2 *> DBGVECB[44]) = (0, 0);
    ( USERCLK2 *> DBGVECB[45]) = (0, 0);
    ( USERCLK2 *> DBGVECB[46]) = (0, 0);
    ( USERCLK2 *> DBGVECB[47]) = (0, 0);
    ( USERCLK2 *> DBGVECB[48]) = (0, 0);
    ( USERCLK2 *> DBGVECB[49]) = (0, 0);
    ( USERCLK2 *> DBGVECB[4]) = (0, 0);
    ( USERCLK2 *> DBGVECB[50]) = (0, 0);
    ( USERCLK2 *> DBGVECB[51]) = (0, 0);
    ( USERCLK2 *> DBGVECB[52]) = (0, 0);
    ( USERCLK2 *> DBGVECB[53]) = (0, 0);
    ( USERCLK2 *> DBGVECB[54]) = (0, 0);
    ( USERCLK2 *> DBGVECB[55]) = (0, 0);
    ( USERCLK2 *> DBGVECB[56]) = (0, 0);
    ( USERCLK2 *> DBGVECB[57]) = (0, 0);
    ( USERCLK2 *> DBGVECB[58]) = (0, 0);
    ( USERCLK2 *> DBGVECB[59]) = (0, 0);
    ( USERCLK2 *> DBGVECB[5]) = (0, 0);
    ( USERCLK2 *> DBGVECB[60]) = (0, 0);
    ( USERCLK2 *> DBGVECB[61]) = (0, 0);
    ( USERCLK2 *> DBGVECB[62]) = (0, 0);
    ( USERCLK2 *> DBGVECB[63]) = (0, 0);
    ( USERCLK2 *> DBGVECB[6]) = (0, 0);
    ( USERCLK2 *> DBGVECB[7]) = (0, 0);
    ( USERCLK2 *> DBGVECB[8]) = (0, 0);
    ( USERCLK2 *> DBGVECB[9]) = (0, 0);
    ( USERCLK2 *> DBGVECC[0]) = (0, 0);
    ( USERCLK2 *> DBGVECC[10]) = (0, 0);
    ( USERCLK2 *> DBGVECC[11]) = (0, 0);
    ( USERCLK2 *> DBGVECC[1]) = (0, 0);
    ( USERCLK2 *> DBGVECC[2]) = (0, 0);
    ( USERCLK2 *> DBGVECC[3]) = (0, 0);
    ( USERCLK2 *> DBGVECC[4]) = (0, 0);
    ( USERCLK2 *> DBGVECC[5]) = (0, 0);
    ( USERCLK2 *> DBGVECC[6]) = (0, 0);
    ( USERCLK2 *> DBGVECC[7]) = (0, 0);
    ( USERCLK2 *> DBGVECC[8]) = (0, 0);
    ( USERCLK2 *> DBGVECC[9]) = (0, 0);
    ( USERCLK2 *> LL2BADDLLPERR) = (0, 0);
    ( USERCLK2 *> LL2BADTLPERR) = (0, 0);
    ( USERCLK2 *> LL2LINKSTATUS[0]) = (0, 0);
    ( USERCLK2 *> LL2LINKSTATUS[1]) = (0, 0);
    ( USERCLK2 *> LL2LINKSTATUS[2]) = (0, 0);
    ( USERCLK2 *> LL2LINKSTATUS[3]) = (0, 0);
    ( USERCLK2 *> LL2LINKSTATUS[4]) = (0, 0);
    ( USERCLK2 *> LL2PROTOCOLERR) = (0, 0);
    ( USERCLK2 *> LL2RECEIVERERR) = (0, 0);
    ( USERCLK2 *> LL2REPLAYROERR) = (0, 0);
    ( USERCLK2 *> LL2REPLAYTOERR) = (0, 0);
    ( USERCLK2 *> LL2SUSPENDOK) = (0, 0);
    ( USERCLK2 *> LL2TFCINIT1SEQ) = (0, 0);
    ( USERCLK2 *> LL2TFCINIT2SEQ) = (0, 0);
    ( USERCLK2 *> LL2TXIDLE) = (0, 0);
    ( USERCLK2 *> PL2L0REQ) = (0, 0);
    ( USERCLK2 *> PL2LINKUP) = (0, 0);
    ( USERCLK2 *> PL2RECEIVERERR) = (0, 0);
    ( USERCLK2 *> PL2RECOVERY) = (0, 0);
    ( USERCLK2 *> PL2RXELECIDLE) = (0, 0);
    ( USERCLK2 *> PL2RXPMSTATE[0]) = (0, 0);
    ( USERCLK2 *> PL2RXPMSTATE[1]) = (0, 0);
    ( USERCLK2 *> PL2SUSPENDOK) = (0, 0);
    ( USERCLK2 *> RECEIVEDFUNCLVLRSTN) = (0, 0);
    ( USERCLK2 *> TL2ASPMSUSPENDCREDITCHECKOK) = (0, 0);
    ( USERCLK2 *> TL2ASPMSUSPENDREQ) = (0, 0);
    ( USERCLK2 *> TL2ERRFCPE) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[0]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[10]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[11]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[12]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[13]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[14]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[15]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[16]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[17]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[18]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[19]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[1]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[20]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[21]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[22]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[23]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[24]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[25]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[26]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[27]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[28]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[29]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[2]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[30]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[31]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[32]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[33]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[34]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[35]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[36]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[37]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[38]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[39]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[3]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[40]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[41]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[42]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[43]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[44]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[45]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[46]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[47]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[48]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[49]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[4]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[50]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[51]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[52]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[53]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[54]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[55]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[56]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[57]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[58]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[59]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[5]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[60]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[61]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[62]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[63]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[6]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[7]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[8]) = (0, 0);
    ( USERCLK2 *> TL2ERRHDR[9]) = (0, 0);
    ( USERCLK2 *> TL2ERRMALFORMED) = (0, 0);
    ( USERCLK2 *> TL2ERRRXOVERFLOW) = (0, 0);
    ( USERCLK2 *> TL2PPMSUSPENDOK) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[0]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[10]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[11]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[1]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[2]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[3]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[4]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[5]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[6]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[7]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[8]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLD[9]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[0]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[1]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[2]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[3]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[4]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[5]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[6]) = (0, 0);
    ( USERCLK2 *> TRNFCCPLH[7]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[0]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[10]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[11]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[1]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[2]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[3]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[4]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[5]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[6]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[7]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[8]) = (0, 0);
    ( USERCLK2 *> TRNFCNPD[9]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[0]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[1]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[2]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[3]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[4]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[5]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[6]) = (0, 0);
    ( USERCLK2 *> TRNFCNPH[7]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[0]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[10]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[11]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[1]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[2]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[3]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[4]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[5]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[6]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[7]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[8]) = (0, 0);
    ( USERCLK2 *> TRNFCPD[9]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[0]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[1]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[2]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[3]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[4]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[5]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[6]) = (0, 0);
    ( USERCLK2 *> TRNFCPH[7]) = (0, 0);
    ( USERCLK2 *> TRNLNKUP) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[0]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[1]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[2]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[3]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[4]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[5]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[6]) = (0, 0);
    ( USERCLK2 *> TRNRBARHIT[7]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[0]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[10]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[11]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[12]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[13]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[14]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[15]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[16]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[17]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[18]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[19]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[1]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[20]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[21]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[22]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[23]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[24]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[25]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[26]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[27]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[28]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[29]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[2]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[30]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[31]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[32]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[33]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[34]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[35]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[36]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[37]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[38]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[39]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[3]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[40]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[41]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[42]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[43]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[44]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[45]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[46]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[47]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[48]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[49]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[4]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[50]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[51]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[52]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[53]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[54]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[55]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[56]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[57]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[58]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[59]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[5]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[60]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[61]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[62]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[63]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[6]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[7]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[8]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPDATA[9]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPSRCRDY[0]) = (0, 0);
    ( USERCLK2 *> TRNRDLLPSRCRDY[1]) = (0, 0);
    ( USERCLK2 *> TRNRD[0]) = (0, 0);
    ( USERCLK2 *> TRNRD[100]) = (0, 0);
    ( USERCLK2 *> TRNRD[101]) = (0, 0);
    ( USERCLK2 *> TRNRD[102]) = (0, 0);
    ( USERCLK2 *> TRNRD[103]) = (0, 0);
    ( USERCLK2 *> TRNRD[104]) = (0, 0);
    ( USERCLK2 *> TRNRD[105]) = (0, 0);
    ( USERCLK2 *> TRNRD[106]) = (0, 0);
    ( USERCLK2 *> TRNRD[107]) = (0, 0);
    ( USERCLK2 *> TRNRD[108]) = (0, 0);
    ( USERCLK2 *> TRNRD[109]) = (0, 0);
    ( USERCLK2 *> TRNRD[10]) = (0, 0);
    ( USERCLK2 *> TRNRD[110]) = (0, 0);
    ( USERCLK2 *> TRNRD[111]) = (0, 0);
    ( USERCLK2 *> TRNRD[112]) = (0, 0);
    ( USERCLK2 *> TRNRD[113]) = (0, 0);
    ( USERCLK2 *> TRNRD[114]) = (0, 0);
    ( USERCLK2 *> TRNRD[115]) = (0, 0);
    ( USERCLK2 *> TRNRD[116]) = (0, 0);
    ( USERCLK2 *> TRNRD[117]) = (0, 0);
    ( USERCLK2 *> TRNRD[118]) = (0, 0);
    ( USERCLK2 *> TRNRD[119]) = (0, 0);
    ( USERCLK2 *> TRNRD[11]) = (0, 0);
    ( USERCLK2 *> TRNRD[120]) = (0, 0);
    ( USERCLK2 *> TRNRD[121]) = (0, 0);
    ( USERCLK2 *> TRNRD[122]) = (0, 0);
    ( USERCLK2 *> TRNRD[123]) = (0, 0);
    ( USERCLK2 *> TRNRD[124]) = (0, 0);
    ( USERCLK2 *> TRNRD[125]) = (0, 0);
    ( USERCLK2 *> TRNRD[126]) = (0, 0);
    ( USERCLK2 *> TRNRD[127]) = (0, 0);
    ( USERCLK2 *> TRNRD[12]) = (0, 0);
    ( USERCLK2 *> TRNRD[13]) = (0, 0);
    ( USERCLK2 *> TRNRD[14]) = (0, 0);
    ( USERCLK2 *> TRNRD[15]) = (0, 0);
    ( USERCLK2 *> TRNRD[16]) = (0, 0);
    ( USERCLK2 *> TRNRD[17]) = (0, 0);
    ( USERCLK2 *> TRNRD[18]) = (0, 0);
    ( USERCLK2 *> TRNRD[19]) = (0, 0);
    ( USERCLK2 *> TRNRD[1]) = (0, 0);
    ( USERCLK2 *> TRNRD[20]) = (0, 0);
    ( USERCLK2 *> TRNRD[21]) = (0, 0);
    ( USERCLK2 *> TRNRD[22]) = (0, 0);
    ( USERCLK2 *> TRNRD[23]) = (0, 0);
    ( USERCLK2 *> TRNRD[24]) = (0, 0);
    ( USERCLK2 *> TRNRD[25]) = (0, 0);
    ( USERCLK2 *> TRNRD[26]) = (0, 0);
    ( USERCLK2 *> TRNRD[27]) = (0, 0);
    ( USERCLK2 *> TRNRD[28]) = (0, 0);
    ( USERCLK2 *> TRNRD[29]) = (0, 0);
    ( USERCLK2 *> TRNRD[2]) = (0, 0);
    ( USERCLK2 *> TRNRD[30]) = (0, 0);
    ( USERCLK2 *> TRNRD[31]) = (0, 0);
    ( USERCLK2 *> TRNRD[32]) = (0, 0);
    ( USERCLK2 *> TRNRD[33]) = (0, 0);
    ( USERCLK2 *> TRNRD[34]) = (0, 0);
    ( USERCLK2 *> TRNRD[35]) = (0, 0);
    ( USERCLK2 *> TRNRD[36]) = (0, 0);
    ( USERCLK2 *> TRNRD[37]) = (0, 0);
    ( USERCLK2 *> TRNRD[38]) = (0, 0);
    ( USERCLK2 *> TRNRD[39]) = (0, 0);
    ( USERCLK2 *> TRNRD[3]) = (0, 0);
    ( USERCLK2 *> TRNRD[40]) = (0, 0);
    ( USERCLK2 *> TRNRD[41]) = (0, 0);
    ( USERCLK2 *> TRNRD[42]) = (0, 0);
    ( USERCLK2 *> TRNRD[43]) = (0, 0);
    ( USERCLK2 *> TRNRD[44]) = (0, 0);
    ( USERCLK2 *> TRNRD[45]) = (0, 0);
    ( USERCLK2 *> TRNRD[46]) = (0, 0);
    ( USERCLK2 *> TRNRD[47]) = (0, 0);
    ( USERCLK2 *> TRNRD[48]) = (0, 0);
    ( USERCLK2 *> TRNRD[49]) = (0, 0);
    ( USERCLK2 *> TRNRD[4]) = (0, 0);
    ( USERCLK2 *> TRNRD[50]) = (0, 0);
    ( USERCLK2 *> TRNRD[51]) = (0, 0);
    ( USERCLK2 *> TRNRD[52]) = (0, 0);
    ( USERCLK2 *> TRNRD[53]) = (0, 0);
    ( USERCLK2 *> TRNRD[54]) = (0, 0);
    ( USERCLK2 *> TRNRD[55]) = (0, 0);
    ( USERCLK2 *> TRNRD[56]) = (0, 0);
    ( USERCLK2 *> TRNRD[57]) = (0, 0);
    ( USERCLK2 *> TRNRD[58]) = (0, 0);
    ( USERCLK2 *> TRNRD[59]) = (0, 0);
    ( USERCLK2 *> TRNRD[5]) = (0, 0);
    ( USERCLK2 *> TRNRD[60]) = (0, 0);
    ( USERCLK2 *> TRNRD[61]) = (0, 0);
    ( USERCLK2 *> TRNRD[62]) = (0, 0);
    ( USERCLK2 *> TRNRD[63]) = (0, 0);
    ( USERCLK2 *> TRNRD[64]) = (0, 0);
    ( USERCLK2 *> TRNRD[65]) = (0, 0);
    ( USERCLK2 *> TRNRD[66]) = (0, 0);
    ( USERCLK2 *> TRNRD[67]) = (0, 0);
    ( USERCLK2 *> TRNRD[68]) = (0, 0);
    ( USERCLK2 *> TRNRD[69]) = (0, 0);
    ( USERCLK2 *> TRNRD[6]) = (0, 0);
    ( USERCLK2 *> TRNRD[70]) = (0, 0);
    ( USERCLK2 *> TRNRD[71]) = (0, 0);
    ( USERCLK2 *> TRNRD[72]) = (0, 0);
    ( USERCLK2 *> TRNRD[73]) = (0, 0);
    ( USERCLK2 *> TRNRD[74]) = (0, 0);
    ( USERCLK2 *> TRNRD[75]) = (0, 0);
    ( USERCLK2 *> TRNRD[76]) = (0, 0);
    ( USERCLK2 *> TRNRD[77]) = (0, 0);
    ( USERCLK2 *> TRNRD[78]) = (0, 0);
    ( USERCLK2 *> TRNRD[79]) = (0, 0);
    ( USERCLK2 *> TRNRD[7]) = (0, 0);
    ( USERCLK2 *> TRNRD[80]) = (0, 0);
    ( USERCLK2 *> TRNRD[81]) = (0, 0);
    ( USERCLK2 *> TRNRD[82]) = (0, 0);
    ( USERCLK2 *> TRNRD[83]) = (0, 0);
    ( USERCLK2 *> TRNRD[84]) = (0, 0);
    ( USERCLK2 *> TRNRD[85]) = (0, 0);
    ( USERCLK2 *> TRNRD[86]) = (0, 0);
    ( USERCLK2 *> TRNRD[87]) = (0, 0);
    ( USERCLK2 *> TRNRD[88]) = (0, 0);
    ( USERCLK2 *> TRNRD[89]) = (0, 0);
    ( USERCLK2 *> TRNRD[8]) = (0, 0);
    ( USERCLK2 *> TRNRD[90]) = (0, 0);
    ( USERCLK2 *> TRNRD[91]) = (0, 0);
    ( USERCLK2 *> TRNRD[92]) = (0, 0);
    ( USERCLK2 *> TRNRD[93]) = (0, 0);
    ( USERCLK2 *> TRNRD[94]) = (0, 0);
    ( USERCLK2 *> TRNRD[95]) = (0, 0);
    ( USERCLK2 *> TRNRD[96]) = (0, 0);
    ( USERCLK2 *> TRNRD[97]) = (0, 0);
    ( USERCLK2 *> TRNRD[98]) = (0, 0);
    ( USERCLK2 *> TRNRD[99]) = (0, 0);
    ( USERCLK2 *> TRNRD[9]) = (0, 0);
    ( USERCLK2 *> TRNRECRCERR) = (0, 0);
    ( USERCLK2 *> TRNREOF) = (0, 0);
    ( USERCLK2 *> TRNRERRFWD) = (0, 0);
    ( USERCLK2 *> TRNRREM[0]) = (0, 0);
    ( USERCLK2 *> TRNRREM[1]) = (0, 0);
    ( USERCLK2 *> TRNRSOF) = (0, 0);
    ( USERCLK2 *> TRNRSRCDSC) = (0, 0);
    ( USERCLK2 *> TRNRSRCRDY) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[0]) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[1]) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[2]) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[3]) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[4]) = (0, 0);
    ( USERCLK2 *> TRNTBUFAV[5]) = (0, 0);
    ( USERCLK2 *> TRNTCFGREQ) = (0, 0);
    ( USERCLK2 *> TRNTDLLPDSTRDY) = (0, 0);
    ( USERCLK2 *> TRNTDSTRDY[0]) = (0, 0);
    ( USERCLK2 *> TRNTDSTRDY[1]) = (0, 0);
    ( USERCLK2 *> TRNTDSTRDY[2]) = (0, 0);
    ( USERCLK2 *> TRNTDSTRDY[3]) = (0, 0);
    ( USERCLK2 *> TRNTERRDROP) = (0, 0);
    ( USERCLK2 *> USERRSTN) = (0, 0);

    specparam PATHPULSE$ = 0;
  endspecify
endmodule
