/*
:name: string_atooct
:description: string.atooct()  tests
:tags: 6.16.9
*/
module top();
	string a = "777";
	int b = a.atooct();
endmodule
