/*
:name: class_member_test_41
:description: Test
:should_fail: 0
:tags: 8.3
*/
class constructible;
function new ();
endfunction : new
endclass