/*
:name: class_member_test_51
:description: Test
:tags: 8.3
*/
class myclass;
function void apply_all();
  foreach (foo[i]) begin
    y = apply_this(foo[i]);
  end
endfunction
endclass