// top.v
// my_incl.vh
// If we have not included file before,
// this symbol _my_incl_vh_ is not defined.

// Start of include contents

// Use parentheses to mitigate any undesired operator precedence issues



  
/*
   mode.vh
*/


   

module top(input clk, input [16-1:0] in1, output [(16 << 2)-1:0] q);
 m1 u1(.clk(clk), .in1(in1), .q(q));
 wire a[10:20];

              reg blob_e; 
      /* wire.h */
reg wire_h;

        

 /* 
  comment
  */ 
endmodule // top
