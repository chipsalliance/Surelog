/*
:name: class_member_test_12
:description: Test
:tags: 8.3
*/
class semaphore;
  local chandle p_handle;
endclass