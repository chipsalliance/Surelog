interface adpcm_if;

logic clk;
logic frame;
logic[3:0] data;
logic bozo;
  
  clocking cb @(posedge clk);
    inout frame;
    //input other;
    inout data;
  endclocking
  
  modport mon_mp (clocking cb);

endinterface: adpcm_if

// This file has been modified from the original.
// Attribution and license:
//----------------------------------------------------------
//   Copyright 2010 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------

