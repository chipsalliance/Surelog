/*
:name: preproc_test_6
:description: Test
:should_fail: 0
:tags: 5.6.4
:type: preprocessing
*/
`define INCEPTION(a, b, c) (a*b-c)
