/*
:name: module_definition
:description: module definition test
:tags: 23.2
*/
module top();

endmodule
