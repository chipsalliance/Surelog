// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: var_local
:description: class with local variable
:tags: 8.18
*/
module class_tb ();
	class a_cls;
		local int a_loc = 2;
	endclass
endmodule
