/*
:name: class_member_test_23
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
extern function void subr(mypkg::foo y[M]);
endclass