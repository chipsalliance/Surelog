/*
:name: class_test_25
:description: Test
:tags: 6.15 8.3
*/
class Foo implements Package::Bar; endclass