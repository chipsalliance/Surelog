module top ();
wire signed [15:0] wire_merged;
endmodule
