module top();
   parameter logic [31:0] P1 = 'x;
   parameter logic [31:0] P2 = 'z;
endmodule // top

