// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: 22.12--line-illegal-4
:description: The level parameter shall be 0, 1, or 2
:should_fail_because: The level parameter shall be 0, 1, or 2
:tags: 22.12
:type: preprocessing
*/
`line 1 "somefile"
