// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: union_test_0
:description: Test
:tags: 7.3
*/
typedef union myunion_fwd;

typedef union { logic a; logic b; } myunion_fwd;

module test;
endmodule
