// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: vector_vectored
:description: vectored vector tests
:tags: 6.9.2
*/
module top();
	tri1 vectored [15:0] a;

endmodule
