// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: typedef_test_0
:description: Test
:tags: 6.18
*/
typedef i_am_a_type_really;

typedef int i_am_a_type_really;

// Multiple forward typedefs are allowed.
typedef i_am_a_type_really;
typedef i_am_a_type_really;

module test;
endmodule
