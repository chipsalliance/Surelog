module dff_diffDataTypes();
input int a;    
input byte b;
input shortint c;
input longint d;
input integer e;
input shortint signed f;

endmodule // dff_diffDataTypes
