/*
:name: variable_assignment
:description: Variable assignment tests
:should_fail: 0
:tags: 6.5
*/
module top();
	int v;

	assign v = 12;
endmodule
