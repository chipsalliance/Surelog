/*
:name: class_test_22
:description: Test
:tags: 6.15 8.3
*/
class Foo extends Package::Bar #(.v1(x),.v2(y)); endclass