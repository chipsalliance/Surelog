// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: localparam_int
:description: localparam integer type
:tags: 6.20.4
*/
module top();
	localparam int p = 123;
endmodule
