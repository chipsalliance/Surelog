/*
:name: class_test_35
:description: Test
:tags: 6.15 8.3
*/
class zzxx;
extern function  void set_port(int ap);
endclass
