/*
:name: associative-arrays-string
:description: Test associative arrays support
:should_fail: 0
:tags: 7.8.2 7.8
*/
module top ();

int arr [ string ];

endmodule
