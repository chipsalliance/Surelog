/*
:name: class_test_13
:description: Test
:tags: 6.15 8.3
*/
class Foo #(int W=8, type Int=int) extends Bar #(x,y,z);
endclass