module top();
   AND and1();
endmodule // top
