module top (input logic b, output logic a);
   assign $root.top.a = b;
endmodule
