/*
:name: 22.11--pragma-basic
:description: Test
:should_fail: 0
:tags: 22.11
:type: preprocessing
*/
`pragma pragma_name "pragma_value"
