module DUT (input i, output o);
  wire i;
  wire o;
  assign o = i;
endmodule
