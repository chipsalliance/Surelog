/*
:name: class_test_26
:description: Test
:should_fail: 0
:tags: 6.15 8.3
*/
class Foo implements Bar#(N); endclass