module nonsynth();

   initial
     #1 a = b;
   

endmodule
