/*
:name: non_blocking_assignment
:description: non-blocking assignment test
:should_fail: 0
:tags: 10.4.2
*/
module top();

logic a;

initial begin
	a <= 2;
end

endmodule
