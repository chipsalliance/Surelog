/*
:name: 22.5.1--define_expansion_23
:description: Test
:should_fail_because: redefinition of `define macro is prohibited
:tags: 22.5.1
:type: preprocessing
*/
`define define "illegal"
