
`include "pack_incl.svh"

module top();
   my_logic a;
   logic b;
   
endmodule
