`ifndef TVIP_AXI_UNDEF_INTERNAL_MACROS_SVH
`define TVIP_AXI_UNDEF_INTERNAL_MACROS_SVH

`undef  tvip_axi_4kb_boundary_mask

`endif
