/*
:name: 22.5.2--undef-basic
:description: Test
:should_fail: 0
:tags: 22.5.2
:type: preprocessing
*/
`define FOO "foo"
`undef FOO
