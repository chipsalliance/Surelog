/*
:name: desc_test_2
:description: Test
:type: preprocessing
:tags: 5.6.4
*/
`ifndef DEBUGGER
`endif
