`ifdef __AST_PKG_SV
`else
`define __AST_PKG_SV

package ast_pkg;
endpackage  // of ast_pkg
`endif  // of __AST_PKG_SV
   
