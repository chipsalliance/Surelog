module top;
   localparam string X = {"abcd", "efgh"};
endmodule
