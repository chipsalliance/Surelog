/*
:name: 22.5.1--define_expansion_22
:description: Test
:tags: 22.5.1
:type: preprocessing
*/
`define max(a,b)((a) > (b) ? (a) : (b))
