/*
:name: preproc_test_11
:description: Test
:tags: 5.6.4
:type: preprocessing
*/
`define LONG_MACRO(
    a,
    b
, c
) \
more text c, b, a \
blah blah macro ends here
