/*
:name: class_test_6
:description: Test
:tags: 6.15 8.3
*/
class Foo extends Bar; endclass