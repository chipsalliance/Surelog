/*
:name: preproc_test_0
:description: Test
:should_fail: 0
:tags: 5.6.4
:type: preprocessing
*/
`define TRUTH
