task iprint_ddr_dq (input integer fd);

   $fdisplay(fd, "INFO: Edge Trigger [%t] ...", $realtime);
   $fdisplay(fd, "i_dqs_pad_bscan_c_1 = %b", i_dqs_pad_bscan_c[1]);
   $fdisplay(fd, "i_dqs_pad_bscan_t_1 = %b", i_dqs_pad_bscan_t[1]);
   $fdisplay(fd, "i_dqs_pad_bscan_c_0 = %b", i_dqs_pad_bscan_c[0]);
   $fdisplay(fd, "i_dqs_pad_bscan_t_0 = %b", i_dqs_pad_bscan_t[0]);
   $fdisplay(fd, "i_dqs_pad_bscan_ie = %b", i_dqs_pad_bscan_ie);
   $fdisplay(fd, "i_dqs_pad_bscan_oe = %b", i_dqs_pad_bscan_oe);
   $fdisplay(fd, "i_dqs_pad_bscan_n = %b", i_dqs_pad_bscan_n);
   $fdisplay(fd, "i_dq_pad_bscan_t_8 = %b", i_dq_pad_bscan_t[8]);
   $fdisplay(fd, "i_dq_pad_bscan_t_7 = %b", i_dq_pad_bscan_t[7]);
   $fdisplay(fd, "i_dq_pad_bscan_t_6 = %b", i_dq_pad_bscan_t[6]);
   $fdisplay(fd, "i_dq_pad_bscan_t_5 = %b", i_dq_pad_bscan_t[5]);
   $fdisplay(fd, "i_dq_pad_bscan_t_4 = %b", i_dq_pad_bscan_t[4]);
   $fdisplay(fd, "i_dq_pad_bscan_t_3 = %b", i_dq_pad_bscan_t[3]);
   $fdisplay(fd, "i_dq_pad_bscan_t_2 = %b", i_dq_pad_bscan_t[2]);
   $fdisplay(fd, "i_dq_pad_bscan_t_1 = %b", i_dq_pad_bscan_t[1]);
   $fdisplay(fd, "i_dq_pad_bscan_t_0 = %b", i_dq_pad_bscan_t[0]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_107 = %b", i_dq_pad_tx_cfg[107]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_106 = %b", i_dq_pad_tx_cfg[106]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_105 = %b", i_dq_pad_tx_cfg[105]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_104 = %b", i_dq_pad_tx_cfg[104]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_103 = %b", i_dq_pad_tx_cfg[103]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_102 = %b", i_dq_pad_tx_cfg[102]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_101 = %b", i_dq_pad_tx_cfg[101]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_99 = %b", i_dq_pad_tx_cfg[99]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_98 = %b", i_dq_pad_tx_cfg[98]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_97 = %b", i_dq_pad_tx_cfg[97]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_96 = %b", i_dq_pad_tx_cfg[96]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_95 = %b", i_dq_pad_tx_cfg[95]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_94 = %b", i_dq_pad_tx_cfg[94]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_93 = %b", i_dq_pad_tx_cfg[93]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_92 = %b", i_dq_pad_tx_cfg[92]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_91 = %b", i_dq_pad_tx_cfg[91]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_90 = %b", i_dq_pad_tx_cfg[90]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_89 = %b", i_dq_pad_tx_cfg[89]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_87 = %b", i_dq_pad_tx_cfg[87]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_86 = %b", i_dq_pad_tx_cfg[86]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_85 = %b", i_dq_pad_tx_cfg[85]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_84 = %b", i_dq_pad_tx_cfg[84]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_83 = %b", i_dq_pad_tx_cfg[83]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_82 = %b", i_dq_pad_tx_cfg[82]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_81 = %b", i_dq_pad_tx_cfg[81]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_80 = %b", i_dq_pad_tx_cfg[80]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_79 = %b", i_dq_pad_tx_cfg[79]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_78 = %b", i_dq_pad_tx_cfg[78]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_77 = %b", i_dq_pad_tx_cfg[77]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_75 = %b", i_dq_pad_tx_cfg[75]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_74 = %b", i_dq_pad_tx_cfg[74]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_73 = %b", i_dq_pad_tx_cfg[73]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_72 = %b", i_dq_pad_tx_cfg[72]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_71 = %b", i_dq_pad_tx_cfg[71]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_70 = %b", i_dq_pad_tx_cfg[70]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_69 = %b", i_dq_pad_tx_cfg[69]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_68 = %b", i_dq_pad_tx_cfg[68]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_67 = %b", i_dq_pad_tx_cfg[67]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_66 = %b", i_dq_pad_tx_cfg[66]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_65 = %b", i_dq_pad_tx_cfg[65]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_63 = %b", i_dq_pad_tx_cfg[63]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_62 = %b", i_dq_pad_tx_cfg[62]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_61 = %b", i_dq_pad_tx_cfg[61]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_60 = %b", i_dq_pad_tx_cfg[60]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_59 = %b", i_dq_pad_tx_cfg[59]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_58 = %b", i_dq_pad_tx_cfg[58]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_57 = %b", i_dq_pad_tx_cfg[57]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_56 = %b", i_dq_pad_tx_cfg[56]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_55 = %b", i_dq_pad_tx_cfg[55]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_54 = %b", i_dq_pad_tx_cfg[54]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_53 = %b", i_dq_pad_tx_cfg[53]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_51 = %b", i_dq_pad_tx_cfg[51]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_50 = %b", i_dq_pad_tx_cfg[50]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_49 = %b", i_dq_pad_tx_cfg[49]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_48 = %b", i_dq_pad_tx_cfg[48]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_47 = %b", i_dq_pad_tx_cfg[47]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_46 = %b", i_dq_pad_tx_cfg[46]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_45 = %b", i_dq_pad_tx_cfg[45]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_44 = %b", i_dq_pad_tx_cfg[44]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_43 = %b", i_dq_pad_tx_cfg[43]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_42 = %b", i_dq_pad_tx_cfg[42]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_41 = %b", i_dq_pad_tx_cfg[41]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_39 = %b", i_dq_pad_tx_cfg[39]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_38 = %b", i_dq_pad_tx_cfg[38]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_37 = %b", i_dq_pad_tx_cfg[37]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_36 = %b", i_dq_pad_tx_cfg[36]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_35 = %b", i_dq_pad_tx_cfg[35]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_34 = %b", i_dq_pad_tx_cfg[34]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_33 = %b", i_dq_pad_tx_cfg[33]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_32 = %b", i_dq_pad_tx_cfg[32]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_31 = %b", i_dq_pad_tx_cfg[31]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_30 = %b", i_dq_pad_tx_cfg[30]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_29 = %b", i_dq_pad_tx_cfg[29]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_27 = %b", i_dq_pad_tx_cfg[27]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_26 = %b", i_dq_pad_tx_cfg[26]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_25 = %b", i_dq_pad_tx_cfg[25]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_24 = %b", i_dq_pad_tx_cfg[24]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_23 = %b", i_dq_pad_tx_cfg[23]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_22 = %b", i_dq_pad_tx_cfg[22]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_21 = %b", i_dq_pad_tx_cfg[21]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_20 = %b", i_dq_pad_tx_cfg[20]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_19 = %b", i_dq_pad_tx_cfg[19]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_18 = %b", i_dq_pad_tx_cfg[18]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_17 = %b", i_dq_pad_tx_cfg[17]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_15 = %b", i_dq_pad_tx_cfg[15]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_14 = %b", i_dq_pad_tx_cfg[14]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_13 = %b", i_dq_pad_tx_cfg[13]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_12 = %b", i_dq_pad_tx_cfg[12]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_11 = %b", i_dq_pad_tx_cfg[11]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_10 = %b", i_dq_pad_tx_cfg[10]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_9 = %b", i_dq_pad_tx_cfg[9]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_8 = %b", i_dq_pad_tx_cfg[8]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_7 = %b", i_dq_pad_tx_cfg[7]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_6 = %b", i_dq_pad_tx_cfg[6]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_5 = %b", i_dq_pad_tx_cfg[5]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_3 = %b", i_dq_pad_tx_cfg[3]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_2 = %b", i_dq_pad_tx_cfg[2]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_1 = %b", i_dq_pad_tx_cfg[1]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_0 = %b", i_dq_pad_tx_cfg[0]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_279 = %b", i_dq_sa_dly_cfg[279]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_278 = %b", i_dq_sa_dly_cfg[278]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_277 = %b", i_dq_sa_dly_cfg[277]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_276 = %b", i_dq_sa_dly_cfg[276]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_275 = %b", i_dq_sa_dly_cfg[275]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_274 = %b", i_dq_sa_dly_cfg[274]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_273 = %b", i_dq_sa_dly_cfg[273]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_272 = %b", i_dq_sa_dly_cfg[272]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_263 = %b", i_dq_sa_dly_cfg[263]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_262 = %b", i_dq_sa_dly_cfg[262]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_261 = %b", i_dq_sa_dly_cfg[261]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_260 = %b", i_dq_sa_dly_cfg[260]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_259 = %b", i_dq_sa_dly_cfg[259]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_258 = %b", i_dq_sa_dly_cfg[258]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_257 = %b", i_dq_sa_dly_cfg[257]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_256 = %b", i_dq_sa_dly_cfg[256]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_247 = %b", i_dq_sa_dly_cfg[247]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_246 = %b", i_dq_sa_dly_cfg[246]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_245 = %b", i_dq_sa_dly_cfg[245]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_244 = %b", i_dq_sa_dly_cfg[244]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_243 = %b", i_dq_sa_dly_cfg[243]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_242 = %b", i_dq_sa_dly_cfg[242]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_241 = %b", i_dq_sa_dly_cfg[241]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_240 = %b", i_dq_sa_dly_cfg[240]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_231 = %b", i_dq_sa_dly_cfg[231]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_230 = %b", i_dq_sa_dly_cfg[230]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_229 = %b", i_dq_sa_dly_cfg[229]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_228 = %b", i_dq_sa_dly_cfg[228]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_227 = %b", i_dq_sa_dly_cfg[227]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_226 = %b", i_dq_sa_dly_cfg[226]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_225 = %b", i_dq_sa_dly_cfg[225]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_224 = %b", i_dq_sa_dly_cfg[224]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_215 = %b", i_dq_sa_dly_cfg[215]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_214 = %b", i_dq_sa_dly_cfg[214]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_213 = %b", i_dq_sa_dly_cfg[213]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_212 = %b", i_dq_sa_dly_cfg[212]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_211 = %b", i_dq_sa_dly_cfg[211]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_210 = %b", i_dq_sa_dly_cfg[210]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_209 = %b", i_dq_sa_dly_cfg[209]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_208 = %b", i_dq_sa_dly_cfg[208]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_199 = %b", i_dq_sa_dly_cfg[199]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_198 = %b", i_dq_sa_dly_cfg[198]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_197 = %b", i_dq_sa_dly_cfg[197]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_196 = %b", i_dq_sa_dly_cfg[196]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_195 = %b", i_dq_sa_dly_cfg[195]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_194 = %b", i_dq_sa_dly_cfg[194]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_193 = %b", i_dq_sa_dly_cfg[193]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_192 = %b", i_dq_sa_dly_cfg[192]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_183 = %b", i_dq_sa_dly_cfg[183]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_182 = %b", i_dq_sa_dly_cfg[182]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_181 = %b", i_dq_sa_dly_cfg[181]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_180 = %b", i_dq_sa_dly_cfg[180]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_179 = %b", i_dq_sa_dly_cfg[179]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_178 = %b", i_dq_sa_dly_cfg[178]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_177 = %b", i_dq_sa_dly_cfg[177]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_176 = %b", i_dq_sa_dly_cfg[176]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_167 = %b", i_dq_sa_dly_cfg[167]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_166 = %b", i_dq_sa_dly_cfg[166]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_165 = %b", i_dq_sa_dly_cfg[165]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_164 = %b", i_dq_sa_dly_cfg[164]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_163 = %b", i_dq_sa_dly_cfg[163]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_162 = %b", i_dq_sa_dly_cfg[162]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_161 = %b", i_dq_sa_dly_cfg[161]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_160 = %b", i_dq_sa_dly_cfg[160]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_151 = %b", i_dq_sa_dly_cfg[151]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_150 = %b", i_dq_sa_dly_cfg[150]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_149 = %b", i_dq_sa_dly_cfg[149]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_148 = %b", i_dq_sa_dly_cfg[148]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_147 = %b", i_dq_sa_dly_cfg[147]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_146 = %b", i_dq_sa_dly_cfg[146]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_145 = %b", i_dq_sa_dly_cfg[145]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_144 = %b", i_dq_sa_dly_cfg[144]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_135 = %b", i_dq_sa_dly_cfg[135]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_134 = %b", i_dq_sa_dly_cfg[134]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_133 = %b", i_dq_sa_dly_cfg[133]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_132 = %b", i_dq_sa_dly_cfg[132]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_131 = %b", i_dq_sa_dly_cfg[131]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_130 = %b", i_dq_sa_dly_cfg[130]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_129 = %b", i_dq_sa_dly_cfg[129]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_128 = %b", i_dq_sa_dly_cfg[128]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_119 = %b", i_dq_sa_dly_cfg[119]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_118 = %b", i_dq_sa_dly_cfg[118]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_117 = %b", i_dq_sa_dly_cfg[117]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_116 = %b", i_dq_sa_dly_cfg[116]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_115 = %b", i_dq_sa_dly_cfg[115]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_114 = %b", i_dq_sa_dly_cfg[114]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_113 = %b", i_dq_sa_dly_cfg[113]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_112 = %b", i_dq_sa_dly_cfg[112]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_103 = %b", i_dq_sa_dly_cfg[103]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_102 = %b", i_dq_sa_dly_cfg[102]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_101 = %b", i_dq_sa_dly_cfg[101]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_100 = %b", i_dq_sa_dly_cfg[100]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_99 = %b", i_dq_sa_dly_cfg[99]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_98 = %b", i_dq_sa_dly_cfg[98]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_97 = %b", i_dq_sa_dly_cfg[97]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_96 = %b", i_dq_sa_dly_cfg[96]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_87 = %b", i_dq_sa_dly_cfg[87]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_86 = %b", i_dq_sa_dly_cfg[86]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_85 = %b", i_dq_sa_dly_cfg[85]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_84 = %b", i_dq_sa_dly_cfg[84]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_83 = %b", i_dq_sa_dly_cfg[83]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_82 = %b", i_dq_sa_dly_cfg[82]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_81 = %b", i_dq_sa_dly_cfg[81]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_80 = %b", i_dq_sa_dly_cfg[80]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_71 = %b", i_dq_sa_dly_cfg[71]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_70 = %b", i_dq_sa_dly_cfg[70]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_69 = %b", i_dq_sa_dly_cfg[69]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_68 = %b", i_dq_sa_dly_cfg[68]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_67 = %b", i_dq_sa_dly_cfg[67]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_66 = %b", i_dq_sa_dly_cfg[66]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_65 = %b", i_dq_sa_dly_cfg[65]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_64 = %b", i_dq_sa_dly_cfg[64]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_55 = %b", i_dq_sa_dly_cfg[55]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_54 = %b", i_dq_sa_dly_cfg[54]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_53 = %b", i_dq_sa_dly_cfg[53]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_52 = %b", i_dq_sa_dly_cfg[52]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_51 = %b", i_dq_sa_dly_cfg[51]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_50 = %b", i_dq_sa_dly_cfg[50]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_49 = %b", i_dq_sa_dly_cfg[49]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_48 = %b", i_dq_sa_dly_cfg[48]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_39 = %b", i_dq_sa_dly_cfg[39]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_38 = %b", i_dq_sa_dly_cfg[38]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_37 = %b", i_dq_sa_dly_cfg[37]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_36 = %b", i_dq_sa_dly_cfg[36]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_35 = %b", i_dq_sa_dly_cfg[35]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_34 = %b", i_dq_sa_dly_cfg[34]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_33 = %b", i_dq_sa_dly_cfg[33]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_32 = %b", i_dq_sa_dly_cfg[32]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_23 = %b", i_dq_sa_dly_cfg[23]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_22 = %b", i_dq_sa_dly_cfg[22]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_21 = %b", i_dq_sa_dly_cfg[21]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_20 = %b", i_dq_sa_dly_cfg[20]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_19 = %b", i_dq_sa_dly_cfg[19]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_18 = %b", i_dq_sa_dly_cfg[18]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_17 = %b", i_dq_sa_dly_cfg[17]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_16 = %b", i_dq_sa_dly_cfg[16]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_7 = %b", i_dq_sa_dly_cfg[7]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_6 = %b", i_dq_sa_dly_cfg[6]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_5 = %b", i_dq_sa_dly_cfg[5]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_4 = %b", i_dq_sa_dly_cfg[4]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_3 = %b", i_dq_sa_dly_cfg[3]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_2 = %b", i_dq_sa_dly_cfg[2]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_1 = %b", i_dq_sa_dly_cfg[1]);
   $fdisplay(fd, "i_dq_sa_dly_cfg_0 = %b", i_dq_sa_dly_cfg[0]);
   $fdisplay(fd, "i_dq_sa_cfg_178 = %b", i_dq_sa_cfg[178]);
   $fdisplay(fd, "i_dq_sa_cfg_176 = %b", i_dq_sa_cfg[176]);
   $fdisplay(fd, "i_dq_sa_cfg_171 = %b", i_dq_sa_cfg[171]);
   $fdisplay(fd, "i_dq_sa_cfg_170 = %b", i_dq_sa_cfg[170]);
   $fdisplay(fd, "i_dq_sa_cfg_169 = %b", i_dq_sa_cfg[169]);
   $fdisplay(fd, "i_dq_sa_cfg_168 = %b", i_dq_sa_cfg[168]);
   $fdisplay(fd, "i_dq_sa_cfg_163 = %b", i_dq_sa_cfg[163]);
   $fdisplay(fd, "i_dq_sa_cfg_162 = %b", i_dq_sa_cfg[162]);
   $fdisplay(fd, "i_dq_sa_cfg_161 = %b", i_dq_sa_cfg[161]);
   $fdisplay(fd, "i_dq_sa_cfg_160 = %b", i_dq_sa_cfg[160]);
   $fdisplay(fd, "i_dq_sa_cfg_158 = %b", i_dq_sa_cfg[158]);
   $fdisplay(fd, "i_dq_sa_cfg_156 = %b", i_dq_sa_cfg[156]);
   $fdisplay(fd, "i_dq_sa_cfg_151 = %b", i_dq_sa_cfg[151]);
   $fdisplay(fd, "i_dq_sa_cfg_150 = %b", i_dq_sa_cfg[150]);
   $fdisplay(fd, "i_dq_sa_cfg_149 = %b", i_dq_sa_cfg[149]);
   $fdisplay(fd, "i_dq_sa_cfg_148 = %b", i_dq_sa_cfg[148]);
   $fdisplay(fd, "i_dq_sa_cfg_143 = %b", i_dq_sa_cfg[143]);
   $fdisplay(fd, "i_dq_sa_cfg_142 = %b", i_dq_sa_cfg[142]);
   $fdisplay(fd, "i_dq_sa_cfg_141 = %b", i_dq_sa_cfg[141]);
   $fdisplay(fd, "i_dq_sa_cfg_140 = %b", i_dq_sa_cfg[140]);
   $fdisplay(fd, "i_dq_sa_cfg_138 = %b", i_dq_sa_cfg[138]);
   $fdisplay(fd, "i_dq_sa_cfg_136 = %b", i_dq_sa_cfg[136]);
   $fdisplay(fd, "i_dq_sa_cfg_131 = %b", i_dq_sa_cfg[131]);
   $fdisplay(fd, "i_dq_sa_cfg_130 = %b", i_dq_sa_cfg[130]);
   $fdisplay(fd, "i_dq_sa_cfg_129 = %b", i_dq_sa_cfg[129]);
   $fdisplay(fd, "i_dq_sa_cfg_128 = %b", i_dq_sa_cfg[128]);
   $fdisplay(fd, "i_dq_sa_cfg_123 = %b", i_dq_sa_cfg[123]);
   $fdisplay(fd, "i_dq_sa_cfg_122 = %b", i_dq_sa_cfg[122]);
   $fdisplay(fd, "i_dq_sa_cfg_121 = %b", i_dq_sa_cfg[121]);
   $fdisplay(fd, "i_dq_sa_cfg_120 = %b", i_dq_sa_cfg[120]);
   $fdisplay(fd, "i_dq_sa_cfg_118 = %b", i_dq_sa_cfg[118]);
   $fdisplay(fd, "i_dq_sa_cfg_116 = %b", i_dq_sa_cfg[116]);
   $fdisplay(fd, "i_dq_sa_cfg_111 = %b", i_dq_sa_cfg[111]);
   $fdisplay(fd, "i_dq_sa_cfg_110 = %b", i_dq_sa_cfg[110]);
   $fdisplay(fd, "i_dq_sa_cfg_109 = %b", i_dq_sa_cfg[109]);
   $fdisplay(fd, "i_dq_sa_cfg_108 = %b", i_dq_sa_cfg[108]);
   $fdisplay(fd, "i_dq_sa_cfg_103 = %b", i_dq_sa_cfg[103]);
   $fdisplay(fd, "i_dq_sa_cfg_102 = %b", i_dq_sa_cfg[102]);
   $fdisplay(fd, "i_dq_sa_cfg_101 = %b", i_dq_sa_cfg[101]);
   $fdisplay(fd, "i_dq_sa_cfg_100 = %b", i_dq_sa_cfg[100]);
   $fdisplay(fd, "i_dq_sa_cfg_98 = %b", i_dq_sa_cfg[98]);
   $fdisplay(fd, "i_dq_sa_cfg_96 = %b", i_dq_sa_cfg[96]);
   $fdisplay(fd, "i_dq_sa_cfg_91 = %b", i_dq_sa_cfg[91]);
   $fdisplay(fd, "i_dq_sa_cfg_90 = %b", i_dq_sa_cfg[90]);
   $fdisplay(fd, "i_dq_sa_cfg_89 = %b", i_dq_sa_cfg[89]);
   $fdisplay(fd, "i_dq_sa_cfg_88 = %b", i_dq_sa_cfg[88]);
   $fdisplay(fd, "i_dq_sa_cfg_83 = %b", i_dq_sa_cfg[83]);
   $fdisplay(fd, "i_dq_sa_cfg_82 = %b", i_dq_sa_cfg[82]);
   $fdisplay(fd, "i_dq_sa_cfg_81 = %b", i_dq_sa_cfg[81]);
   $fdisplay(fd, "i_dq_sa_cfg_80 = %b", i_dq_sa_cfg[80]);
   $fdisplay(fd, "i_dq_sa_cfg_78 = %b", i_dq_sa_cfg[78]);
   $fdisplay(fd, "i_dq_sa_cfg_76 = %b", i_dq_sa_cfg[76]);
   $fdisplay(fd, "i_dq_sa_cfg_71 = %b", i_dq_sa_cfg[71]);
   $fdisplay(fd, "i_dq_sa_cfg_70 = %b", i_dq_sa_cfg[70]);
   $fdisplay(fd, "i_dq_sa_cfg_69 = %b", i_dq_sa_cfg[69]);
   $fdisplay(fd, "i_dq_sa_cfg_68 = %b", i_dq_sa_cfg[68]);
   $fdisplay(fd, "i_dq_sa_cfg_63 = %b", i_dq_sa_cfg[63]);
   $fdisplay(fd, "i_dq_sa_cfg_62 = %b", i_dq_sa_cfg[62]);
   $fdisplay(fd, "i_dq_sa_cfg_61 = %b", i_dq_sa_cfg[61]);
   $fdisplay(fd, "i_dq_sa_cfg_60 = %b", i_dq_sa_cfg[60]);
   $fdisplay(fd, "i_dq_sa_cfg_58 = %b", i_dq_sa_cfg[58]);
   $fdisplay(fd, "i_dq_sa_cfg_56 = %b", i_dq_sa_cfg[56]);
   $fdisplay(fd, "i_dq_sa_cfg_51 = %b", i_dq_sa_cfg[51]);
   $fdisplay(fd, "i_dq_sa_cfg_50 = %b", i_dq_sa_cfg[50]);
   $fdisplay(fd, "i_dq_sa_cfg_49 = %b", i_dq_sa_cfg[49]);
   $fdisplay(fd, "i_dq_sa_cfg_48 = %b", i_dq_sa_cfg[48]);
   $fdisplay(fd, "i_dq_sa_cfg_43 = %b", i_dq_sa_cfg[43]);
   $fdisplay(fd, "i_dq_sa_cfg_42 = %b", i_dq_sa_cfg[42]);
   $fdisplay(fd, "i_dq_sa_cfg_41 = %b", i_dq_sa_cfg[41]);
   $fdisplay(fd, "i_dq_sa_cfg_40 = %b", i_dq_sa_cfg[40]);
   $fdisplay(fd, "i_dq_sa_cfg_38 = %b", i_dq_sa_cfg[38]);
   $fdisplay(fd, "i_dq_sa_cfg_36 = %b", i_dq_sa_cfg[36]);
   $fdisplay(fd, "i_dq_sa_cfg_31 = %b", i_dq_sa_cfg[31]);
   $fdisplay(fd, "i_dq_sa_cfg_30 = %b", i_dq_sa_cfg[30]);
   $fdisplay(fd, "i_dq_sa_cfg_29 = %b", i_dq_sa_cfg[29]);
   $fdisplay(fd, "i_dq_sa_cfg_28 = %b", i_dq_sa_cfg[28]);
   $fdisplay(fd, "i_dq_sa_cfg_23 = %b", i_dq_sa_cfg[23]);
   $fdisplay(fd, "i_dq_sa_cfg_22 = %b", i_dq_sa_cfg[22]);
   $fdisplay(fd, "i_dq_sa_cfg_21 = %b", i_dq_sa_cfg[21]);
   $fdisplay(fd, "i_dq_sa_cfg_20 = %b", i_dq_sa_cfg[20]);
   $fdisplay(fd, "i_dq_sa_cfg_18 = %b", i_dq_sa_cfg[18]);
   $fdisplay(fd, "i_dq_sa_cfg_16 = %b", i_dq_sa_cfg[16]);
   $fdisplay(fd, "i_dq_sa_cfg_11 = %b", i_dq_sa_cfg[11]);
   $fdisplay(fd, "i_dq_sa_cfg_10 = %b", i_dq_sa_cfg[10]);
   $fdisplay(fd, "i_dq_sa_cfg_9 = %b", i_dq_sa_cfg[9]);
   $fdisplay(fd, "i_dq_sa_cfg_8 = %b", i_dq_sa_cfg[8]);
   $fdisplay(fd, "i_dq_sa_cfg_3 = %b", i_dq_sa_cfg[3]);
   $fdisplay(fd, "i_dq_sa_cfg_2 = %b", i_dq_sa_cfg[2]);
   $fdisplay(fd, "i_dq_sa_cfg_1 = %b", i_dq_sa_cfg[1]);
   $fdisplay(fd, "i_dq_sa_cfg_0 = %b", i_dq_sa_cfg[0]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_13 = %b", i_dqs_pad_tx_cmn_cfg[13]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_12 = %b", i_dqs_pad_tx_cmn_cfg[12]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_11 = %b", i_dqs_pad_tx_cmn_cfg[11]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_10 = %b", i_dqs_pad_tx_cmn_cfg[10]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_9 = %b", i_dqs_pad_tx_cmn_cfg[9]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_8 = %b", i_dqs_pad_tx_cmn_cfg[8]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_7 = %b", i_dqs_pad_tx_cmn_cfg[7]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_6 = %b", i_dqs_pad_tx_cmn_cfg[6]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_5 = %b", i_dqs_pad_tx_cmn_cfg[5]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_4 = %b", i_dqs_pad_tx_cmn_cfg[4]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_3 = %b", i_dqs_pad_tx_cmn_cfg[3]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_2 = %b", i_dqs_pad_tx_cmn_cfg[2]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_1 = %b", i_dqs_pad_tx_cmn_cfg[1]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_0 = %b", i_dqs_pad_tx_cmn_cfg[0]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_23 = %b", i_dqs_pad_tx_cfg[23]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_22 = %b", i_dqs_pad_tx_cfg[22]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_21 = %b", i_dqs_pad_tx_cfg[21]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_20 = %b", i_dqs_pad_tx_cfg[20]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_19 = %b", i_dqs_pad_tx_cfg[19]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_18 = %b", i_dqs_pad_tx_cfg[18]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_17 = %b", i_dqs_pad_tx_cfg[17]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_16 = %b", i_dqs_pad_tx_cfg[16]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_15 = %b", i_dqs_pad_tx_cfg[15]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_14 = %b", i_dqs_pad_tx_cfg[14]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_13 = %b", i_dqs_pad_tx_cfg[13]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_12 = %b", i_dqs_pad_tx_cfg[12]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_11 = %b", i_dqs_pad_tx_cfg[11]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_10 = %b", i_dqs_pad_tx_cfg[10]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_9 = %b", i_dqs_pad_tx_cfg[9]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_8 = %b", i_dqs_pad_tx_cfg[8]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_7 = %b", i_dqs_pad_tx_cfg[7]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_6 = %b", i_dqs_pad_tx_cfg[6]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_5 = %b", i_dqs_pad_tx_cfg[5]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_4 = %b", i_dqs_pad_tx_cfg[4]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_3 = %b", i_dqs_pad_tx_cfg[3]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_2 = %b", i_dqs_pad_tx_cfg[2]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_1 = %b", i_dqs_pad_tx_cfg[1]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_0 = %b", i_dqs_pad_tx_cfg[0]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_25 = %b", i_dqs_pad_rx_cmn_cfg[25]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_24 = %b", i_dqs_pad_rx_cmn_cfg[24]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_23 = %b", i_dqs_pad_rx_cmn_cfg[23]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_22 = %b", i_dqs_pad_rx_cmn_cfg[22]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_21 = %b", i_dqs_pad_rx_cmn_cfg[21]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_20 = %b", i_dqs_pad_rx_cmn_cfg[20]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_19 = %b", i_dqs_pad_rx_cmn_cfg[19]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_18 = %b", i_dqs_pad_rx_cmn_cfg[18]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_17 = %b", i_dqs_pad_rx_cmn_cfg[17]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_16 = %b", i_dqs_pad_rx_cmn_cfg[16]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_15 = %b", i_dqs_pad_rx_cmn_cfg[15]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_14 = %b", i_dqs_pad_rx_cmn_cfg[14]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_13 = %b", i_dqs_pad_rx_cmn_cfg[13]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_12 = %b", i_dqs_pad_rx_cmn_cfg[12]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_11 = %b", i_dqs_pad_rx_cmn_cfg[11]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_10 = %b", i_dqs_pad_rx_cmn_cfg[10]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_9 = %b", i_dqs_pad_rx_cmn_cfg[9]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_8 = %b", i_dqs_pad_rx_cmn_cfg[8]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_7 = %b", i_dqs_pad_rx_cmn_cfg[7]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_6 = %b", i_dqs_pad_rx_cmn_cfg[6]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_5 = %b", i_dqs_pad_rx_cmn_cfg[5]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_4 = %b", i_dqs_pad_rx_cmn_cfg[4]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_3 = %b", i_dqs_pad_rx_cmn_cfg[3]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_2 = %b", i_dqs_pad_rx_cmn_cfg[2]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_1 = %b", i_dqs_pad_rx_cmn_cfg[1]);
   $fdisplay(fd, "i_dqs_pad_rx_cmn_cfg_0 = %b", i_dqs_pad_rx_cmn_cfg[0]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_31 = %b", i_dqs_pad_rx_cfg[31]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_30 = %b", i_dqs_pad_rx_cfg[30]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_29 = %b", i_dqs_pad_rx_cfg[29]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_28 = %b", i_dqs_pad_rx_cfg[28]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_27 = %b", i_dqs_pad_rx_cfg[27]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_26 = %b", i_dqs_pad_rx_cfg[26]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_25 = %b", i_dqs_pad_rx_cfg[25]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_24 = %b", i_dqs_pad_rx_cfg[24]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_23 = %b", i_dqs_pad_rx_cfg[23]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_22 = %b", i_dqs_pad_rx_cfg[22]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_21 = %b", i_dqs_pad_rx_cfg[21]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_20 = %b", i_dqs_pad_rx_cfg[20]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_19 = %b", i_dqs_pad_rx_cfg[19]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_18 = %b", i_dqs_pad_rx_cfg[18]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_17 = %b", i_dqs_pad_rx_cfg[17]);
   $fdisplay(fd, "i_dqs_pad_rx_cfg_16 = %b", i_dqs_pad_rx_cfg[16]);
   $fdisplay(fd, "i_dqs_sa_cmn_cfg_4 = %b", i_dqs_sa_cmn_cfg[4]);
   $fdisplay(fd, "i_dqs_sa_cmn_cfg_1 = %b", i_dqs_sa_cmn_cfg[1]);
   $fdisplay(fd, "i_dqs_sa_cmn_cfg_0 = %b", i_dqs_sa_cmn_cfg[0]);
   $fdisplay(fd, "i_dqs_hiz_n = %b", i_dqs_hiz_n);
   //`display( "i_dqs_freeze_n = %b", i_dqs_freeze_n); // 20201230 release
   $fdisplay(fd, "i_dq_cmn_freeze_n = %b", i_dq_cmn_freeze_n);
   //`display( "i_dq_freeze_n_hv = %b", i_dq_freeze_n_hv);
   $fdisplay(fd, "ana_vref_in = %b", ana_vref_in);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_33 = %b", i_dqs_rdqs_pi_0_cfg[33]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_32 = %b", i_dqs_rdqs_pi_0_cfg[32]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_31 = %b", i_dqs_rdqs_pi_0_cfg[31]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_30 = %b", i_dqs_rdqs_pi_0_cfg[30]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_29 = %b", i_dqs_rdqs_pi_0_cfg[29]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_28 = %b", i_dqs_rdqs_pi_0_cfg[28]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_27 = %b", i_dqs_rdqs_pi_0_cfg[27]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_26 = %b", i_dqs_rdqs_pi_0_cfg[26]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_25 = %b", i_dqs_rdqs_pi_0_cfg[25]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_24 = %b", i_dqs_rdqs_pi_0_cfg[24]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_23 = %b", i_dqs_rdqs_pi_0_cfg[23]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_22 = %b", i_dqs_rdqs_pi_0_cfg[22]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_21 = %b", i_dqs_rdqs_pi_0_cfg[21]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_20 = %b", i_dqs_rdqs_pi_0_cfg[20]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_19 = %b", i_dqs_rdqs_pi_0_cfg[19]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_18 = %b", i_dqs_rdqs_pi_0_cfg[18]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_17 = %b", i_dqs_rdqs_pi_0_cfg[17]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_16 = %b", i_dqs_rdqs_pi_0_cfg[16]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_14 = %b", i_dqs_rdqs_pi_0_cfg[14]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_13 = %b", i_dqs_rdqs_pi_0_cfg[13]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_12 = %b", i_dqs_rdqs_pi_0_cfg[12]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_11 = %b", i_dqs_rdqs_pi_0_cfg[11]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_10 = %b", i_dqs_rdqs_pi_0_cfg[10]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_9 = %b", i_dqs_rdqs_pi_0_cfg[9]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_8 = %b", i_dqs_rdqs_pi_0_cfg[8]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_7 = %b", i_dqs_rdqs_pi_0_cfg[7]);
   $fdisplay(fd, "i_dqs_rdqs_pi_0_cfg_6 = %b", i_dqs_rdqs_pi_0_cfg[6]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_33 = %b", i_dqs_rcs_pi_cfg[33]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_32 = %b", i_dqs_rcs_pi_cfg[32]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_31 = %b", i_dqs_rcs_pi_cfg[31]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_30 = %b", i_dqs_rcs_pi_cfg[30]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_29 = %b", i_dqs_rcs_pi_cfg[29]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_28 = %b", i_dqs_rcs_pi_cfg[28]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_27 = %b", i_dqs_rcs_pi_cfg[27]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_26 = %b", i_dqs_rcs_pi_cfg[26]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_25 = %b", i_dqs_rcs_pi_cfg[25]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_24 = %b", i_dqs_rcs_pi_cfg[24]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_23 = %b", i_dqs_rcs_pi_cfg[23]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_22 = %b", i_dqs_rcs_pi_cfg[22]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_21 = %b", i_dqs_rcs_pi_cfg[21]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_20 = %b", i_dqs_rcs_pi_cfg[20]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_19 = %b", i_dqs_rcs_pi_cfg[19]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_18 = %b", i_dqs_rcs_pi_cfg[18]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_17 = %b", i_dqs_rcs_pi_cfg[17]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_16 = %b", i_dqs_rcs_pi_cfg[16]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_14 = %b", i_dqs_rcs_pi_cfg[14]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_13 = %b", i_dqs_rcs_pi_cfg[13]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_12 = %b", i_dqs_rcs_pi_cfg[12]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_11 = %b", i_dqs_rcs_pi_cfg[11]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_10 = %b", i_dqs_rcs_pi_cfg[10]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_9 = %b", i_dqs_rcs_pi_cfg[9]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_8 = %b", i_dqs_rcs_pi_cfg[8]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_7 = %b", i_dqs_rcs_pi_cfg[7]);
   $fdisplay(fd, "i_dqs_rcs_pi_cfg_6 = %b", i_dqs_rcs_pi_cfg[6]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_33 = %b", i_dqs_ren_pi_cfg[33]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_32 = %b", i_dqs_ren_pi_cfg[32]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_31 = %b", i_dqs_ren_pi_cfg[31]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_30 = %b", i_dqs_ren_pi_cfg[30]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_29 = %b", i_dqs_ren_pi_cfg[29]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_28 = %b", i_dqs_ren_pi_cfg[28]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_27 = %b", i_dqs_ren_pi_cfg[27]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_26 = %b", i_dqs_ren_pi_cfg[26]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_25 = %b", i_dqs_ren_pi_cfg[25]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_24 = %b", i_dqs_ren_pi_cfg[24]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_23 = %b", i_dqs_ren_pi_cfg[23]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_22 = %b", i_dqs_ren_pi_cfg[22]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_21 = %b", i_dqs_ren_pi_cfg[21]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_20 = %b", i_dqs_ren_pi_cfg[20]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_19 = %b", i_dqs_ren_pi_cfg[19]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_18 = %b", i_dqs_ren_pi_cfg[18]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_17 = %b", i_dqs_ren_pi_cfg[17]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_16 = %b", i_dqs_ren_pi_cfg[16]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_14 = %b", i_dqs_ren_pi_cfg[14]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_13 = %b", i_dqs_ren_pi_cfg[13]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_12 = %b", i_dqs_ren_pi_cfg[12]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_11 = %b", i_dqs_ren_pi_cfg[11]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_10 = %b", i_dqs_ren_pi_cfg[10]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_9 = %b", i_dqs_ren_pi_cfg[9]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_8 = %b", i_dqs_ren_pi_cfg[8]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_7 = %b", i_dqs_ren_pi_cfg[7]);
   $fdisplay(fd, "i_dqs_ren_pi_cfg_6 = %b", i_dqs_ren_pi_cfg[6]);
   $fdisplay(fd, "i_dqs_pre_filter_sel_1 = %b", i_dqs_pre_filter_sel[1]);
   $fdisplay(fd, "i_dqs_pre_filter_sel_0 = %b", i_dqs_pre_filter_sel[0]);
   $fdisplay(fd, "i_dqs_wck_mode = %b", i_dqs_wck_mode);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_8 = %b", i_dqs_sdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_7 = %b", i_dqs_sdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_6 = %b", i_dqs_sdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_5 = %b", i_dqs_sdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_4 = %b", i_dqs_sdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_3 = %b", i_dqs_sdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_2 = %b", i_dqs_sdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_1 = %b", i_dqs_sdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_0 = %b", i_dqs_sdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dqs_rgb_mode_7 = %b", i_dqs_rgb_mode[7]);
   $fdisplay(fd, "i_dqs_rgb_mode_6 = %b", i_dqs_rgb_mode[6]);
   $fdisplay(fd, "i_dqs_rgb_mode_5 = %b", i_dqs_rgb_mode[5]);
   $fdisplay(fd, "i_dqs_rgb_mode_4 = %b", i_dqs_rgb_mode[4]);
   $fdisplay(fd, "i_dqs_rgb_mode_3 = %b", i_dqs_rgb_mode[3]);
   $fdisplay(fd, "i_dqs_rgb_mode_2 = %b", i_dqs_rgb_mode[2]);
   $fdisplay(fd, "i_dqs_rgb_mode_1 = %b", i_dqs_rgb_mode[1]);
   $fdisplay(fd, "i_dqs_rgb_mode_0 = %b", i_dqs_rgb_mode[0]);
   $fdisplay(fd, "i_dqs_sdr_71 = %b", i_dqs_sdr[71]);
   $fdisplay(fd, "i_dqs_sdr_70 = %b", i_dqs_sdr[70]);
   $fdisplay(fd, "i_dqs_sdr_69 = %b", i_dqs_sdr[69]);
   $fdisplay(fd, "i_dqs_sdr_68 = %b", i_dqs_sdr[68]);
   $fdisplay(fd, "i_dqs_sdr_67 = %b", i_dqs_sdr[67]);
   $fdisplay(fd, "i_dqs_sdr_66 = %b", i_dqs_sdr[66]);
   $fdisplay(fd, "i_dqs_sdr_65 = %b", i_dqs_sdr[65]);
   $fdisplay(fd, "i_dqs_sdr_64 = %b", i_dqs_sdr[64]);
   $fdisplay(fd, "i_dqs_sdr_63 = %b", i_dqs_sdr[63]);
   $fdisplay(fd, "i_dqs_sdr_62 = %b", i_dqs_sdr[62]);
   $fdisplay(fd, "i_dqs_sdr_61 = %b", i_dqs_sdr[61]);
   $fdisplay(fd, "i_dqs_sdr_60 = %b", i_dqs_sdr[60]);
   $fdisplay(fd, "i_dqs_sdr_59 = %b", i_dqs_sdr[59]);
   $fdisplay(fd, "i_dqs_sdr_58 = %b", i_dqs_sdr[58]);
   $fdisplay(fd, "i_dqs_sdr_57 = %b", i_dqs_sdr[57]);
   $fdisplay(fd, "i_dqs_sdr_56 = %b", i_dqs_sdr[56]);
   $fdisplay(fd, "i_dqs_sdr_55 = %b", i_dqs_sdr[55]);
   $fdisplay(fd, "i_dqs_sdr_54 = %b", i_dqs_sdr[54]);
   $fdisplay(fd, "i_dqs_sdr_53 = %b", i_dqs_sdr[53]);
   $fdisplay(fd, "i_dqs_sdr_52 = %b", i_dqs_sdr[52]);
   $fdisplay(fd, "i_dqs_sdr_51 = %b", i_dqs_sdr[51]);
   $fdisplay(fd, "i_dqs_sdr_50 = %b", i_dqs_sdr[50]);
   $fdisplay(fd, "i_dqs_sdr_49 = %b", i_dqs_sdr[49]);
   $fdisplay(fd, "i_dqs_sdr_48 = %b", i_dqs_sdr[48]);
   $fdisplay(fd, "i_dqs_sdr_47 = %b", i_dqs_sdr[47]);
   $fdisplay(fd, "i_dqs_sdr_46 = %b", i_dqs_sdr[46]);
   $fdisplay(fd, "i_dqs_sdr_45 = %b", i_dqs_sdr[45]);
   $fdisplay(fd, "i_dqs_sdr_44 = %b", i_dqs_sdr[44]);
   $fdisplay(fd, "i_dqs_sdr_43 = %b", i_dqs_sdr[43]);
   $fdisplay(fd, "i_dqs_sdr_42 = %b", i_dqs_sdr[42]);
   $fdisplay(fd, "i_dqs_sdr_41 = %b", i_dqs_sdr[41]);
   $fdisplay(fd, "i_dqs_sdr_40 = %b", i_dqs_sdr[40]);
   $fdisplay(fd, "i_dqs_sdr_39 = %b", i_dqs_sdr[39]);
   $fdisplay(fd, "i_dqs_sdr_38 = %b", i_dqs_sdr[38]);
   $fdisplay(fd, "i_dqs_sdr_37 = %b", i_dqs_sdr[37]);
   $fdisplay(fd, "i_dqs_sdr_36 = %b", i_dqs_sdr[36]);
   $fdisplay(fd, "i_dqs_sdr_35 = %b", i_dqs_sdr[35]);
   $fdisplay(fd, "i_dqs_sdr_34 = %b", i_dqs_sdr[34]);
   $fdisplay(fd, "i_dqs_sdr_33 = %b", i_dqs_sdr[33]);
   $fdisplay(fd, "i_dqs_sdr_32 = %b", i_dqs_sdr[32]);
   $fdisplay(fd, "i_dqs_sdr_31 = %b", i_dqs_sdr[31]);
   $fdisplay(fd, "i_dqs_sdr_30 = %b", i_dqs_sdr[30]);
   $fdisplay(fd, "i_dqs_sdr_29 = %b", i_dqs_sdr[29]);
   $fdisplay(fd, "i_dqs_sdr_28 = %b", i_dqs_sdr[28]);
   $fdisplay(fd, "i_dqs_sdr_27 = %b", i_dqs_sdr[27]);
   $fdisplay(fd, "i_dqs_sdr_26 = %b", i_dqs_sdr[26]);
   $fdisplay(fd, "i_dqs_sdr_25 = %b", i_dqs_sdr[25]);
   $fdisplay(fd, "i_dqs_sdr_24 = %b", i_dqs_sdr[24]);
   $fdisplay(fd, "i_dqs_sdr_23 = %b", i_dqs_sdr[23]);
   $fdisplay(fd, "i_dqs_sdr_22 = %b", i_dqs_sdr[22]);
   $fdisplay(fd, "i_dqs_sdr_21 = %b", i_dqs_sdr[21]);
   $fdisplay(fd, "i_dqs_sdr_20 = %b", i_dqs_sdr[20]);
   $fdisplay(fd, "i_dqs_sdr_19 = %b", i_dqs_sdr[19]);
   $fdisplay(fd, "i_dqs_sdr_18 = %b", i_dqs_sdr[18]);
   $fdisplay(fd, "i_dqs_sdr_17 = %b", i_dqs_sdr[17]);
   $fdisplay(fd, "i_dqs_sdr_16 = %b", i_dqs_sdr[16]);
   $fdisplay(fd, "i_dqs_sdr_15 = %b", i_dqs_sdr[15]);
   $fdisplay(fd, "i_dqs_sdr_14 = %b", i_dqs_sdr[14]);
   $fdisplay(fd, "i_dqs_sdr_13 = %b", i_dqs_sdr[13]);
   $fdisplay(fd, "i_dqs_sdr_12 = %b", i_dqs_sdr[12]);
   $fdisplay(fd, "i_dqs_sdr_11 = %b", i_dqs_sdr[11]);
   $fdisplay(fd, "i_dqs_sdr_10 = %b", i_dqs_sdr[10]);
   $fdisplay(fd, "i_dqs_sdr_9 = %b", i_dqs_sdr[9]);
   $fdisplay(fd, "i_dqs_sdr_8 = %b", i_dqs_sdr[8]);
   $fdisplay(fd, "i_dqs_sdr_7 = %b", i_dqs_sdr[7]);
   $fdisplay(fd, "i_dqs_sdr_6 = %b", i_dqs_sdr[6]);
   $fdisplay(fd, "i_dqs_sdr_5 = %b", i_dqs_sdr[5]);
   $fdisplay(fd, "i_dqs_sdr_4 = %b", i_dqs_sdr[4]);
   $fdisplay(fd, "i_dqs_sdr_3 = %b", i_dqs_sdr[3]);
   $fdisplay(fd, "i_dqs_sdr_2 = %b", i_dqs_sdr[2]);
   $fdisplay(fd, "i_dqs_sdr_1 = %b", i_dqs_sdr[1]);
   $fdisplay(fd, "i_dqs_sdr_0 = %b", i_dqs_sdr[0]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_33 = %b", i_dqs_sdr_rt_pi_cfg[33]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_32 = %b", i_dqs_sdr_rt_pi_cfg[32]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_31 = %b", i_dqs_sdr_rt_pi_cfg[31]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_30 = %b", i_dqs_sdr_rt_pi_cfg[30]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_29 = %b", i_dqs_sdr_rt_pi_cfg[29]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_28 = %b", i_dqs_sdr_rt_pi_cfg[28]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_27 = %b", i_dqs_sdr_rt_pi_cfg[27]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_26 = %b", i_dqs_sdr_rt_pi_cfg[26]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_25 = %b", i_dqs_sdr_rt_pi_cfg[25]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_24 = %b", i_dqs_sdr_rt_pi_cfg[24]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_23 = %b", i_dqs_sdr_rt_pi_cfg[23]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_22 = %b", i_dqs_sdr_rt_pi_cfg[22]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_21 = %b", i_dqs_sdr_rt_pi_cfg[21]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_20 = %b", i_dqs_sdr_rt_pi_cfg[20]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_19 = %b", i_dqs_sdr_rt_pi_cfg[19]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_18 = %b", i_dqs_sdr_rt_pi_cfg[18]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_17 = %b", i_dqs_sdr_rt_pi_cfg[17]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_16 = %b", i_dqs_sdr_rt_pi_cfg[16]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_14 = %b", i_dqs_sdr_rt_pi_cfg[14]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_13 = %b", i_dqs_sdr_rt_pi_cfg[13]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_12 = %b", i_dqs_sdr_rt_pi_cfg[12]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_11 = %b", i_dqs_sdr_rt_pi_cfg[11]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_10 = %b", i_dqs_sdr_rt_pi_cfg[10]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_9 = %b", i_dqs_sdr_rt_pi_cfg[9]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_8 = %b", i_dqs_sdr_rt_pi_cfg[8]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_7 = %b", i_dqs_sdr_rt_pi_cfg[7]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_6 = %b", i_dqs_sdr_rt_pi_cfg[6]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_33 = %b", i_dqs_ddr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_32 = %b", i_dqs_ddr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_31 = %b", i_dqs_ddr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_30 = %b", i_dqs_ddr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_29 = %b", i_dqs_ddr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_28 = %b", i_dqs_ddr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_27 = %b", i_dqs_ddr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_26 = %b", i_dqs_ddr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_25 = %b", i_dqs_ddr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_24 = %b", i_dqs_ddr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_23 = %b", i_dqs_ddr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_22 = %b", i_dqs_ddr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_21 = %b", i_dqs_ddr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_20 = %b", i_dqs_ddr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_19 = %b", i_dqs_ddr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_18 = %b", i_dqs_ddr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_17 = %b", i_dqs_ddr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_16 = %b", i_dqs_ddr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_14 = %b", i_dqs_ddr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_13 = %b", i_dqs_ddr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_12 = %b", i_dqs_ddr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_11 = %b", i_dqs_ddr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_10 = %b", i_dqs_ddr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_9 = %b", i_dqs_ddr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_8 = %b", i_dqs_ddr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_7 = %b", i_dqs_ddr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_6 = %b", i_dqs_ddr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_33 = %b", i_dqs_qdr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_32 = %b", i_dqs_qdr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_31 = %b", i_dqs_qdr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_30 = %b", i_dqs_qdr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_29 = %b", i_dqs_qdr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_28 = %b", i_dqs_qdr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_27 = %b", i_dqs_qdr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_26 = %b", i_dqs_qdr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_25 = %b", i_dqs_qdr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_24 = %b", i_dqs_qdr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_23 = %b", i_dqs_qdr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_22 = %b", i_dqs_qdr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_21 = %b", i_dqs_qdr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_20 = %b", i_dqs_qdr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_19 = %b", i_dqs_qdr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_18 = %b", i_dqs_qdr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_17 = %b", i_dqs_qdr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_16 = %b", i_dqs_qdr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_14 = %b", i_dqs_qdr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_13 = %b", i_dqs_qdr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_12 = %b", i_dqs_qdr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_11 = %b", i_dqs_qdr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_10 = %b", i_dqs_qdr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_9 = %b", i_dqs_qdr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_8 = %b", i_dqs_qdr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_7 = %b", i_dqs_qdr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_6 = %b", i_dqs_qdr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_17 = %b", i_dqs_xdr_lpde_cfg[17]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_16 = %b", i_dqs_xdr_lpde_cfg[16]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_15 = %b", i_dqs_xdr_lpde_cfg[15]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_14 = %b", i_dqs_xdr_lpde_cfg[14]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_13 = %b", i_dqs_xdr_lpde_cfg[13]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_12 = %b", i_dqs_xdr_lpde_cfg[12]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_11 = %b", i_dqs_xdr_lpde_cfg[11]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_10 = %b", i_dqs_xdr_lpde_cfg[10]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_9 = %b", i_dqs_xdr_lpde_cfg[9]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_8 = %b", i_dqs_xdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_7 = %b", i_dqs_xdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_6 = %b", i_dqs_xdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_5 = %b", i_dqs_xdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_4 = %b", i_dqs_xdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_3 = %b", i_dqs_xdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_2 = %b", i_dqs_xdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_1 = %b", i_dqs_xdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_0 = %b", i_dqs_xdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_8 = %b", i_dqs_ddr_1_pipe_en[8]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_7 = %b", i_dqs_ddr_1_pipe_en[7]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_6 = %b", i_dqs_ddr_1_pipe_en[6]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_5 = %b", i_dqs_ddr_1_pipe_en[5]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_4 = %b", i_dqs_ddr_1_pipe_en[4]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_3 = %b", i_dqs_ddr_1_pipe_en[3]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_2 = %b", i_dqs_ddr_1_pipe_en[2]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_1 = %b", i_dqs_ddr_1_pipe_en[1]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_0 = %b", i_dqs_ddr_1_pipe_en[0]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_16 = %b", i_dqs_ddr_1_x_sel[16]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_14 = %b", i_dqs_ddr_1_x_sel[14]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_12 = %b", i_dqs_ddr_1_x_sel[12]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_10 = %b", i_dqs_ddr_1_x_sel[10]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_8 = %b", i_dqs_ddr_1_x_sel[8]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_6 = %b", i_dqs_ddr_1_x_sel[6]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_4 = %b", i_dqs_ddr_1_x_sel[4]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_2 = %b", i_dqs_ddr_1_x_sel[2]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_0 = %b", i_dqs_ddr_1_x_sel[0]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_8 = %b", i_dqs_ddr_0_pipe_en[8]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_7 = %b", i_dqs_ddr_0_pipe_en[7]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_6 = %b", i_dqs_ddr_0_pipe_en[6]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_5 = %b", i_dqs_ddr_0_pipe_en[5]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_4 = %b", i_dqs_ddr_0_pipe_en[4]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_3 = %b", i_dqs_ddr_0_pipe_en[3]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_2 = %b", i_dqs_ddr_0_pipe_en[2]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_1 = %b", i_dqs_ddr_0_pipe_en[1]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_0 = %b", i_dqs_ddr_0_pipe_en[0]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_16 = %b", i_dqs_ddr_0_x_sel[16]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_14 = %b", i_dqs_ddr_0_x_sel[14]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_12 = %b", i_dqs_ddr_0_x_sel[12]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_10 = %b", i_dqs_ddr_0_x_sel[10]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_8 = %b", i_dqs_ddr_0_x_sel[8]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_6 = %b", i_dqs_ddr_0_x_sel[6]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_4 = %b", i_dqs_ddr_0_x_sel[4]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_2 = %b", i_dqs_ddr_0_x_sel[2]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_0 = %b", i_dqs_ddr_0_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_8 = %b", i_dqs_sdr_3_pipe_en[8]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_7 = %b", i_dqs_sdr_3_pipe_en[7]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_6 = %b", i_dqs_sdr_3_pipe_en[6]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_5 = %b", i_dqs_sdr_3_pipe_en[5]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_4 = %b", i_dqs_sdr_3_pipe_en[4]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_3 = %b", i_dqs_sdr_3_pipe_en[3]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_2 = %b", i_dqs_sdr_3_pipe_en[2]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_1 = %b", i_dqs_sdr_3_pipe_en[1]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_0 = %b", i_dqs_sdr_3_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_25 = %b", i_dqs_sdr_3_x_sel[25]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_24 = %b", i_dqs_sdr_3_x_sel[24]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_22 = %b", i_dqs_sdr_3_x_sel[22]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_21 = %b", i_dqs_sdr_3_x_sel[21]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_19 = %b", i_dqs_sdr_3_x_sel[19]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_18 = %b", i_dqs_sdr_3_x_sel[18]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_16 = %b", i_dqs_sdr_3_x_sel[16]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_15 = %b", i_dqs_sdr_3_x_sel[15]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_13 = %b", i_dqs_sdr_3_x_sel[13]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_12 = %b", i_dqs_sdr_3_x_sel[12]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_10 = %b", i_dqs_sdr_3_x_sel[10]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_9 = %b", i_dqs_sdr_3_x_sel[9]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_7 = %b", i_dqs_sdr_3_x_sel[7]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_6 = %b", i_dqs_sdr_3_x_sel[6]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_4 = %b", i_dqs_sdr_3_x_sel[4]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_3 = %b", i_dqs_sdr_3_x_sel[3]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_1 = %b", i_dqs_sdr_3_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_0 = %b", i_dqs_sdr_3_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_17 = %b", i_dqs_sdr_3_fc_dly[17]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_16 = %b", i_dqs_sdr_3_fc_dly[16]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_15 = %b", i_dqs_sdr_3_fc_dly[15]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_14 = %b", i_dqs_sdr_3_fc_dly[14]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_13 = %b", i_dqs_sdr_3_fc_dly[13]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_12 = %b", i_dqs_sdr_3_fc_dly[12]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_11 = %b", i_dqs_sdr_3_fc_dly[11]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_10 = %b", i_dqs_sdr_3_fc_dly[10]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_9 = %b", i_dqs_sdr_3_fc_dly[9]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_8 = %b", i_dqs_sdr_3_fc_dly[8]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_7 = %b", i_dqs_sdr_3_fc_dly[7]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_6 = %b", i_dqs_sdr_3_fc_dly[6]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_5 = %b", i_dqs_sdr_3_fc_dly[5]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_4 = %b", i_dqs_sdr_3_fc_dly[4]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_3 = %b", i_dqs_sdr_3_fc_dly[3]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_2 = %b", i_dqs_sdr_3_fc_dly[2]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_1 = %b", i_dqs_sdr_3_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_0 = %b", i_dqs_sdr_3_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_8 = %b", i_dqs_sdr_2_pipe_en[8]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_7 = %b", i_dqs_sdr_2_pipe_en[7]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_6 = %b", i_dqs_sdr_2_pipe_en[6]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_5 = %b", i_dqs_sdr_2_pipe_en[5]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_4 = %b", i_dqs_sdr_2_pipe_en[4]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_3 = %b", i_dqs_sdr_2_pipe_en[3]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_2 = %b", i_dqs_sdr_2_pipe_en[2]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_1 = %b", i_dqs_sdr_2_pipe_en[1]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_0 = %b", i_dqs_sdr_2_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_25 = %b", i_dqs_sdr_2_x_sel[25]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_24 = %b", i_dqs_sdr_2_x_sel[24]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_22 = %b", i_dqs_sdr_2_x_sel[22]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_21 = %b", i_dqs_sdr_2_x_sel[21]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_19 = %b", i_dqs_sdr_2_x_sel[19]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_18 = %b", i_dqs_sdr_2_x_sel[18]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_16 = %b", i_dqs_sdr_2_x_sel[16]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_15 = %b", i_dqs_sdr_2_x_sel[15]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_13 = %b", i_dqs_sdr_2_x_sel[13]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_12 = %b", i_dqs_sdr_2_x_sel[12]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_10 = %b", i_dqs_sdr_2_x_sel[10]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_9 = %b", i_dqs_sdr_2_x_sel[9]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_7 = %b", i_dqs_sdr_2_x_sel[7]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_6 = %b", i_dqs_sdr_2_x_sel[6]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_4 = %b", i_dqs_sdr_2_x_sel[4]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_3 = %b", i_dqs_sdr_2_x_sel[3]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_1 = %b", i_dqs_sdr_2_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_0 = %b", i_dqs_sdr_2_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_17 = %b", i_dqs_sdr_2_fc_dly[17]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_16 = %b", i_dqs_sdr_2_fc_dly[16]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_15 = %b", i_dqs_sdr_2_fc_dly[15]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_14 = %b", i_dqs_sdr_2_fc_dly[14]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_13 = %b", i_dqs_sdr_2_fc_dly[13]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_12 = %b", i_dqs_sdr_2_fc_dly[12]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_11 = %b", i_dqs_sdr_2_fc_dly[11]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_10 = %b", i_dqs_sdr_2_fc_dly[10]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_9 = %b", i_dqs_sdr_2_fc_dly[9]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_8 = %b", i_dqs_sdr_2_fc_dly[8]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_7 = %b", i_dqs_sdr_2_fc_dly[7]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_6 = %b", i_dqs_sdr_2_fc_dly[6]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_5 = %b", i_dqs_sdr_2_fc_dly[5]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_4 = %b", i_dqs_sdr_2_fc_dly[4]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_3 = %b", i_dqs_sdr_2_fc_dly[3]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_2 = %b", i_dqs_sdr_2_fc_dly[2]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_1 = %b", i_dqs_sdr_2_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_0 = %b", i_dqs_sdr_2_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_8 = %b", i_dqs_sdr_1_pipe_en[8]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_7 = %b", i_dqs_sdr_1_pipe_en[7]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_6 = %b", i_dqs_sdr_1_pipe_en[6]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_5 = %b", i_dqs_sdr_1_pipe_en[5]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_4 = %b", i_dqs_sdr_1_pipe_en[4]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_3 = %b", i_dqs_sdr_1_pipe_en[3]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_2 = %b", i_dqs_sdr_1_pipe_en[2]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_1 = %b", i_dqs_sdr_1_pipe_en[1]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_0 = %b", i_dqs_sdr_1_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_25 = %b", i_dqs_sdr_1_x_sel[25]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_24 = %b", i_dqs_sdr_1_x_sel[24]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_22 = %b", i_dqs_sdr_1_x_sel[22]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_21 = %b", i_dqs_sdr_1_x_sel[21]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_19 = %b", i_dqs_sdr_1_x_sel[19]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_18 = %b", i_dqs_sdr_1_x_sel[18]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_16 = %b", i_dqs_sdr_1_x_sel[16]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_15 = %b", i_dqs_sdr_1_x_sel[15]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_13 = %b", i_dqs_sdr_1_x_sel[13]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_12 = %b", i_dqs_sdr_1_x_sel[12]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_10 = %b", i_dqs_sdr_1_x_sel[10]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_9 = %b", i_dqs_sdr_1_x_sel[9]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_7 = %b", i_dqs_sdr_1_x_sel[7]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_6 = %b", i_dqs_sdr_1_x_sel[6]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_4 = %b", i_dqs_sdr_1_x_sel[4]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_3 = %b", i_dqs_sdr_1_x_sel[3]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_1 = %b", i_dqs_sdr_1_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_0 = %b", i_dqs_sdr_1_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_17 = %b", i_dqs_sdr_1_fc_dly[17]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_16 = %b", i_dqs_sdr_1_fc_dly[16]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_15 = %b", i_dqs_sdr_1_fc_dly[15]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_14 = %b", i_dqs_sdr_1_fc_dly[14]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_13 = %b", i_dqs_sdr_1_fc_dly[13]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_12 = %b", i_dqs_sdr_1_fc_dly[12]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_11 = %b", i_dqs_sdr_1_fc_dly[11]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_10 = %b", i_dqs_sdr_1_fc_dly[10]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_9 = %b", i_dqs_sdr_1_fc_dly[9]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_8 = %b", i_dqs_sdr_1_fc_dly[8]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_7 = %b", i_dqs_sdr_1_fc_dly[7]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_6 = %b", i_dqs_sdr_1_fc_dly[6]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_5 = %b", i_dqs_sdr_1_fc_dly[5]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_4 = %b", i_dqs_sdr_1_fc_dly[4]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_3 = %b", i_dqs_sdr_1_fc_dly[3]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_2 = %b", i_dqs_sdr_1_fc_dly[2]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_1 = %b", i_dqs_sdr_1_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_0 = %b", i_dqs_sdr_1_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_8 = %b", i_dqs_sdr_0_pipe_en[8]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_7 = %b", i_dqs_sdr_0_pipe_en[7]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_6 = %b", i_dqs_sdr_0_pipe_en[6]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_5 = %b", i_dqs_sdr_0_pipe_en[5]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_4 = %b", i_dqs_sdr_0_pipe_en[4]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_3 = %b", i_dqs_sdr_0_pipe_en[3]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_2 = %b", i_dqs_sdr_0_pipe_en[2]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_1 = %b", i_dqs_sdr_0_pipe_en[1]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_0 = %b", i_dqs_sdr_0_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_25 = %b", i_dqs_sdr_0_x_sel[25]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_24 = %b", i_dqs_sdr_0_x_sel[24]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_22 = %b", i_dqs_sdr_0_x_sel[22]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_21 = %b", i_dqs_sdr_0_x_sel[21]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_19 = %b", i_dqs_sdr_0_x_sel[19]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_18 = %b", i_dqs_sdr_0_x_sel[18]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_16 = %b", i_dqs_sdr_0_x_sel[16]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_15 = %b", i_dqs_sdr_0_x_sel[15]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_13 = %b", i_dqs_sdr_0_x_sel[13]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_12 = %b", i_dqs_sdr_0_x_sel[12]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_10 = %b", i_dqs_sdr_0_x_sel[10]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_9 = %b", i_dqs_sdr_0_x_sel[9]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_7 = %b", i_dqs_sdr_0_x_sel[7]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_6 = %b", i_dqs_sdr_0_x_sel[6]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_4 = %b", i_dqs_sdr_0_x_sel[4]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_3 = %b", i_dqs_sdr_0_x_sel[3]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_1 = %b", i_dqs_sdr_0_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_0 = %b", i_dqs_sdr_0_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_17 = %b", i_dqs_sdr_0_fc_dly[17]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_16 = %b", i_dqs_sdr_0_fc_dly[16]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_15 = %b", i_dqs_sdr_0_fc_dly[15]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_14 = %b", i_dqs_sdr_0_fc_dly[14]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_13 = %b", i_dqs_sdr_0_fc_dly[13]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_12 = %b", i_dqs_sdr_0_fc_dly[12]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_11 = %b", i_dqs_sdr_0_fc_dly[11]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_10 = %b", i_dqs_sdr_0_fc_dly[10]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_9 = %b", i_dqs_sdr_0_fc_dly[9]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_8 = %b", i_dqs_sdr_0_fc_dly[8]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_7 = %b", i_dqs_sdr_0_fc_dly[7]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_6 = %b", i_dqs_sdr_0_fc_dly[6]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_5 = %b", i_dqs_sdr_0_fc_dly[5]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_4 = %b", i_dqs_sdr_0_fc_dly[4]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_3 = %b", i_dqs_sdr_0_fc_dly[3]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_2 = %b", i_dqs_sdr_0_fc_dly[2]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_1 = %b", i_dqs_sdr_0_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_0 = %b", i_dqs_sdr_0_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_8 = %b", i_dqs_sdr_rt_pipe_en[8]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_7 = %b", i_dqs_sdr_rt_pipe_en[7]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_6 = %b", i_dqs_sdr_rt_pipe_en[6]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_5 = %b", i_dqs_sdr_rt_pipe_en[5]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_4 = %b", i_dqs_sdr_rt_pipe_en[4]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_3 = %b", i_dqs_sdr_rt_pipe_en[3]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_2 = %b", i_dqs_sdr_rt_pipe_en[2]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_1 = %b", i_dqs_sdr_rt_pipe_en[1]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_0 = %b", i_dqs_sdr_rt_pipe_en[0]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_3 = %b", i_dfirdclk_en_pulse_ext[3]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_2 = %b", i_dfirdclk_en_pulse_ext[2]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_1 = %b", i_dfirdclk_en_pulse_ext[1]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_0 = %b", i_dfirdclk_en_pulse_ext[0]);
   $fdisplay(fd, "i_dfirdclk_en = %b", i_dfirdclk_en);
   $fdisplay(fd, "i_dq_dfi_wrtraffic = %b", i_dq_dfi_wrtraffic);
   $fdisplay(fd, "i_dqs_dfi_wrtraffic = %b", i_dqs_dfi_wrtraffic);
   $fdisplay(fd, "i_csp_div_rst_n %b", i_csp_div_rst_n);
   $fdisplay(fd, "i_dqs_ck2wck_ratio_2 = %b", i_dqs_ck2wck_ratio[2]);
   $fdisplay(fd, "i_dqs_ck2wck_ratio_1 = %b", i_dqs_ck2wck_ratio[1]);
   $fdisplay(fd, "i_dqs_wgb_mode_8 = %b", i_dqs_wgb_mode[8]);
   $fdisplay(fd, "i_dqs_tgb_mode_7 = %b", i_dqs_tgb_mode[7]);
   $fdisplay(fd, "i_dqs_tgb_mode_6 = %b", i_dqs_tgb_mode[6]);
   $fdisplay(fd, "i_dqs_tgb_mode_4 = %b", i_dqs_tgb_mode[4]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_62 = %b", i_dqs_egress_mode_dig[62]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_57 = %b", i_dqs_egress_mode_dig[57]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_56 = %b", i_dqs_egress_mode_dig[56]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_55 = %b", i_dqs_egress_mode_dig[55]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_50 = %b", i_dqs_egress_mode_dig[50]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_49 = %b", i_dqs_egress_mode_dig[49]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_48 = %b", i_dqs_egress_mode_dig[48]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_43 = %b", i_dqs_egress_mode_dig[43]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_42 = %b", i_dqs_egress_mode_dig[42]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_41 = %b", i_dqs_egress_mode_dig[41]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_36 = %b", i_dqs_egress_mode_dig[36]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_35 = %b", i_dqs_egress_mode_dig[35]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_34 = %b", i_dqs_egress_mode_dig[34]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_29 = %b", i_dqs_egress_mode_dig[29]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_28 = %b", i_dqs_egress_mode_dig[28]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_27 = %b", i_dqs_egress_mode_dig[27]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_22 = %b", i_dqs_egress_mode_dig[22]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_21 = %b", i_dqs_egress_mode_dig[21]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_20 = %b", i_dqs_egress_mode_dig[20]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_15 = %b", i_dqs_egress_mode_dig[15]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_14 = %b", i_dqs_egress_mode_dig[14]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_13 = %b", i_dqs_egress_mode_dig[13]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_8 = %b", i_dqs_egress_mode_dig[8]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_7 = %b", i_dqs_egress_mode_dig[7]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_6 = %b", i_dqs_egress_mode_dig[6]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_1 = %b", i_dqs_egress_mode_dig[1]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_0 = %b", i_dqs_egress_mode_dig[0]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_50 = %b", i_dqs_egress_mode_ana[50]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_49 = %b", i_dqs_egress_mode_ana[49]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_48 = %b", i_dqs_egress_mode_ana[48]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_44 = %b", i_dqs_egress_mode_ana[44]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_43 = %b", i_dqs_egress_mode_ana[43]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_42 = %b", i_dqs_egress_mode_ana[42]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_38 = %b", i_dqs_egress_mode_ana[38]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_37 = %b", i_dqs_egress_mode_ana[37]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_36 = %b", i_dqs_egress_mode_ana[36]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_32 = %b", i_dqs_egress_mode_ana[32]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_31 = %b", i_dqs_egress_mode_ana[31]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_30 = %b", i_dqs_egress_mode_ana[30]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_26 = %b", i_dqs_egress_mode_ana[26]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_25 = %b", i_dqs_egress_mode_ana[25]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_24 = %b", i_dqs_egress_mode_ana[24]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_20 = %b", i_dqs_egress_mode_ana[20]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_19 = %b", i_dqs_egress_mode_ana[19]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_18 = %b", i_dqs_egress_mode_ana[18]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_14 = %b", i_dqs_egress_mode_ana[14]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_13 = %b", i_dqs_egress_mode_ana[13]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_12 = %b", i_dqs_egress_mode_ana[12]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_8 = %b", i_dqs_egress_mode_ana[8]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_7 = %b", i_dqs_egress_mode_ana[7]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_6 = %b", i_dqs_egress_mode_ana[6]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_2 = %b", i_dqs_egress_mode_ana[2]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_1 = %b", i_dqs_egress_mode_ana[1]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_0 = %b", i_dqs_egress_mode_ana[0]);
   $fdisplay(fd, "i_dq_sdr_71 = %b", i_dq_sdr[71]);
   $fdisplay(fd, "i_dq_sdr_70 = %b", i_dq_sdr[70]);
   $fdisplay(fd, "i_dq_sdr_69 = %b", i_dq_sdr[69]);
   $fdisplay(fd, "i_dq_sdr_68 = %b", i_dq_sdr[68]);
   $fdisplay(fd, "i_dq_sdr_67 = %b", i_dq_sdr[67]);
   $fdisplay(fd, "i_dq_sdr_66 = %b", i_dq_sdr[66]);
   $fdisplay(fd, "i_dq_sdr_65 = %b", i_dq_sdr[65]);
   $fdisplay(fd, "i_dq_sdr_64 = %b", i_dq_sdr[64]);
   $fdisplay(fd, "i_dq_sdr_63 = %b", i_dq_sdr[63]);
   $fdisplay(fd, "i_dq_sdr_62 = %b", i_dq_sdr[62]);
   $fdisplay(fd, "i_dq_sdr_61 = %b", i_dq_sdr[61]);
   $fdisplay(fd, "i_dq_sdr_60 = %b", i_dq_sdr[60]);
   $fdisplay(fd, "i_dq_sdr_59 = %b", i_dq_sdr[59]);
   $fdisplay(fd, "i_dq_sdr_58 = %b", i_dq_sdr[58]);
   $fdisplay(fd, "i_dq_sdr_57 = %b", i_dq_sdr[57]);
   $fdisplay(fd, "i_dq_sdr_56 = %b", i_dq_sdr[56]);
   $fdisplay(fd, "i_dq_sdr_55 = %b", i_dq_sdr[55]);
   $fdisplay(fd, "i_dq_sdr_54 = %b", i_dq_sdr[54]);
   $fdisplay(fd, "i_dq_sdr_53 = %b", i_dq_sdr[53]);
   $fdisplay(fd, "i_dq_sdr_52 = %b", i_dq_sdr[52]);
   $fdisplay(fd, "i_dq_sdr_51 = %b", i_dq_sdr[51]);
   $fdisplay(fd, "i_dq_sdr_50 = %b", i_dq_sdr[50]);
   $fdisplay(fd, "i_dq_sdr_49 = %b", i_dq_sdr[49]);
   $fdisplay(fd, "i_dq_sdr_48 = %b", i_dq_sdr[48]);
   $fdisplay(fd, "i_dq_sdr_47 = %b", i_dq_sdr[47]);
   $fdisplay(fd, "i_dq_sdr_46 = %b", i_dq_sdr[46]);
   $fdisplay(fd, "i_dq_sdr_45 = %b", i_dq_sdr[45]);
   $fdisplay(fd, "i_dq_sdr_44 = %b", i_dq_sdr[44]);
   $fdisplay(fd, "i_dq_sdr_43 = %b", i_dq_sdr[43]);
   $fdisplay(fd, "i_dq_sdr_42 = %b", i_dq_sdr[42]);
   $fdisplay(fd, "i_dq_sdr_41 = %b", i_dq_sdr[41]);
   $fdisplay(fd, "i_dq_sdr_40 = %b", i_dq_sdr[40]);
   $fdisplay(fd, "i_dq_sdr_39 = %b", i_dq_sdr[39]);
   $fdisplay(fd, "i_dq_sdr_38 = %b", i_dq_sdr[38]);
   $fdisplay(fd, "i_dq_sdr_37 = %b", i_dq_sdr[37]);
   $fdisplay(fd, "i_dq_sdr_36 = %b", i_dq_sdr[36]);
   $fdisplay(fd, "i_dq_sdr_35 = %b", i_dq_sdr[35]);
   $fdisplay(fd, "i_dq_sdr_34 = %b", i_dq_sdr[34]);
   $fdisplay(fd, "i_dq_sdr_33 = %b", i_dq_sdr[33]);
   $fdisplay(fd, "i_dq_sdr_32 = %b", i_dq_sdr[32]);
   $fdisplay(fd, "i_dq_sdr_31 = %b", i_dq_sdr[31]);
   $fdisplay(fd, "i_dq_sdr_30 = %b", i_dq_sdr[30]);
   $fdisplay(fd, "i_dq_sdr_29 = %b", i_dq_sdr[29]);
   $fdisplay(fd, "i_dq_sdr_28 = %b", i_dq_sdr[28]);
   $fdisplay(fd, "i_dq_sdr_27 = %b", i_dq_sdr[27]);
   $fdisplay(fd, "i_dq_sdr_26 = %b", i_dq_sdr[26]);
   $fdisplay(fd, "i_dq_sdr_25 = %b", i_dq_sdr[25]);
   $fdisplay(fd, "i_dq_sdr_24 = %b", i_dq_sdr[24]);
   $fdisplay(fd, "i_dq_sdr_23 = %b", i_dq_sdr[23]);
   $fdisplay(fd, "i_dq_sdr_22 = %b", i_dq_sdr[22]);
   $fdisplay(fd, "i_dq_sdr_21 = %b", i_dq_sdr[21]);
   $fdisplay(fd, "i_dq_sdr_20 = %b", i_dq_sdr[20]);
   $fdisplay(fd, "i_dq_sdr_19 = %b", i_dq_sdr[19]);
   $fdisplay(fd, "i_dq_sdr_18 = %b", i_dq_sdr[18]);
   $fdisplay(fd, "i_dq_sdr_17 = %b", i_dq_sdr[17]);
   $fdisplay(fd, "i_dq_sdr_16 = %b", i_dq_sdr[16]);
   $fdisplay(fd, "i_dq_sdr_15 = %b", i_dq_sdr[15]);
   $fdisplay(fd, "i_dq_sdr_14 = %b", i_dq_sdr[14]);
   $fdisplay(fd, "i_dq_sdr_13 = %b", i_dq_sdr[13]);
   $fdisplay(fd, "i_dq_sdr_12 = %b", i_dq_sdr[12]);
   $fdisplay(fd, "i_dq_sdr_11 = %b", i_dq_sdr[11]);
   $fdisplay(fd, "i_dq_sdr_10 = %b", i_dq_sdr[10]);
   $fdisplay(fd, "i_dq_sdr_9 = %b", i_dq_sdr[9]);
   $fdisplay(fd, "i_dq_sdr_8 = %b", i_dq_sdr[8]);
   $fdisplay(fd, "i_dq_sdr_7 = %b", i_dq_sdr[7]);
   $fdisplay(fd, "i_dq_sdr_6 = %b", i_dq_sdr[6]);
   $fdisplay(fd, "i_dq_sdr_5 = %b", i_dq_sdr[5]);
   $fdisplay(fd, "i_dq_sdr_4 = %b", i_dq_sdr[4]);
   $fdisplay(fd, "i_dq_sdr_3 = %b", i_dq_sdr[3]);
   $fdisplay(fd, "i_dq_sdr_2 = %b", i_dq_sdr[2]);
   $fdisplay(fd, "i_dq_sdr_1 = %b", i_dq_sdr[1]);
   $fdisplay(fd, "i_dq_sdr_0 = %b", i_dq_sdr[0]);
   $fdisplay(fd, "i_dfi_pi_cfg_14 = %b", i_dfi_pi_cfg[14]);
   $fdisplay(fd, "i_dfi_pi_cfg_13 = %b", i_dfi_pi_cfg[13]);
   $fdisplay(fd, "i_dfi_pi_cfg_12 = %b", i_dfi_pi_cfg[12]);
   $fdisplay(fd, "i_dfi_pi_cfg_11 = %b", i_dfi_pi_cfg[11]);
   $fdisplay(fd, "i_dfi_pi_cfg_10 = %b", i_dfi_pi_cfg[10]);
   $fdisplay(fd, "i_dfi_pi_cfg_9 = %b", i_dfi_pi_cfg[9]);
   $fdisplay(fd, "i_dfi_pi_cfg_8 = %b", i_dfi_pi_cfg[8]);
   $fdisplay(fd, "i_dfi_pi_cfg_7 = %b", i_dfi_pi_cfg[7]);
   $fdisplay(fd, "i_dfi_pi_cfg_6 = %b", i_dfi_pi_cfg[6]);
   $fdisplay(fd, "i_sdr_pi_cfg_14 = %b", i_sdr_pi_cfg[14]);
   $fdisplay(fd, "i_sdr_pi_cfg_13 = %b", i_sdr_pi_cfg[13]);
   $fdisplay(fd, "i_sdr_pi_cfg_12 = %b", i_sdr_pi_cfg[12]);
   $fdisplay(fd, "i_sdr_pi_cfg_11 = %b", i_sdr_pi_cfg[11]);
   $fdisplay(fd, "i_sdr_pi_cfg_10 = %b", i_sdr_pi_cfg[10]);
   $fdisplay(fd, "i_sdr_pi_cfg_9 = %b", i_sdr_pi_cfg[9]);
   $fdisplay(fd, "i_sdr_pi_cfg_8 = %b", i_sdr_pi_cfg[8]);
   $fdisplay(fd, "i_sdr_pi_cfg_7 = %b", i_sdr_pi_cfg[7]);
   $fdisplay(fd, "i_sdr_pi_cfg_6 = %b", i_sdr_pi_cfg[6]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_33 = %b", i_dq_sdr_rt_pi_cfg[33]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_32 = %b", i_dq_sdr_rt_pi_cfg[32]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_31 = %b", i_dq_sdr_rt_pi_cfg[31]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_30 = %b", i_dq_sdr_rt_pi_cfg[30]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_29 = %b", i_dq_sdr_rt_pi_cfg[29]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_28 = %b", i_dq_sdr_rt_pi_cfg[28]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_27 = %b", i_dq_sdr_rt_pi_cfg[27]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_26 = %b", i_dq_sdr_rt_pi_cfg[26]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_25 = %b", i_dq_sdr_rt_pi_cfg[25]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_24 = %b", i_dq_sdr_rt_pi_cfg[24]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_23 = %b", i_dq_sdr_rt_pi_cfg[23]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_22 = %b", i_dq_sdr_rt_pi_cfg[22]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_21 = %b", i_dq_sdr_rt_pi_cfg[21]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_20 = %b", i_dq_sdr_rt_pi_cfg[20]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_19 = %b", i_dq_sdr_rt_pi_cfg[19]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_18 = %b", i_dq_sdr_rt_pi_cfg[18]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_17 = %b", i_dq_sdr_rt_pi_cfg[17]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_16 = %b", i_dq_sdr_rt_pi_cfg[16]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_14 = %b", i_dq_sdr_rt_pi_cfg[14]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_13 = %b", i_dq_sdr_rt_pi_cfg[13]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_12 = %b", i_dq_sdr_rt_pi_cfg[12]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_11 = %b", i_dq_sdr_rt_pi_cfg[11]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_10 = %b", i_dq_sdr_rt_pi_cfg[10]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_9 = %b", i_dq_sdr_rt_pi_cfg[9]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_8 = %b", i_dq_sdr_rt_pi_cfg[8]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_7 = %b", i_dq_sdr_rt_pi_cfg[7]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_6 = %b", i_dq_sdr_rt_pi_cfg[6]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_33 = %b", i_dq_ddr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_32 = %b", i_dq_ddr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_31 = %b", i_dq_ddr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_30 = %b", i_dq_ddr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_29 = %b", i_dq_ddr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_28 = %b", i_dq_ddr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_27 = %b", i_dq_ddr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_26 = %b", i_dq_ddr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_25 = %b", i_dq_ddr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_24 = %b", i_dq_ddr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_23 = %b", i_dq_ddr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_22 = %b", i_dq_ddr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_21 = %b", i_dq_ddr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_20 = %b", i_dq_ddr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_19 = %b", i_dq_ddr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_18 = %b", i_dq_ddr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_17 = %b", i_dq_ddr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_16 = %b", i_dq_ddr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_14 = %b", i_dq_ddr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_13 = %b", i_dq_ddr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_12 = %b", i_dq_ddr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_11 = %b", i_dq_ddr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_10 = %b", i_dq_ddr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_9 = %b", i_dq_ddr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_8 = %b", i_dq_ddr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_7 = %b", i_dq_ddr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_6 = %b", i_dq_ddr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_33 = %b", i_dq_qdr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_32 = %b", i_dq_qdr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_31 = %b", i_dq_qdr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_30 = %b", i_dq_qdr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_29 = %b", i_dq_qdr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_28 = %b", i_dq_qdr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_27 = %b", i_dq_qdr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_26 = %b", i_dq_qdr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_25 = %b", i_dq_qdr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_24 = %b", i_dq_qdr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_23 = %b", i_dq_qdr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_22 = %b", i_dq_qdr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_21 = %b", i_dq_qdr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_20 = %b", i_dq_qdr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_19 = %b", i_dq_qdr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_18 = %b", i_dq_qdr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_17 = %b", i_dq_qdr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_16 = %b", i_dq_qdr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_14 = %b", i_dq_qdr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_13 = %b", i_dq_qdr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_12 = %b", i_dq_qdr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_11 = %b", i_dq_qdr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_10 = %b", i_dq_qdr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_9 = %b", i_dq_qdr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_8 = %b", i_dq_qdr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_7 = %b", i_dq_qdr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_6 = %b", i_dq_qdr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_80 = %b", i_dq_xdr_lpde_cfg[80]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_79 = %b", i_dq_xdr_lpde_cfg[79]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_78 = %b", i_dq_xdr_lpde_cfg[78]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_77 = %b", i_dq_xdr_lpde_cfg[77]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_76 = %b", i_dq_xdr_lpde_cfg[76]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_75 = %b", i_dq_xdr_lpde_cfg[75]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_74 = %b", i_dq_xdr_lpde_cfg[74]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_73 = %b", i_dq_xdr_lpde_cfg[73]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_72 = %b", i_dq_xdr_lpde_cfg[72]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_71 = %b", i_dq_xdr_lpde_cfg[71]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_70 = %b", i_dq_xdr_lpde_cfg[70]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_69 = %b", i_dq_xdr_lpde_cfg[69]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_68 = %b", i_dq_xdr_lpde_cfg[68]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_67 = %b", i_dq_xdr_lpde_cfg[67]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_66 = %b", i_dq_xdr_lpde_cfg[66]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_65 = %b", i_dq_xdr_lpde_cfg[65]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_64 = %b", i_dq_xdr_lpde_cfg[64]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_63 = %b", i_dq_xdr_lpde_cfg[63]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_62 = %b", i_dq_xdr_lpde_cfg[62]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_61 = %b", i_dq_xdr_lpde_cfg[61]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_60 = %b", i_dq_xdr_lpde_cfg[60]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_59 = %b", i_dq_xdr_lpde_cfg[59]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_58 = %b", i_dq_xdr_lpde_cfg[58]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_57 = %b", i_dq_xdr_lpde_cfg[57]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_56 = %b", i_dq_xdr_lpde_cfg[56]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_55 = %b", i_dq_xdr_lpde_cfg[55]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_54 = %b", i_dq_xdr_lpde_cfg[54]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_53 = %b", i_dq_xdr_lpde_cfg[53]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_52 = %b", i_dq_xdr_lpde_cfg[52]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_51 = %b", i_dq_xdr_lpde_cfg[51]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_50 = %b", i_dq_xdr_lpde_cfg[50]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_49 = %b", i_dq_xdr_lpde_cfg[49]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_48 = %b", i_dq_xdr_lpde_cfg[48]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_47 = %b", i_dq_xdr_lpde_cfg[47]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_46 = %b", i_dq_xdr_lpde_cfg[46]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_45 = %b", i_dq_xdr_lpde_cfg[45]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_44 = %b", i_dq_xdr_lpde_cfg[44]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_43 = %b", i_dq_xdr_lpde_cfg[43]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_42 = %b", i_dq_xdr_lpde_cfg[42]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_41 = %b", i_dq_xdr_lpde_cfg[41]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_40 = %b", i_dq_xdr_lpde_cfg[40]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_39 = %b", i_dq_xdr_lpde_cfg[39]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_38 = %b", i_dq_xdr_lpde_cfg[38]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_37 = %b", i_dq_xdr_lpde_cfg[37]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_36 = %b", i_dq_xdr_lpde_cfg[36]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_35 = %b", i_dq_xdr_lpde_cfg[35]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_34 = %b", i_dq_xdr_lpde_cfg[34]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_33 = %b", i_dq_xdr_lpde_cfg[33]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_32 = %b", i_dq_xdr_lpde_cfg[32]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_31 = %b", i_dq_xdr_lpde_cfg[31]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_30 = %b", i_dq_xdr_lpde_cfg[30]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_29 = %b", i_dq_xdr_lpde_cfg[29]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_28 = %b", i_dq_xdr_lpde_cfg[28]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_27 = %b", i_dq_xdr_lpde_cfg[27]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_26 = %b", i_dq_xdr_lpde_cfg[26]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_25 = %b", i_dq_xdr_lpde_cfg[25]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_24 = %b", i_dq_xdr_lpde_cfg[24]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_23 = %b", i_dq_xdr_lpde_cfg[23]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_22 = %b", i_dq_xdr_lpde_cfg[22]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_21 = %b", i_dq_xdr_lpde_cfg[21]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_20 = %b", i_dq_xdr_lpde_cfg[20]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_19 = %b", i_dq_xdr_lpde_cfg[19]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_18 = %b", i_dq_xdr_lpde_cfg[18]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_17 = %b", i_dq_xdr_lpde_cfg[17]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_16 = %b", i_dq_xdr_lpde_cfg[16]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_15 = %b", i_dq_xdr_lpde_cfg[15]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_14 = %b", i_dq_xdr_lpde_cfg[14]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_13 = %b", i_dq_xdr_lpde_cfg[13]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_12 = %b", i_dq_xdr_lpde_cfg[12]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_11 = %b", i_dq_xdr_lpde_cfg[11]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_10 = %b", i_dq_xdr_lpde_cfg[10]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_9 = %b", i_dq_xdr_lpde_cfg[9]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_8 = %b", i_dq_xdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_7 = %b", i_dq_xdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_6 = %b", i_dq_xdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_5 = %b", i_dq_xdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_4 = %b", i_dq_xdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_3 = %b", i_dq_xdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_2 = %b", i_dq_xdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_1 = %b", i_dq_xdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_0 = %b", i_dq_xdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_8 = %b", i_dq_ddr_1_pipe_en[8]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_7 = %b", i_dq_ddr_1_pipe_en[7]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_6 = %b", i_dq_ddr_1_pipe_en[6]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_5 = %b", i_dq_ddr_1_pipe_en[5]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_4 = %b", i_dq_ddr_1_pipe_en[4]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_3 = %b", i_dq_ddr_1_pipe_en[3]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_2 = %b", i_dq_ddr_1_pipe_en[2]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_1 = %b", i_dq_ddr_1_pipe_en[1]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_0 = %b", i_dq_ddr_1_pipe_en[0]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_16 = %b", i_dq_ddr_1_x_sel[16]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_14 = %b", i_dq_ddr_1_x_sel[14]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_12 = %b", i_dq_ddr_1_x_sel[12]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_10 = %b", i_dq_ddr_1_x_sel[10]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_8 = %b", i_dq_ddr_1_x_sel[8]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_6 = %b", i_dq_ddr_1_x_sel[6]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_4 = %b", i_dq_ddr_1_x_sel[4]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_2 = %b", i_dq_ddr_1_x_sel[2]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_0 = %b", i_dq_ddr_1_x_sel[0]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_8 = %b", i_dq_ddr_0_pipe_en[8]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_7 = %b", i_dq_ddr_0_pipe_en[7]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_6 = %b", i_dq_ddr_0_pipe_en[6]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_5 = %b", i_dq_ddr_0_pipe_en[5]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_4 = %b", i_dq_ddr_0_pipe_en[4]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_3 = %b", i_dq_ddr_0_pipe_en[3]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_2 = %b", i_dq_ddr_0_pipe_en[2]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_1 = %b", i_dq_ddr_0_pipe_en[1]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_0 = %b", i_dq_ddr_0_pipe_en[0]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_16 = %b", i_dq_ddr_0_x_sel[16]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_14 = %b", i_dq_ddr_0_x_sel[14]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_12 = %b", i_dq_ddr_0_x_sel[12]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_10 = %b", i_dq_ddr_0_x_sel[10]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_8 = %b", i_dq_ddr_0_x_sel[8]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_6 = %b", i_dq_ddr_0_x_sel[6]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_4 = %b", i_dq_ddr_0_x_sel[4]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_2 = %b", i_dq_ddr_0_x_sel[2]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_0 = %b", i_dq_ddr_0_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_8 = %b", i_dq_sdr_3_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_7 = %b", i_dq_sdr_3_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_6 = %b", i_dq_sdr_3_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_5 = %b", i_dq_sdr_3_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_4 = %b", i_dq_sdr_3_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_3 = %b", i_dq_sdr_3_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_2 = %b", i_dq_sdr_3_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_1 = %b", i_dq_sdr_3_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_0 = %b", i_dq_sdr_3_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_25 = %b", i_dq_sdr_3_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_24 = %b", i_dq_sdr_3_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_22 = %b", i_dq_sdr_3_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_21 = %b", i_dq_sdr_3_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_19 = %b", i_dq_sdr_3_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_18 = %b", i_dq_sdr_3_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_16 = %b", i_dq_sdr_3_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_15 = %b", i_dq_sdr_3_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_13 = %b", i_dq_sdr_3_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_12 = %b", i_dq_sdr_3_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_10 = %b", i_dq_sdr_3_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_9 = %b", i_dq_sdr_3_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_7 = %b", i_dq_sdr_3_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_6 = %b", i_dq_sdr_3_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_4 = %b", i_dq_sdr_3_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_3 = %b", i_dq_sdr_3_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_1 = %b", i_dq_sdr_3_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_0 = %b", i_dq_sdr_3_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_17 = %b", i_dq_sdr_3_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_16 = %b", i_dq_sdr_3_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_15 = %b", i_dq_sdr_3_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_14 = %b", i_dq_sdr_3_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_13 = %b", i_dq_sdr_3_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_12 = %b", i_dq_sdr_3_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_11 = %b", i_dq_sdr_3_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_10 = %b", i_dq_sdr_3_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_9 = %b", i_dq_sdr_3_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_8 = %b", i_dq_sdr_3_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_7 = %b", i_dq_sdr_3_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_6 = %b", i_dq_sdr_3_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_5 = %b", i_dq_sdr_3_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_4 = %b", i_dq_sdr_3_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_3 = %b", i_dq_sdr_3_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_2 = %b", i_dq_sdr_3_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_1 = %b", i_dq_sdr_3_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_0 = %b", i_dq_sdr_3_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_8 = %b", i_dq_sdr_2_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_7 = %b", i_dq_sdr_2_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_6 = %b", i_dq_sdr_2_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_5 = %b", i_dq_sdr_2_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_4 = %b", i_dq_sdr_2_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_3 = %b", i_dq_sdr_2_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_2 = %b", i_dq_sdr_2_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_1 = %b", i_dq_sdr_2_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_0 = %b", i_dq_sdr_2_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_25 = %b", i_dq_sdr_2_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_24 = %b", i_dq_sdr_2_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_22 = %b", i_dq_sdr_2_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_21 = %b", i_dq_sdr_2_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_19 = %b", i_dq_sdr_2_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_18 = %b", i_dq_sdr_2_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_16 = %b", i_dq_sdr_2_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_15 = %b", i_dq_sdr_2_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_13 = %b", i_dq_sdr_2_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_12 = %b", i_dq_sdr_2_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_10 = %b", i_dq_sdr_2_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_9 = %b", i_dq_sdr_2_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_7 = %b", i_dq_sdr_2_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_6 = %b", i_dq_sdr_2_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_4 = %b", i_dq_sdr_2_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_3 = %b", i_dq_sdr_2_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_1 = %b", i_dq_sdr_2_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_0 = %b", i_dq_sdr_2_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_17 = %b", i_dq_sdr_2_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_16 = %b", i_dq_sdr_2_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_15 = %b", i_dq_sdr_2_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_14 = %b", i_dq_sdr_2_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_13 = %b", i_dq_sdr_2_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_12 = %b", i_dq_sdr_2_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_11 = %b", i_dq_sdr_2_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_10 = %b", i_dq_sdr_2_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_9 = %b", i_dq_sdr_2_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_8 = %b", i_dq_sdr_2_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_7 = %b", i_dq_sdr_2_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_6 = %b", i_dq_sdr_2_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_5 = %b", i_dq_sdr_2_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_4 = %b", i_dq_sdr_2_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_3 = %b", i_dq_sdr_2_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_2 = %b", i_dq_sdr_2_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_1 = %b", i_dq_sdr_2_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_0 = %b", i_dq_sdr_2_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_8 = %b", i_dq_sdr_1_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_7 = %b", i_dq_sdr_1_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_6 = %b", i_dq_sdr_1_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_5 = %b", i_dq_sdr_1_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_4 = %b", i_dq_sdr_1_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_3 = %b", i_dq_sdr_1_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_2 = %b", i_dq_sdr_1_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_1 = %b", i_dq_sdr_1_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_0 = %b", i_dq_sdr_1_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_25 = %b", i_dq_sdr_1_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_24 = %b", i_dq_sdr_1_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_22 = %b", i_dq_sdr_1_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_21 = %b", i_dq_sdr_1_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_19 = %b", i_dq_sdr_1_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_18 = %b", i_dq_sdr_1_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_16 = %b", i_dq_sdr_1_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_15 = %b", i_dq_sdr_1_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_13 = %b", i_dq_sdr_1_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_12 = %b", i_dq_sdr_1_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_10 = %b", i_dq_sdr_1_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_9 = %b", i_dq_sdr_1_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_7 = %b", i_dq_sdr_1_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_6 = %b", i_dq_sdr_1_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_4 = %b", i_dq_sdr_1_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_3 = %b", i_dq_sdr_1_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_1 = %b", i_dq_sdr_1_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_0 = %b", i_dq_sdr_1_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_17 = %b", i_dq_sdr_1_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_16 = %b", i_dq_sdr_1_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_15 = %b", i_dq_sdr_1_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_14 = %b", i_dq_sdr_1_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_13 = %b", i_dq_sdr_1_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_12 = %b", i_dq_sdr_1_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_11 = %b", i_dq_sdr_1_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_10 = %b", i_dq_sdr_1_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_9 = %b", i_dq_sdr_1_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_8 = %b", i_dq_sdr_1_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_7 = %b", i_dq_sdr_1_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_6 = %b", i_dq_sdr_1_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_5 = %b", i_dq_sdr_1_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_4 = %b", i_dq_sdr_1_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_3 = %b", i_dq_sdr_1_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_2 = %b", i_dq_sdr_1_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_1 = %b", i_dq_sdr_1_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_0 = %b", i_dq_sdr_1_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_8 = %b", i_dq_sdr_0_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_7 = %b", i_dq_sdr_0_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_6 = %b", i_dq_sdr_0_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_5 = %b", i_dq_sdr_0_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_4 = %b", i_dq_sdr_0_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_3 = %b", i_dq_sdr_0_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_2 = %b", i_dq_sdr_0_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_1 = %b", i_dq_sdr_0_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_0 = %b", i_dq_sdr_0_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_25 = %b", i_dq_sdr_0_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_24 = %b", i_dq_sdr_0_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_22 = %b", i_dq_sdr_0_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_21 = %b", i_dq_sdr_0_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_19 = %b", i_dq_sdr_0_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_18 = %b", i_dq_sdr_0_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_16 = %b", i_dq_sdr_0_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_15 = %b", i_dq_sdr_0_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_13 = %b", i_dq_sdr_0_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_12 = %b", i_dq_sdr_0_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_10 = %b", i_dq_sdr_0_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_9 = %b", i_dq_sdr_0_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_7 = %b", i_dq_sdr_0_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_6 = %b", i_dq_sdr_0_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_4 = %b", i_dq_sdr_0_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_3 = %b", i_dq_sdr_0_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_1 = %b", i_dq_sdr_0_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_0 = %b", i_dq_sdr_0_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_17 = %b", i_dq_sdr_0_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_16 = %b", i_dq_sdr_0_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_15 = %b", i_dq_sdr_0_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_14 = %b", i_dq_sdr_0_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_13 = %b", i_dq_sdr_0_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_12 = %b", i_dq_sdr_0_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_11 = %b", i_dq_sdr_0_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_10 = %b", i_dq_sdr_0_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_9 = %b", i_dq_sdr_0_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_8 = %b", i_dq_sdr_0_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_7 = %b", i_dq_sdr_0_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_6 = %b", i_dq_sdr_0_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_5 = %b", i_dq_sdr_0_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_4 = %b", i_dq_sdr_0_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_3 = %b", i_dq_sdr_0_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_2 = %b", i_dq_sdr_0_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_1 = %b", i_dq_sdr_0_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_0 = %b", i_dq_sdr_0_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_8 = %b", i_dq_sdr_rt_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_7 = %b", i_dq_sdr_rt_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_6 = %b", i_dq_sdr_rt_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_5 = %b", i_dq_sdr_rt_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_4 = %b", i_dq_sdr_rt_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_3 = %b", i_dq_sdr_rt_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_2 = %b", i_dq_sdr_rt_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_1 = %b", i_dq_sdr_rt_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_0 = %b", i_dq_sdr_rt_pipe_en[0]);
   $fdisplay(fd, "i_dq_egress_mode_dig_62 = %b", i_dq_egress_mode_dig[62]);
   $fdisplay(fd, "i_dq_egress_mode_dig_57 = %b", i_dq_egress_mode_dig[57]);
   $fdisplay(fd, "i_dq_egress_mode_dig_56 = %b", i_dq_egress_mode_dig[56]);
   $fdisplay(fd, "i_dq_egress_mode_dig_55 = %b", i_dq_egress_mode_dig[55]);
   $fdisplay(fd, "i_dq_egress_mode_dig_50 = %b", i_dq_egress_mode_dig[50]);
   $fdisplay(fd, "i_dq_egress_mode_dig_49 = %b", i_dq_egress_mode_dig[49]);
   $fdisplay(fd, "i_dq_egress_mode_dig_48 = %b", i_dq_egress_mode_dig[48]);
   $fdisplay(fd, "i_dq_egress_mode_dig_43 = %b", i_dq_egress_mode_dig[43]);
   $fdisplay(fd, "i_dq_egress_mode_dig_42 = %b", i_dq_egress_mode_dig[42]);
   $fdisplay(fd, "i_dq_egress_mode_dig_41 = %b", i_dq_egress_mode_dig[41]);
   $fdisplay(fd, "i_dq_egress_mode_dig_36 = %b", i_dq_egress_mode_dig[36]);
   $fdisplay(fd, "i_dq_egress_mode_dig_35 = %b", i_dq_egress_mode_dig[35]);
   $fdisplay(fd, "i_dq_egress_mode_dig_34 = %b", i_dq_egress_mode_dig[34]);
   $fdisplay(fd, "i_dq_egress_mode_dig_29 = %b", i_dq_egress_mode_dig[29]);
   $fdisplay(fd, "i_dq_egress_mode_dig_28 = %b", i_dq_egress_mode_dig[28]);
   $fdisplay(fd, "i_dq_egress_mode_dig_27 = %b", i_dq_egress_mode_dig[27]);
   $fdisplay(fd, "i_dq_egress_mode_dig_22 = %b", i_dq_egress_mode_dig[22]);
   $fdisplay(fd, "i_dq_egress_mode_dig_21 = %b", i_dq_egress_mode_dig[21]);
   $fdisplay(fd, "i_dq_egress_mode_dig_20 = %b", i_dq_egress_mode_dig[20]);
   $fdisplay(fd, "i_dq_egress_mode_dig_15 = %b", i_dq_egress_mode_dig[15]);
   $fdisplay(fd, "i_dq_egress_mode_dig_14 = %b", i_dq_egress_mode_dig[14]);
   $fdisplay(fd, "i_dq_egress_mode_dig_13 = %b", i_dq_egress_mode_dig[13]);
   $fdisplay(fd, "i_dq_egress_mode_dig_8 = %b", i_dq_egress_mode_dig[8]);
   $fdisplay(fd, "i_dq_egress_mode_dig_7 = %b", i_dq_egress_mode_dig[7]);
   $fdisplay(fd, "i_dq_egress_mode_dig_6 = %b", i_dq_egress_mode_dig[6]);
   $fdisplay(fd, "i_dq_egress_mode_dig_1 = %b", i_dq_egress_mode_dig[1]);
   $fdisplay(fd, "i_dq_egress_mode_dig_0 = %b", i_dq_egress_mode_dig[0]);
   $fdisplay(fd, "i_dq_egress_mode_ana_50 = %b", i_dq_egress_mode_ana[50]);
   $fdisplay(fd, "i_dq_egress_mode_ana_49 = %b", i_dq_egress_mode_ana[49]);
   $fdisplay(fd, "i_dq_egress_mode_ana_48 = %b", i_dq_egress_mode_ana[48]);
   $fdisplay(fd, "i_dq_egress_mode_ana_44 = %b", i_dq_egress_mode_ana[44]);
   $fdisplay(fd, "i_dq_egress_mode_ana_43 = %b", i_dq_egress_mode_ana[43]);
   $fdisplay(fd, "i_dq_egress_mode_ana_42 = %b", i_dq_egress_mode_ana[42]);
   $fdisplay(fd, "i_dq_egress_mode_ana_38 = %b", i_dq_egress_mode_ana[38]);
   $fdisplay(fd, "i_dq_egress_mode_ana_37 = %b", i_dq_egress_mode_ana[37]);
   $fdisplay(fd, "i_dq_egress_mode_ana_36 = %b", i_dq_egress_mode_ana[36]);
   $fdisplay(fd, "i_dq_egress_mode_ana_32 = %b", i_dq_egress_mode_ana[32]);
   $fdisplay(fd, "i_dq_egress_mode_ana_31 = %b", i_dq_egress_mode_ana[31]);
   $fdisplay(fd, "i_dq_egress_mode_ana_30 = %b", i_dq_egress_mode_ana[30]);
   $fdisplay(fd, "i_dq_egress_mode_ana_26 = %b", i_dq_egress_mode_ana[26]);
   $fdisplay(fd, "i_dq_egress_mode_ana_25 = %b", i_dq_egress_mode_ana[25]);
   $fdisplay(fd, "i_dq_egress_mode_ana_24 = %b", i_dq_egress_mode_ana[24]);
   $fdisplay(fd, "i_dq_egress_mode_ana_20 = %b", i_dq_egress_mode_ana[20]);
   $fdisplay(fd, "i_dq_egress_mode_ana_19 = %b", i_dq_egress_mode_ana[19]);
   $fdisplay(fd, "i_dq_egress_mode_ana_18 = %b", i_dq_egress_mode_ana[18]);
   $fdisplay(fd, "i_dq_egress_mode_ana_14 = %b", i_dq_egress_mode_ana[14]);
   $fdisplay(fd, "i_dq_egress_mode_ana_13 = %b", i_dq_egress_mode_ana[13]);
   $fdisplay(fd, "i_dq_egress_mode_ana_12 = %b", i_dq_egress_mode_ana[12]);
   $fdisplay(fd, "i_dq_egress_mode_ana_8 = %b", i_dq_egress_mode_ana[8]);
   $fdisplay(fd, "i_dq_egress_mode_ana_7 = %b", i_dq_egress_mode_ana[7]);
   $fdisplay(fd, "i_dq_egress_mode_ana_6 = %b", i_dq_egress_mode_ana[6]);
   $fdisplay(fd, "i_dq_egress_mode_ana_2 = %b", i_dq_egress_mode_ana[2]);
   $fdisplay(fd, "i_dq_egress_mode_ana_1 = %b", i_dq_egress_mode_ana[1]);
   $fdisplay(fd, "i_dq_egress_mode_ana_0 = %b", i_dq_egress_mode_ana[0]);
   $fdisplay(fd, "i_pll_clk_270 = %b", i_pll_clk_270);
   $fdisplay(fd, "i_pll_clk_180 = %b", i_pll_clk_180);
   $fdisplay(fd, "i_pll_clk_90 = %b", i_pll_clk_90);
   $fdisplay(fd, "i_pll_clk_0 = %b", i_pll_clk_0);
   $fdisplay(fd, "i_rst = %b", i_rst);
   $fdisplay(fd, "i_scan_mode = %b", i_scan_mode);
   $fdisplay(fd, "i_scan_clk = %b", i_scan_clk);

endtask

task oprint_ddr_dq (input integer fd);

   $fdisplay(fd, "INFO: Edge Trigger [%t] ...", $realtime);

   $fdisplay(fd, "o_dqs_pad_bscan_c_1 = %b", o_dqs_pad_bscan_c[1]);
   $fdisplay(fd, "o_dqs_pad_bscan_c_0 = %b", o_dqs_pad_bscan_c[0]);
   $fdisplay(fd, "o_dqs_pad_bscan_t_1 = %b", o_dqs_pad_bscan_t[1]);
   $fdisplay(fd, "o_dqs_pad_bscan_t_0 = %b", o_dqs_pad_bscan_t[0]);
   $fdisplay(fd, "o_dq_pad_bscan_t_8 = %b", o_dq_pad_bscan_t[8]);
   $fdisplay(fd, "o_dq_pad_bscan_t_7 = %b", o_dq_pad_bscan_t[7]);
   $fdisplay(fd, "o_dq_pad_bscan_t_6 = %b", o_dq_pad_bscan_t[6]);
   $fdisplay(fd, "o_dq_pad_bscan_t_5 = %b", o_dq_pad_bscan_t[5]);
   $fdisplay(fd, "o_dq_pad_bscan_t_4 = %b", o_dq_pad_bscan_t[4]);
   $fdisplay(fd, "o_dq_pad_bscan_t_3 = %b", o_dq_pad_bscan_t[3]);
   $fdisplay(fd, "o_dq_pad_bscan_t_2 = %b", o_dq_pad_bscan_t[2]);
   $fdisplay(fd, "o_dq_pad_bscan_t_1 = %b", o_dq_pad_bscan_t[1]);
   $fdisplay(fd, "o_dq_pad_bscan_t_0 = %b", o_dq_pad_bscan_t[0]);
   $fdisplay(fd, "o_dq_core_eg_8 = %b", o_dq_core_eg[8]);
   $fdisplay(fd, "o_dq_core_eg_7 = %b", o_dq_core_eg[7]);
   $fdisplay(fd, "o_dq_core_eg_6 = %b", o_dq_core_eg[6]);
   $fdisplay(fd, "o_dq_core_eg_5 = %b", o_dq_core_eg[5]);
   $fdisplay(fd, "o_dq_core_eg_4 = %b", o_dq_core_eg[4]);
   $fdisplay(fd, "o_dq_core_eg_3 = %b", o_dq_core_eg[3]);
   $fdisplay(fd, "o_dq_core_eg_2 = %b", o_dq_core_eg[2]);
   $fdisplay(fd, "o_dq_core_eg_1 = %b", o_dq_core_eg[1]);
   $fdisplay(fd, "o_dq_core_eg_0 = %b", o_dq_core_eg[0]);
   $fdisplay(fd, "o_dq_core_ig_8 = %b", o_dq_core_ig[8]);
   $fdisplay(fd, "o_dq_core_ig_7 = %b", o_dq_core_ig[7]);
   $fdisplay(fd, "o_dq_core_ig_6 = %b", o_dq_core_ig[6]);
   $fdisplay(fd, "o_dq_core_ig_5 = %b", o_dq_core_ig[5]);
   $fdisplay(fd, "o_dq_core_ig_4 = %b", o_dq_core_ig[4]);
   $fdisplay(fd, "o_dq_core_ig_3 = %b", o_dq_core_ig[3]);
   $fdisplay(fd, "o_dq_core_ig_2 = %b", o_dq_core_ig[2]);
   $fdisplay(fd, "o_dq_core_ig_1 = %b", o_dq_core_ig[1]);
   $fdisplay(fd, "o_dq_core_ig_0 = %b", o_dq_core_ig[0]);
   $fdisplay(fd, "o_dqs_core_eg_8 = %b", o_dqs_core_eg[8]);
   $fdisplay(fd, "o_dqs_core_eg_7 = %b", o_dqs_core_eg[7]);
   $fdisplay(fd, "o_dqs_core_eg_6 = %b", o_dqs_core_eg[6]);
   $fdisplay(fd, "o_dqs_core_eg_5 = %b", o_dqs_core_eg[5]);
   $fdisplay(fd, "o_dqs_core_eg_4 = %b", o_dqs_core_eg[4]);
   $fdisplay(fd, "o_dqs_core_eg_3 = %b", o_dqs_core_eg[3]);
   $fdisplay(fd, "o_dqs_core_eg_2 = %b", o_dqs_core_eg[2]);
   $fdisplay(fd, "o_dqs_core_eg_1 = %b", o_dqs_core_eg[1]);
   $fdisplay(fd, "o_dqs_core_eg_0 = %b", o_dqs_core_eg[0]);
   $fdisplay(fd, "o_dqs_core_ig_8 = %b", o_dqs_core_ig[8]);
   $fdisplay(fd, "o_dqs_core_ig_7 = %b", o_dqs_core_ig[7]);
   $fdisplay(fd, "o_dqs_core_ig_6 = %b", o_dqs_core_ig[6]);
   $fdisplay(fd, "o_dqs_core_ig_5 = %b", o_dqs_core_ig[5]);
   $fdisplay(fd, "o_dqs_core_ig_4 = %b", o_dqs_core_ig[4]);
   $fdisplay(fd, "o_dqs_core_ig_3 = %b", o_dqs_core_ig[3]);
   $fdisplay(fd, "o_dqs_core_ig_2 = %b", o_dqs_core_ig[2]);
   $fdisplay(fd, "o_dqs_core_ig_1 = %b", o_dqs_core_ig[1]);
   $fdisplay(fd, "o_dqs_core_ig_0 = %b", o_dqs_core_ig[0]);
   $fdisplay(fd, "o_dqs_ren_pi_phase_sta = %b", o_dqs_ren_pi_phase_sta);
   $fdisplay(fd, "o_dqs_rcs_pi_phase_sta = %b", o_dqs_rcs_pi_phase_sta);
   $fdisplay(fd, "o_dq_sdr_35 = %b", o_dq_sdr[35]);
   $fdisplay(fd, "o_dq_sdr_34 = %b", o_dq_sdr[34]);
   $fdisplay(fd, "o_dq_sdr_33 = %b", o_dq_sdr[33]);
   $fdisplay(fd, "o_dq_sdr_32 = %b", o_dq_sdr[32]);
   $fdisplay(fd, "o_dq_sdr_31 = %b", o_dq_sdr[31]);
   $fdisplay(fd, "o_dq_sdr_30 = %b", o_dq_sdr[30]);
   $fdisplay(fd, "o_dq_sdr_29 = %b", o_dq_sdr[29]);
   $fdisplay(fd, "o_dq_sdr_28 = %b", o_dq_sdr[28]);
   $fdisplay(fd, "o_dq_sdr_27 = %b", o_dq_sdr[27]);
   $fdisplay(fd, "o_dq_sdr_26 = %b", o_dq_sdr[26]);
   $fdisplay(fd, "o_dq_sdr_25 = %b", o_dq_sdr[25]);
   $fdisplay(fd, "o_dq_sdr_24 = %b", o_dq_sdr[24]);
   $fdisplay(fd, "o_dq_sdr_23 = %b", o_dq_sdr[23]);
   $fdisplay(fd, "o_dq_sdr_22 = %b", o_dq_sdr[22]);
   $fdisplay(fd, "o_dq_sdr_21 = %b", o_dq_sdr[21]);
   $fdisplay(fd, "o_dq_sdr_20 = %b", o_dq_sdr[20]);
   $fdisplay(fd, "o_dq_sdr_19 = %b", o_dq_sdr[19]);
   $fdisplay(fd, "o_dq_sdr_18 = %b", o_dq_sdr[18]);
   $fdisplay(fd, "o_dq_sdr_17 = %b", o_dq_sdr[17]);
   $fdisplay(fd, "o_dq_sdr_16 = %b", o_dq_sdr[16]);
   $fdisplay(fd, "o_dq_sdr_15 = %b", o_dq_sdr[15]);
   $fdisplay(fd, "o_dq_sdr_14 = %b", o_dq_sdr[14]);
   $fdisplay(fd, "o_dq_sdr_13 = %b", o_dq_sdr[13]);
   $fdisplay(fd, "o_dq_sdr_12 = %b", o_dq_sdr[12]);
   $fdisplay(fd, "o_dq_sdr_11 = %b", o_dq_sdr[11]);
   $fdisplay(fd, "o_dq_sdr_10 = %b", o_dq_sdr[10]);
   $fdisplay(fd, "o_dq_sdr_9 = %b", o_dq_sdr[9]);
   $fdisplay(fd, "o_dq_sdr_8 = %b", o_dq_sdr[8]);
   $fdisplay(fd, "o_dq_sdr_7 = %b", o_dq_sdr[7]);
   $fdisplay(fd, "o_dq_sdr_6 = %b", o_dq_sdr[6]);
   $fdisplay(fd, "o_dq_sdr_5 = %b", o_dq_sdr[5]);
   $fdisplay(fd, "o_dq_sdr_4 = %b", o_dq_sdr[4]);
   $fdisplay(fd, "o_dq_sdr_3 = %b", o_dq_sdr[3]);
   $fdisplay(fd, "o_dq_sdr_2 = %b", o_dq_sdr[2]);
   $fdisplay(fd, "o_dq_sdr_1 = %b", o_dq_sdr[1]);
   $fdisplay(fd, "o_dq_sdr_0 = %b", o_dq_sdr[0]);
   $fdisplay(fd, "o_dq_sa_35 = %b", o_dq_sa[35]);
   $fdisplay(fd, "o_dq_sa_34 = %b", o_dq_sa[34]);
   $fdisplay(fd, "o_dq_sa_33 = %b", o_dq_sa[33]);
   $fdisplay(fd, "o_dq_sa_32 = %b", o_dq_sa[32]);
   $fdisplay(fd, "o_dq_sa_31 = %b", o_dq_sa[31]);
   $fdisplay(fd, "o_dq_sa_30 = %b", o_dq_sa[30]);
   $fdisplay(fd, "o_dq_sa_29 = %b", o_dq_sa[29]);
   $fdisplay(fd, "o_dq_sa_28 = %b", o_dq_sa[28]);
   $fdisplay(fd, "o_dq_sa_27 = %b", o_dq_sa[27]);
   $fdisplay(fd, "o_dq_sa_26 = %b", o_dq_sa[26]);
   $fdisplay(fd, "o_dq_sa_25 = %b", o_dq_sa[25]);
   $fdisplay(fd, "o_dq_sa_24 = %b", o_dq_sa[24]);
   $fdisplay(fd, "o_dq_sa_23 = %b", o_dq_sa[23]);
   $fdisplay(fd, "o_dq_sa_22 = %b", o_dq_sa[22]);
   $fdisplay(fd, "o_dq_sa_21 = %b", o_dq_sa[21]);
   $fdisplay(fd, "o_dq_sa_20 = %b", o_dq_sa[20]);
   $fdisplay(fd, "o_dq_sa_19 = %b", o_dq_sa[19]);
   $fdisplay(fd, "o_dq_sa_18 = %b", o_dq_sa[18]);
   $fdisplay(fd, "o_dq_sa_17 = %b", o_dq_sa[17]);
   $fdisplay(fd, "o_dq_sa_16 = %b", o_dq_sa[16]);
   $fdisplay(fd, "o_dq_sa_15 = %b", o_dq_sa[15]);
   $fdisplay(fd, "o_dq_sa_14 = %b", o_dq_sa[14]);
   $fdisplay(fd, "o_dq_sa_13 = %b", o_dq_sa[13]);
   $fdisplay(fd, "o_dq_sa_12 = %b", o_dq_sa[12]);
   $fdisplay(fd, "o_dq_sa_11 = %b", o_dq_sa[11]);
   $fdisplay(fd, "o_dq_sa_10 = %b", o_dq_sa[10]);
   $fdisplay(fd, "o_dq_sa_9 = %b", o_dq_sa[9]);
   $fdisplay(fd, "o_dq_sa_8 = %b", o_dq_sa[8]);
   $fdisplay(fd, "o_dq_sa_7 = %b", o_dq_sa[7]);
   $fdisplay(fd, "o_dq_sa_6 = %b", o_dq_sa[6]);
   $fdisplay(fd, "o_dq_sa_5 = %b", o_dq_sa[5]);
   $fdisplay(fd, "o_dq_sa_4 = %b", o_dq_sa[4]);
   $fdisplay(fd, "o_dq_sa_3 = %b", o_dq_sa[3]);
   $fdisplay(fd, "o_dq_sa_2 = %b", o_dq_sa[2]);
   $fdisplay(fd, "o_dq_sa_1 = %b", o_dq_sa[1]);
   $fdisplay(fd, "o_dq_sa_0 = %b", o_dq_sa[0]);
   $fdisplay(fd, "o_rcs = %b", o_rcs);
   $fdisplay(fd, "o_dfird_clk_2 = %b", o_dfird_clk_2);
   $fdisplay(fd, "o_dfird_clk_1 = %b", o_dfird_clk_1);
   $fdisplay(fd, "o_dfiwr_clk_2 = %b", o_dfiwr_clk_2);
   $fdisplay(fd, "o_dfiwr_clk_1 = %b", o_dfiwr_clk_1);
   $fdisplay(fd, "o_rx_sdr__clk = %b", o_rx_sdr_clk);
   $fdisplay(fd, "o_phy_clk = %b", o_phy_clk);
   $fdisplay(fd, "o_tst_clk_1 = %b", o_tst_clk[1]);
   $fdisplay(fd, "o_tst_clk_0 = %b", o_tst_clk[0]);

endtask

task iprint_ddr_ca (input integer fd);

   $fdisplay(fd, "INFO: Edge Trigger [%t] ...", $realtime);
   $fdisplay(fd, "i_dqs_pad_bscan_c_0 = %b", i_dqs_pad_bscan_c[0]);
   $fdisplay(fd, "i_dqs_pad_bscan_t_0 = %b", i_dqs_pad_bscan_t[0]);
   $fdisplay(fd, "i_dqs_pad_bscan_ie = %b", i_dqs_pad_bscan_ie);
   $fdisplay(fd, "i_dqs_pad_bscan_oe = %b", i_dqs_pad_bscan_oe);
   $fdisplay(fd, "i_dqs_pad_bscan_n = %b", i_dqs_pad_bscan_n);
   $fdisplay(fd, "i_dq_pad_bscan_t_10 = %b", i_dq_pad_bscan_t[10]);
   $fdisplay(fd, "i_dq_pad_bscan_t_9 = %b", i_dq_pad_bscan_t[9]);
   $fdisplay(fd, "i_dq_pad_bscan_t_8 = %b", i_dq_pad_bscan_t[8]);
   $fdisplay(fd, "i_dq_pad_bscan_t_7 = %b", i_dq_pad_bscan_t[7]);
   $fdisplay(fd, "i_dq_pad_bscan_t_6 = %b", i_dq_pad_bscan_t[6]);
   $fdisplay(fd, "i_dq_pad_bscan_t_5 = %b", i_dq_pad_bscan_t[5]);
   $fdisplay(fd, "i_dq_pad_bscan_t_4 = %b", i_dq_pad_bscan_t[4]);
   $fdisplay(fd, "i_dq_pad_bscan_t_3 = %b", i_dq_pad_bscan_t[3]);
   $fdisplay(fd, "i_dq_pad_bscan_t_2 = %b", i_dq_pad_bscan_t[2]);
   $fdisplay(fd, "i_dq_pad_bscan_t_1 = %b", i_dq_pad_bscan_t[1]);
   $fdisplay(fd, "i_dq_pad_bscan_t_0 = %b", i_dq_pad_bscan_t[0]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_125 = %b", i_dq_pad_tx_cfg[125]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_123 = %b", i_dq_pad_tx_cfg[123]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_122 = %b", i_dq_pad_tx_cfg[122]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_121 = %b", i_dq_pad_tx_cfg[121]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_120 = %b", i_dq_pad_tx_cfg[120]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_113 = %b", i_dq_pad_tx_cfg[113]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_111 = %b", i_dq_pad_tx_cfg[111]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_110 = %b", i_dq_pad_tx_cfg[110]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_109 = %b", i_dq_pad_tx_cfg[109]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_108 = %b", i_dq_pad_tx_cfg[108]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_107 = %b", i_dq_pad_tx_cfg[107]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_106 = %b", i_dq_pad_tx_cfg[106]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_105 = %b", i_dq_pad_tx_cfg[105]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_104 = %b", i_dq_pad_tx_cfg[104]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_103 = %b", i_dq_pad_tx_cfg[103]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_102 = %b", i_dq_pad_tx_cfg[102]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_101 = %b", i_dq_pad_tx_cfg[101]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_99 = %b", i_dq_pad_tx_cfg[99]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_98 = %b", i_dq_pad_tx_cfg[98]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_97 = %b", i_dq_pad_tx_cfg[97]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_96 = %b", i_dq_pad_tx_cfg[96]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_95 = %b", i_dq_pad_tx_cfg[95]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_94 = %b", i_dq_pad_tx_cfg[94]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_93 = %b", i_dq_pad_tx_cfg[93]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_92 = %b", i_dq_pad_tx_cfg[92]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_91 = %b", i_dq_pad_tx_cfg[91]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_90 = %b", i_dq_pad_tx_cfg[90]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_89 = %b", i_dq_pad_tx_cfg[89]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_87 = %b", i_dq_pad_tx_cfg[87]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_86 = %b", i_dq_pad_tx_cfg[86]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_85 = %b", i_dq_pad_tx_cfg[85]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_84 = %b", i_dq_pad_tx_cfg[84]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_83 = %b", i_dq_pad_tx_cfg[83]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_82 = %b", i_dq_pad_tx_cfg[82]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_81 = %b", i_dq_pad_tx_cfg[81]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_80 = %b", i_dq_pad_tx_cfg[80]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_79 = %b", i_dq_pad_tx_cfg[79]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_78 = %b", i_dq_pad_tx_cfg[78]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_77 = %b", i_dq_pad_tx_cfg[77]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_75 = %b", i_dq_pad_tx_cfg[75]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_74 = %b", i_dq_pad_tx_cfg[74]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_73 = %b", i_dq_pad_tx_cfg[73]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_72 = %b", i_dq_pad_tx_cfg[72]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_71 = %b", i_dq_pad_tx_cfg[71]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_70 = %b", i_dq_pad_tx_cfg[70]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_69 = %b", i_dq_pad_tx_cfg[69]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_68 = %b", i_dq_pad_tx_cfg[68]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_67 = %b", i_dq_pad_tx_cfg[67]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_66 = %b", i_dq_pad_tx_cfg[66]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_65 = %b", i_dq_pad_tx_cfg[65]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_63 = %b", i_dq_pad_tx_cfg[63]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_62 = %b", i_dq_pad_tx_cfg[62]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_61 = %b", i_dq_pad_tx_cfg[61]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_60 = %b", i_dq_pad_tx_cfg[60]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_59 = %b", i_dq_pad_tx_cfg[59]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_58 = %b", i_dq_pad_tx_cfg[58]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_57 = %b", i_dq_pad_tx_cfg[57]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_56 = %b", i_dq_pad_tx_cfg[56]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_55 = %b", i_dq_pad_tx_cfg[55]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_54 = %b", i_dq_pad_tx_cfg[54]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_53 = %b", i_dq_pad_tx_cfg[53]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_51 = %b", i_dq_pad_tx_cfg[51]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_50 = %b", i_dq_pad_tx_cfg[50]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_49 = %b", i_dq_pad_tx_cfg[49]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_48 = %b", i_dq_pad_tx_cfg[48]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_47 = %b", i_dq_pad_tx_cfg[47]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_46 = %b", i_dq_pad_tx_cfg[46]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_45 = %b", i_dq_pad_tx_cfg[45]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_44 = %b", i_dq_pad_tx_cfg[44]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_43 = %b", i_dq_pad_tx_cfg[43]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_42 = %b", i_dq_pad_tx_cfg[42]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_41 = %b", i_dq_pad_tx_cfg[41]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_39 = %b", i_dq_pad_tx_cfg[39]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_38 = %b", i_dq_pad_tx_cfg[38]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_37 = %b", i_dq_pad_tx_cfg[37]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_36 = %b", i_dq_pad_tx_cfg[36]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_35 = %b", i_dq_pad_tx_cfg[35]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_34 = %b", i_dq_pad_tx_cfg[34]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_33 = %b", i_dq_pad_tx_cfg[33]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_32 = %b", i_dq_pad_tx_cfg[32]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_31 = %b", i_dq_pad_tx_cfg[31]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_30 = %b", i_dq_pad_tx_cfg[30]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_29 = %b", i_dq_pad_tx_cfg[29]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_27 = %b", i_dq_pad_tx_cfg[27]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_26 = %b", i_dq_pad_tx_cfg[26]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_25 = %b", i_dq_pad_tx_cfg[25]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_24 = %b", i_dq_pad_tx_cfg[24]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_23 = %b", i_dq_pad_tx_cfg[23]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_22 = %b", i_dq_pad_tx_cfg[22]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_21 = %b", i_dq_pad_tx_cfg[21]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_20 = %b", i_dq_pad_tx_cfg[20]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_19 = %b", i_dq_pad_tx_cfg[19]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_18 = %b", i_dq_pad_tx_cfg[18]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_17 = %b", i_dq_pad_tx_cfg[17]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_15 = %b", i_dq_pad_tx_cfg[15]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_14 = %b", i_dq_pad_tx_cfg[14]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_13 = %b", i_dq_pad_tx_cfg[13]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_12 = %b", i_dq_pad_tx_cfg[12]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_11 = %b", i_dq_pad_tx_cfg[11]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_10 = %b", i_dq_pad_tx_cfg[10]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_9 = %b", i_dq_pad_tx_cfg[9]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_8 = %b", i_dq_pad_tx_cfg[8]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_7 = %b", i_dq_pad_tx_cfg[7]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_6 = %b", i_dq_pad_tx_cfg[6]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_5 = %b", i_dq_pad_tx_cfg[5]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_3 = %b", i_dq_pad_tx_cfg[3]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_2 = %b", i_dq_pad_tx_cfg[2]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_1 = %b", i_dq_pad_tx_cfg[1]);
   $fdisplay(fd, "i_dq_pad_tx_cfg_0 = %b", i_dq_pad_tx_cfg[0]);
   $fdisplay(fd, "i_dq_freeze_n_hv = %b", i_dq_freeze_n_hv);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_13 = %b", i_dqs_pad_tx_cmn_cfg[13]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_12 = %b", i_dqs_pad_tx_cmn_cfg[12]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_11 = %b", i_dqs_pad_tx_cmn_cfg[11]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_10 = %b", i_dqs_pad_tx_cmn_cfg[10]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_9 = %b", i_dqs_pad_tx_cmn_cfg[9]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_8 = %b", i_dqs_pad_tx_cmn_cfg[8]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_7 = %b", i_dqs_pad_tx_cmn_cfg[7]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_6 = %b", i_dqs_pad_tx_cmn_cfg[6]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_5 = %b", i_dqs_pad_tx_cmn_cfg[5]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_4 = %b", i_dqs_pad_tx_cmn_cfg[4]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_3 = %b", i_dqs_pad_tx_cmn_cfg[3]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_2 = %b", i_dqs_pad_tx_cmn_cfg[2]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_1 = %b", i_dqs_pad_tx_cmn_cfg[1]);
   $fdisplay(fd, "i_dqs_pad_tx_cmn_cfg_0 = %b", i_dqs_pad_tx_cmn_cfg[0]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_11 = %b", i_dqs_pad_tx_cfg[11]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_10 = %b", i_dqs_pad_tx_cfg[10]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_9 = %b", i_dqs_pad_tx_cfg[9]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_8 = %b", i_dqs_pad_tx_cfg[8]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_7 = %b", i_dqs_pad_tx_cfg[7]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_6 = %b", i_dqs_pad_tx_cfg[6]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_5 = %b", i_dqs_pad_tx_cfg[5]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_4 = %b", i_dqs_pad_tx_cfg[4]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_3 = %b", i_dqs_pad_tx_cfg[3]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_2 = %b", i_dqs_pad_tx_cfg[2]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_1 = %b", i_dqs_pad_tx_cfg[1]);
   $fdisplay(fd, "i_dqs_pad_tx_cfg_0 = %b", i_dqs_pad_tx_cfg[0]);
   $fdisplay(fd, "i_dqs_hiz_n = %b", i_dqs_hiz_n);
   $fdisplay(fd, "i_dq_cmn_freeze_n = %b", i_dq_cmn_freeze_n);
   $fdisplay(fd, "i_dqs_pre_filter_sel_1 = %b", i_dqs_pre_filter_sel[1]);
   $fdisplay(fd, "i_dqs_pre_filter_sel_0 = %b", i_dqs_pre_filter_sel[0]);
   $fdisplay(fd, "i_dqs_wck_mode = %b", i_dqs_wck_mode);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_8 = %b", i_dqs_sdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_7 = %b", i_dqs_sdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_6 = %b", i_dqs_sdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_5 = %b", i_dqs_sdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_4 = %b", i_dqs_sdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_3 = %b", i_dqs_sdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_2 = %b", i_dqs_sdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_1 = %b", i_dqs_sdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dqs_sdr_lpde_cfg_0 = %b", i_dqs_sdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dqs_rgb_mode_7 = %b", i_dqs_rgb_mode[7]);
   $fdisplay(fd, "i_dqs_rgb_mode_6 = %b", i_dqs_rgb_mode[6]);
   $fdisplay(fd, "i_dqs_rgb_mode_5 = %b", i_dqs_rgb_mode[5]);
   $fdisplay(fd, "i_dqs_rgb_mode_4 = %b", i_dqs_rgb_mode[4]);
   $fdisplay(fd, "i_dqs_rgb_mode_3 = %b", i_dqs_rgb_mode[3]);
   $fdisplay(fd, "i_dqs_rgb_mode_2 = %b", i_dqs_rgb_mode[2]);
   $fdisplay(fd, "i_dqs_rgb_mode_1 = %b", i_dqs_rgb_mode[1]);
   $fdisplay(fd, "i_dqs_rgb_mode_0 = %b", i_dqs_rgb_mode[0]);
   $fdisplay(fd, "i_dqs_sdr_64 = %b", i_dqs_sdr[64]);
   $fdisplay(fd, "i_dqs_sdr_56 = %b", i_dqs_sdr[56]);
   $fdisplay(fd, "i_dqs_sdr_48 = %b", i_dqs_sdr[48]);
   $fdisplay(fd, "i_dqs_sdr_40 = %b", i_dqs_sdr[40]);
   $fdisplay(fd, "i_dqs_sdr_32 = %b", i_dqs_sdr[32]);
   $fdisplay(fd, "i_dqs_sdr_24 = %b", i_dqs_sdr[24]);
   $fdisplay(fd, "i_dqs_sdr_16 = %b", i_dqs_sdr[16]);
   $fdisplay(fd, "i_dqs_sdr_8 = %b", i_dqs_sdr[8]);
   $fdisplay(fd, "i_dqs_sdr_7 = %b", i_dqs_sdr[7]);
   $fdisplay(fd, "i_dqs_sdr_6 = %b", i_dqs_sdr[6]);
   $fdisplay(fd, "i_dqs_sdr_5 = %b", i_dqs_sdr[5]);
   $fdisplay(fd, "i_dqs_sdr_4 = %b", i_dqs_sdr[4]);
   $fdisplay(fd, "i_dqs_sdr_3 = %b", i_dqs_sdr[3]);
   $fdisplay(fd, "i_dqs_sdr_2 = %b", i_dqs_sdr[2]);
   $fdisplay(fd, "i_dqs_sdr_1 = %b", i_dqs_sdr[1]);
   $fdisplay(fd, "i_dqs_sdr_0 = %b", i_dqs_sdr[0]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_33 = %b", i_dqs_sdr_rt_pi_cfg[33]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_32 = %b", i_dqs_sdr_rt_pi_cfg[32]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_31 = %b", i_dqs_sdr_rt_pi_cfg[31]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_30 = %b", i_dqs_sdr_rt_pi_cfg[30]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_29 = %b", i_dqs_sdr_rt_pi_cfg[29]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_28 = %b", i_dqs_sdr_rt_pi_cfg[28]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_27 = %b", i_dqs_sdr_rt_pi_cfg[27]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_26 = %b", i_dqs_sdr_rt_pi_cfg[26]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_25 = %b", i_dqs_sdr_rt_pi_cfg[25]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_24 = %b", i_dqs_sdr_rt_pi_cfg[24]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_23 = %b", i_dqs_sdr_rt_pi_cfg[23]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_22 = %b", i_dqs_sdr_rt_pi_cfg[22]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_21 = %b", i_dqs_sdr_rt_pi_cfg[21]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_20 = %b", i_dqs_sdr_rt_pi_cfg[20]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_19 = %b", i_dqs_sdr_rt_pi_cfg[19]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_18 = %b", i_dqs_sdr_rt_pi_cfg[18]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_17 = %b", i_dqs_sdr_rt_pi_cfg[17]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_16 = %b", i_dqs_sdr_rt_pi_cfg[16]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_14 = %b", i_dqs_sdr_rt_pi_cfg[14]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_13 = %b", i_dqs_sdr_rt_pi_cfg[13]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_12 = %b", i_dqs_sdr_rt_pi_cfg[12]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_11 = %b", i_dqs_sdr_rt_pi_cfg[11]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_10 = %b", i_dqs_sdr_rt_pi_cfg[10]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_9 = %b", i_dqs_sdr_rt_pi_cfg[9]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_8 = %b", i_dqs_sdr_rt_pi_cfg[8]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_7 = %b", i_dqs_sdr_rt_pi_cfg[7]);
   $fdisplay(fd, "i_dqs_sdr_rt_pi_cfg_6 = %b", i_dqs_sdr_rt_pi_cfg[6]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_33 = %b", i_dqs_ddr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_32 = %b", i_dqs_ddr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_31 = %b", i_dqs_ddr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_30 = %b", i_dqs_ddr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_29 = %b", i_dqs_ddr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_28 = %b", i_dqs_ddr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_27 = %b", i_dqs_ddr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_26 = %b", i_dqs_ddr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_25 = %b", i_dqs_ddr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_24 = %b", i_dqs_ddr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_23 = %b", i_dqs_ddr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_22 = %b", i_dqs_ddr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_21 = %b", i_dqs_ddr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_20 = %b", i_dqs_ddr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_19 = %b", i_dqs_ddr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_18 = %b", i_dqs_ddr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_17 = %b", i_dqs_ddr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_16 = %b", i_dqs_ddr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_14 = %b", i_dqs_ddr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_13 = %b", i_dqs_ddr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_12 = %b", i_dqs_ddr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_11 = %b", i_dqs_ddr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_10 = %b", i_dqs_ddr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_9 = %b", i_dqs_ddr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_8 = %b", i_dqs_ddr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_7 = %b", i_dqs_ddr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dqs_ddr_pi_0_cfg_6 = %b", i_dqs_ddr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_33 = %b", i_dqs_qdr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_32 = %b", i_dqs_qdr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_31 = %b", i_dqs_qdr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_30 = %b", i_dqs_qdr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_29 = %b", i_dqs_qdr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_28 = %b", i_dqs_qdr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_27 = %b", i_dqs_qdr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_26 = %b", i_dqs_qdr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_25 = %b", i_dqs_qdr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_24 = %b", i_dqs_qdr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_23 = %b", i_dqs_qdr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_22 = %b", i_dqs_qdr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_21 = %b", i_dqs_qdr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_20 = %b", i_dqs_qdr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_19 = %b", i_dqs_qdr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_18 = %b", i_dqs_qdr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_17 = %b", i_dqs_qdr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_16 = %b", i_dqs_qdr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_14 = %b", i_dqs_qdr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_13 = %b", i_dqs_qdr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_12 = %b", i_dqs_qdr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_11 = %b", i_dqs_qdr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_10 = %b", i_dqs_qdr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_9 = %b", i_dqs_qdr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_8 = %b", i_dqs_qdr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_7 = %b", i_dqs_qdr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dqs_qdr_pi_0_cfg_6 = %b", i_dqs_qdr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_8 = %b", i_dqs_xdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_7 = %b", i_dqs_xdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_6 = %b", i_dqs_xdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_5 = %b", i_dqs_xdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_4 = %b", i_dqs_xdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_3 = %b", i_dqs_xdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_2 = %b", i_dqs_xdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_1 = %b", i_dqs_xdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dqs_xdr_lpde_cfg_0 = %b", i_dqs_xdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dqs_ddr_1_pipe_en_0 = %b", i_dqs_ddr_1_pipe_en[0]);
   $fdisplay(fd, "i_dqs_ddr_1_x_sel_0 = %b", i_dqs_ddr_1_x_sel[0]);
   $fdisplay(fd, "i_dqs_ddr_0_pipe_en_0 = %b", i_dqs_ddr_0_pipe_en[0]);
   $fdisplay(fd, "i_dqs_ddr_0_x_sel_0 = %b", i_dqs_ddr_0_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_3_pipe_en_0 = %b", i_dqs_sdr_3_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_1 = %b", i_dqs_sdr_3_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_3_x_sel_0 = %b", i_dqs_sdr_3_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_1 = %b", i_dqs_sdr_3_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_3_fc_dly_0 = %b", i_dqs_sdr_3_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_2_pipe_en_0 = %b", i_dqs_sdr_2_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_1 = %b", i_dqs_sdr_2_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_2_x_sel_0 = %b", i_dqs_sdr_2_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_1 = %b", i_dqs_sdr_2_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_2_fc_dly_0 = %b", i_dqs_sdr_2_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_1_pipe_en_0 = %b", i_dqs_sdr_1_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_1 = %b", i_dqs_sdr_1_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_1_x_sel_0 = %b", i_dqs_sdr_1_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_1 = %b", i_dqs_sdr_1_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_1_fc_dly_0 = %b", i_dqs_sdr_1_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_0_pipe_en_0 = %b", i_dqs_sdr_0_pipe_en[0]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_1 = %b", i_dqs_sdr_0_x_sel[1]);
   $fdisplay(fd, "i_dqs_sdr_0_x_sel_0 = %b", i_dqs_sdr_0_x_sel[0]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_1 = %b", i_dqs_sdr_0_fc_dly[1]);
   $fdisplay(fd, "i_dqs_sdr_0_fc_dly_0 = %b", i_dqs_sdr_0_fc_dly[0]);
   $fdisplay(fd, "i_dqs_sdr_rt_pipe_en_0 = %b", i_dqs_sdr_rt_pipe_en[0]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_3 = %b", i_dfirdclk_en_pulse_ext[3]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_2 = %b", i_dfirdclk_en_pulse_ext[2]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_1 = %b", i_dfirdclk_en_pulse_ext[1]);
   $fdisplay(fd, "i_dfirdclk_en_pulse_ext_0 = %b", i_dfirdclk_en_pulse_ext[0]);
   $fdisplay(fd, "i_dfirdclk_en = %b", i_dfirdclk_en);
   $fdisplay(fd, "i_dq_dfi_wrtraffic = %b", i_dq_dfi_wrtraffic);
   $fdisplay(fd, "i_dqs_dfi_wrtraffic = %b", i_dqs_dfi_wrtraffic);
   $fdisplay(fd, "i_csp_div_rst_n = %b", i_csp_div_rst_n);
   $fdisplay(fd, "i_dqs_ck2wck_ratio_2 = %b", i_dqs_ck2wck_ratio[2]);
   $fdisplay(fd, "i_dqs_ck2wck_ratio_1 = %b", i_dqs_ck2wck_ratio[1]);
   $fdisplay(fd, "i_dqs_wgb_mode_8 = %b", i_dqs_wgb_mode[8]);
   $fdisplay(fd, "i_dqs_tgb_mode_7 = %b", i_dqs_tgb_mode[7]);
   $fdisplay(fd, "i_dqs_tgb_mode_6 = %b", i_dqs_tgb_mode[6]);
   $fdisplay(fd, "i_dqs_tgb_mode_4 = %b", i_dqs_tgb_mode[4]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_6 = %b", i_dqs_egress_mode_dig[6]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_1 = %b", i_dqs_egress_mode_dig[1]);
   $fdisplay(fd, "i_dqs_egress_mode_dig_0 = %b", i_dqs_egress_mode_dig[0]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_2 = %b", i_dqs_egress_mode_ana[2]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_1 = %b", i_dqs_egress_mode_ana[1]);
   $fdisplay(fd, "i_dqs_egress_mode_ana_0 = %b", i_dqs_egress_mode_ana[0]);
   $fdisplay(fd, "i_dq_sdr_87 = %b", i_dq_sdr[87]);
   $fdisplay(fd, "i_dq_sdr_86 = %b", i_dq_sdr[86]);
   $fdisplay(fd, "i_dq_sdr_85 = %b", i_dq_sdr[85]);
   $fdisplay(fd, "i_dq_sdr_84 = %b", i_dq_sdr[84]);
   $fdisplay(fd, "i_dq_sdr_83 = %b", i_dq_sdr[83]);
   $fdisplay(fd, "i_dq_sdr_82 = %b", i_dq_sdr[82]);
   $fdisplay(fd, "i_dq_sdr_81 = %b", i_dq_sdr[81]);
   $fdisplay(fd, "i_dq_sdr_80 = %b", i_dq_sdr[80]);
   $fdisplay(fd, "i_dq_sdr_79 = %b", i_dq_sdr[79]);
   $fdisplay(fd, "i_dq_sdr_78 = %b", i_dq_sdr[78]);
   $fdisplay(fd, "i_dq_sdr_77 = %b", i_dq_sdr[77]);
   $fdisplay(fd, "i_dq_sdr_76 = %b", i_dq_sdr[76]);
   $fdisplay(fd, "i_dq_sdr_75 = %b", i_dq_sdr[75]);
   $fdisplay(fd, "i_dq_sdr_74 = %b", i_dq_sdr[74]);
   $fdisplay(fd, "i_dq_sdr_73 = %b", i_dq_sdr[73]);
   $fdisplay(fd, "i_dq_sdr_72 = %b", i_dq_sdr[72]);
   $fdisplay(fd, "i_dq_sdr_71 = %b", i_dq_sdr[71]);
   $fdisplay(fd, "i_dq_sdr_70 = %b", i_dq_sdr[70]);
   $fdisplay(fd, "i_dq_sdr_69 = %b", i_dq_sdr[69]);
   $fdisplay(fd, "i_dq_sdr_68 = %b", i_dq_sdr[68]);
   $fdisplay(fd, "i_dq_sdr_67 = %b", i_dq_sdr[67]);
   $fdisplay(fd, "i_dq_sdr_66 = %b", i_dq_sdr[66]);
   $fdisplay(fd, "i_dq_sdr_65 = %b", i_dq_sdr[65]);
   $fdisplay(fd, "i_dq_sdr_64 = %b", i_dq_sdr[64]);
   $fdisplay(fd, "i_dq_sdr_63 = %b", i_dq_sdr[63]);
   $fdisplay(fd, "i_dq_sdr_62 = %b", i_dq_sdr[62]);
   $fdisplay(fd, "i_dq_sdr_61 = %b", i_dq_sdr[61]);
   $fdisplay(fd, "i_dq_sdr_60 = %b", i_dq_sdr[60]);
   $fdisplay(fd, "i_dq_sdr_59 = %b", i_dq_sdr[59]);
   $fdisplay(fd, "i_dq_sdr_58 = %b", i_dq_sdr[58]);
   $fdisplay(fd, "i_dq_sdr_57 = %b", i_dq_sdr[57]);
   $fdisplay(fd, "i_dq_sdr_56 = %b", i_dq_sdr[56]);
   $fdisplay(fd, "i_dq_sdr_55 = %b", i_dq_sdr[55]);
   $fdisplay(fd, "i_dq_sdr_54 = %b", i_dq_sdr[54]);
   $fdisplay(fd, "i_dq_sdr_53 = %b", i_dq_sdr[53]);
   $fdisplay(fd, "i_dq_sdr_52 = %b", i_dq_sdr[52]);
   $fdisplay(fd, "i_dq_sdr_51 = %b", i_dq_sdr[51]);
   $fdisplay(fd, "i_dq_sdr_50 = %b", i_dq_sdr[50]);
   $fdisplay(fd, "i_dq_sdr_49 = %b", i_dq_sdr[49]);
   $fdisplay(fd, "i_dq_sdr_48 = %b", i_dq_sdr[48]);
   $fdisplay(fd, "i_dq_sdr_47 = %b", i_dq_sdr[47]);
   $fdisplay(fd, "i_dq_sdr_46 = %b", i_dq_sdr[46]);
   $fdisplay(fd, "i_dq_sdr_45 = %b", i_dq_sdr[45]);
   $fdisplay(fd, "i_dq_sdr_44 = %b", i_dq_sdr[44]);
   $fdisplay(fd, "i_dq_sdr_43 = %b", i_dq_sdr[43]);
   $fdisplay(fd, "i_dq_sdr_42 = %b", i_dq_sdr[42]);
   $fdisplay(fd, "i_dq_sdr_41 = %b", i_dq_sdr[41]);
   $fdisplay(fd, "i_dq_sdr_40 = %b", i_dq_sdr[40]);
   $fdisplay(fd, "i_dq_sdr_39 = %b", i_dq_sdr[39]);
   $fdisplay(fd, "i_dq_sdr_38 = %b", i_dq_sdr[38]);
   $fdisplay(fd, "i_dq_sdr_37 = %b", i_dq_sdr[37]);
   $fdisplay(fd, "i_dq_sdr_36 = %b", i_dq_sdr[36]);
   $fdisplay(fd, "i_dq_sdr_35 = %b", i_dq_sdr[35]);
   $fdisplay(fd, "i_dq_sdr_34 = %b", i_dq_sdr[34]);
   $fdisplay(fd, "i_dq_sdr_33 = %b", i_dq_sdr[33]);
   $fdisplay(fd, "i_dq_sdr_32 = %b", i_dq_sdr[32]);
   $fdisplay(fd, "i_dq_sdr_31 = %b", i_dq_sdr[31]);
   $fdisplay(fd, "i_dq_sdr_30 = %b", i_dq_sdr[30]);
   $fdisplay(fd, "i_dq_sdr_29 = %b", i_dq_sdr[29]);
   $fdisplay(fd, "i_dq_sdr_28 = %b", i_dq_sdr[28]);
   $fdisplay(fd, "i_dq_sdr_27 = %b", i_dq_sdr[27]);
   $fdisplay(fd, "i_dq_sdr_26 = %b", i_dq_sdr[26]);
   $fdisplay(fd, "i_dq_sdr_25 = %b", i_dq_sdr[25]);
   $fdisplay(fd, "i_dq_sdr_24 = %b", i_dq_sdr[24]);
   $fdisplay(fd, "i_dq_sdr_23 = %b", i_dq_sdr[23]);
   $fdisplay(fd, "i_dq_sdr_22 = %b", i_dq_sdr[22]);
   $fdisplay(fd, "i_dq_sdr_21 = %b", i_dq_sdr[21]);
   $fdisplay(fd, "i_dq_sdr_20 = %b", i_dq_sdr[20]);
   $fdisplay(fd, "i_dq_sdr_19 = %b", i_dq_sdr[19]);
   $fdisplay(fd, "i_dq_sdr_18 = %b", i_dq_sdr[18]);
   $fdisplay(fd, "i_dq_sdr_17 = %b", i_dq_sdr[17]);
   $fdisplay(fd, "i_dq_sdr_16 = %b", i_dq_sdr[16]);
   $fdisplay(fd, "i_dq_sdr_15 = %b", i_dq_sdr[15]);
   $fdisplay(fd, "i_dq_sdr_14 = %b", i_dq_sdr[14]);
   $fdisplay(fd, "i_dq_sdr_13 = %b", i_dq_sdr[13]);
   $fdisplay(fd, "i_dq_sdr_12 = %b", i_dq_sdr[12]);
   $fdisplay(fd, "i_dq_sdr_11 = %b", i_dq_sdr[11]);
   $fdisplay(fd, "i_dq_sdr_10 = %b", i_dq_sdr[10]);
   $fdisplay(fd, "i_dq_sdr_9 = %b", i_dq_sdr[9]);
   $fdisplay(fd, "i_dq_sdr_8 = %b", i_dq_sdr[8]);
   $fdisplay(fd, "i_dq_sdr_7 = %b", i_dq_sdr[7]);
   $fdisplay(fd, "i_dq_sdr_6 = %b", i_dq_sdr[6]);
   $fdisplay(fd, "i_dq_sdr_5 = %b", i_dq_sdr[5]);
   $fdisplay(fd, "i_dq_sdr_4 = %b", i_dq_sdr[4]);
   $fdisplay(fd, "i_dq_sdr_3 = %b", i_dq_sdr[3]);
   $fdisplay(fd, "i_dq_sdr_2 = %b", i_dq_sdr[2]);
   $fdisplay(fd, "i_dq_sdr_1 = %b", i_dq_sdr[1]);
   $fdisplay(fd, "i_dq_sdr_0 = %b", i_dq_sdr[0]);
   $fdisplay(fd, "i_dfi_pi_cfg_14 = %b", i_dfi_pi_cfg[14]);
   $fdisplay(fd, "i_dfi_pi_cfg_13 = %b", i_dfi_pi_cfg[13]);
   $fdisplay(fd, "i_dfi_pi_cfg_12 = %b", i_dfi_pi_cfg[12]);
   $fdisplay(fd, "i_dfi_pi_cfg_11 = %b", i_dfi_pi_cfg[11]);
   $fdisplay(fd, "i_dfi_pi_cfg_10 = %b", i_dfi_pi_cfg[10]);
   $fdisplay(fd, "i_dfi_pi_cfg_9 = %b", i_dfi_pi_cfg[9]);
   $fdisplay(fd, "i_dfi_pi_cfg_8 = %b", i_dfi_pi_cfg[8]);
   $fdisplay(fd, "i_dfi_pi_cfg_7 = %b", i_dfi_pi_cfg[7]);
   $fdisplay(fd, "i_dfi_pi_cfg_6 = %b", i_dfi_pi_cfg[6]);
   $fdisplay(fd, "i_sdr_pi_cfg_14 = %b", i_sdr_pi_cfg[14]);
   $fdisplay(fd, "i_sdr_pi_cfg_13 = %b", i_sdr_pi_cfg[13]);
   $fdisplay(fd, "i_sdr_pi_cfg_12 = %b", i_sdr_pi_cfg[12]);
   $fdisplay(fd, "i_sdr_pi_cfg_11 = %b", i_sdr_pi_cfg[11]);
   $fdisplay(fd, "i_sdr_pi_cfg_10 = %b", i_sdr_pi_cfg[10]);
   $fdisplay(fd, "i_sdr_pi_cfg_9 = %b", i_sdr_pi_cfg[9]);
   $fdisplay(fd, "i_sdr_pi_cfg_8 = %b", i_sdr_pi_cfg[8]);
   $fdisplay(fd, "i_sdr_pi_cfg_7 = %b", i_sdr_pi_cfg[7]);
   $fdisplay(fd, "i_sdr_pi_cfg_6 = %b", i_sdr_pi_cfg[6]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_33 = %b", i_dq_sdr_rt_pi_cfg[33]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_32 = %b", i_dq_sdr_rt_pi_cfg[32]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_31 = %b", i_dq_sdr_rt_pi_cfg[31]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_30 = %b", i_dq_sdr_rt_pi_cfg[30]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_29 = %b", i_dq_sdr_rt_pi_cfg[29]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_28 = %b", i_dq_sdr_rt_pi_cfg[28]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_27 = %b", i_dq_sdr_rt_pi_cfg[27]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_26 = %b", i_dq_sdr_rt_pi_cfg[26]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_25 = %b", i_dq_sdr_rt_pi_cfg[25]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_24 = %b", i_dq_sdr_rt_pi_cfg[24]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_23 = %b", i_dq_sdr_rt_pi_cfg[23]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_22 = %b", i_dq_sdr_rt_pi_cfg[22]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_21 = %b", i_dq_sdr_rt_pi_cfg[21]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_20 = %b", i_dq_sdr_rt_pi_cfg[20]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_19 = %b", i_dq_sdr_rt_pi_cfg[19]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_18 = %b", i_dq_sdr_rt_pi_cfg[18]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_17 = %b", i_dq_sdr_rt_pi_cfg[17]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_16 = %b", i_dq_sdr_rt_pi_cfg[16]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_14 = %b", i_dq_sdr_rt_pi_cfg[14]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_13 = %b", i_dq_sdr_rt_pi_cfg[13]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_12 = %b", i_dq_sdr_rt_pi_cfg[12]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_11 = %b", i_dq_sdr_rt_pi_cfg[11]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_10 = %b", i_dq_sdr_rt_pi_cfg[10]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_9 = %b", i_dq_sdr_rt_pi_cfg[9]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_8 = %b", i_dq_sdr_rt_pi_cfg[8]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_7 = %b", i_dq_sdr_rt_pi_cfg[7]);
   $fdisplay(fd, "i_dq_sdr_rt_pi_cfg_6 = %b", i_dq_sdr_rt_pi_cfg[6]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_33 = %b", i_dq_ddr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_32 = %b", i_dq_ddr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_31 = %b", i_dq_ddr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_30 = %b", i_dq_ddr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_29 = %b", i_dq_ddr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_28 = %b", i_dq_ddr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_27 = %b", i_dq_ddr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_26 = %b", i_dq_ddr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_25 = %b", i_dq_ddr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_24 = %b", i_dq_ddr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_23 = %b", i_dq_ddr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_22 = %b", i_dq_ddr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_21 = %b", i_dq_ddr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_20 = %b", i_dq_ddr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_19 = %b", i_dq_ddr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_18 = %b", i_dq_ddr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_17 = %b", i_dq_ddr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_16 = %b", i_dq_ddr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_14 = %b", i_dq_ddr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_13 = %b", i_dq_ddr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_12 = %b", i_dq_ddr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_11 = %b", i_dq_ddr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_10 = %b", i_dq_ddr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_9 = %b", i_dq_ddr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_8 = %b", i_dq_ddr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_7 = %b", i_dq_ddr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dq_ddr_pi_0_cfg_6 = %b", i_dq_ddr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_33 = %b", i_dq_qdr_pi_0_cfg[33]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_32 = %b", i_dq_qdr_pi_0_cfg[32]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_31 = %b", i_dq_qdr_pi_0_cfg[31]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_30 = %b", i_dq_qdr_pi_0_cfg[30]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_29 = %b", i_dq_qdr_pi_0_cfg[29]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_28 = %b", i_dq_qdr_pi_0_cfg[28]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_27 = %b", i_dq_qdr_pi_0_cfg[27]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_26 = %b", i_dq_qdr_pi_0_cfg[26]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_25 = %b", i_dq_qdr_pi_0_cfg[25]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_24 = %b", i_dq_qdr_pi_0_cfg[24]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_23 = %b", i_dq_qdr_pi_0_cfg[23]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_22 = %b", i_dq_qdr_pi_0_cfg[22]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_21 = %b", i_dq_qdr_pi_0_cfg[21]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_20 = %b", i_dq_qdr_pi_0_cfg[20]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_19 = %b", i_dq_qdr_pi_0_cfg[19]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_18 = %b", i_dq_qdr_pi_0_cfg[18]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_17 = %b", i_dq_qdr_pi_0_cfg[17]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_16 = %b", i_dq_qdr_pi_0_cfg[16]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_14 = %b", i_dq_qdr_pi_0_cfg[14]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_13 = %b", i_dq_qdr_pi_0_cfg[13]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_12 = %b", i_dq_qdr_pi_0_cfg[12]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_11 = %b", i_dq_qdr_pi_0_cfg[11]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_10 = %b", i_dq_qdr_pi_0_cfg[10]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_9 = %b", i_dq_qdr_pi_0_cfg[9]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_8 = %b", i_dq_qdr_pi_0_cfg[8]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_7 = %b", i_dq_qdr_pi_0_cfg[7]);
   $fdisplay(fd, "i_dq_qdr_pi_0_cfg_6 = %b", i_dq_qdr_pi_0_cfg[6]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_98 = %b", i_dq_xdr_lpde_cfg[98]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_97 = %b", i_dq_xdr_lpde_cfg[97]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_96 = %b", i_dq_xdr_lpde_cfg[96]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_95 = %b", i_dq_xdr_lpde_cfg[95]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_94 = %b", i_dq_xdr_lpde_cfg[94]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_93 = %b", i_dq_xdr_lpde_cfg[93]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_92 = %b", i_dq_xdr_lpde_cfg[92]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_91 = %b", i_dq_xdr_lpde_cfg[91]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_90 = %b", i_dq_xdr_lpde_cfg[90]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_89 = %b", i_dq_xdr_lpde_cfg[89]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_88 = %b", i_dq_xdr_lpde_cfg[88]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_87 = %b", i_dq_xdr_lpde_cfg[87]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_86 = %b", i_dq_xdr_lpde_cfg[86]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_85 = %b", i_dq_xdr_lpde_cfg[85]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_84 = %b", i_dq_xdr_lpde_cfg[84]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_83 = %b", i_dq_xdr_lpde_cfg[83]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_82 = %b", i_dq_xdr_lpde_cfg[82]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_81 = %b", i_dq_xdr_lpde_cfg[81]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_80 = %b", i_dq_xdr_lpde_cfg[80]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_79 = %b", i_dq_xdr_lpde_cfg[79]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_78 = %b", i_dq_xdr_lpde_cfg[78]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_77 = %b", i_dq_xdr_lpde_cfg[77]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_76 = %b", i_dq_xdr_lpde_cfg[76]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_75 = %b", i_dq_xdr_lpde_cfg[75]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_74 = %b", i_dq_xdr_lpde_cfg[74]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_73 = %b", i_dq_xdr_lpde_cfg[73]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_72 = %b", i_dq_xdr_lpde_cfg[72]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_71 = %b", i_dq_xdr_lpde_cfg[71]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_70 = %b", i_dq_xdr_lpde_cfg[70]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_69 = %b", i_dq_xdr_lpde_cfg[69]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_68 = %b", i_dq_xdr_lpde_cfg[68]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_67 = %b", i_dq_xdr_lpde_cfg[67]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_66 = %b", i_dq_xdr_lpde_cfg[66]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_65 = %b", i_dq_xdr_lpde_cfg[65]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_64 = %b", i_dq_xdr_lpde_cfg[64]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_63 = %b", i_dq_xdr_lpde_cfg[63]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_62 = %b", i_dq_xdr_lpde_cfg[62]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_61 = %b", i_dq_xdr_lpde_cfg[61]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_60 = %b", i_dq_xdr_lpde_cfg[60]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_59 = %b", i_dq_xdr_lpde_cfg[59]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_58 = %b", i_dq_xdr_lpde_cfg[58]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_57 = %b", i_dq_xdr_lpde_cfg[57]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_56 = %b", i_dq_xdr_lpde_cfg[56]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_55 = %b", i_dq_xdr_lpde_cfg[55]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_54 = %b", i_dq_xdr_lpde_cfg[54]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_53 = %b", i_dq_xdr_lpde_cfg[53]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_52 = %b", i_dq_xdr_lpde_cfg[52]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_51 = %b", i_dq_xdr_lpde_cfg[51]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_50 = %b", i_dq_xdr_lpde_cfg[50]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_49 = %b", i_dq_xdr_lpde_cfg[49]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_48 = %b", i_dq_xdr_lpde_cfg[48]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_47 = %b", i_dq_xdr_lpde_cfg[47]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_46 = %b", i_dq_xdr_lpde_cfg[46]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_45 = %b", i_dq_xdr_lpde_cfg[45]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_44 = %b", i_dq_xdr_lpde_cfg[44]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_43 = %b", i_dq_xdr_lpde_cfg[43]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_42 = %b", i_dq_xdr_lpde_cfg[42]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_41 = %b", i_dq_xdr_lpde_cfg[41]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_40 = %b", i_dq_xdr_lpde_cfg[40]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_39 = %b", i_dq_xdr_lpde_cfg[39]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_38 = %b", i_dq_xdr_lpde_cfg[38]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_37 = %b", i_dq_xdr_lpde_cfg[37]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_36 = %b", i_dq_xdr_lpde_cfg[36]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_35 = %b", i_dq_xdr_lpde_cfg[35]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_34 = %b", i_dq_xdr_lpde_cfg[34]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_33 = %b", i_dq_xdr_lpde_cfg[33]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_32 = %b", i_dq_xdr_lpde_cfg[32]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_31 = %b", i_dq_xdr_lpde_cfg[31]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_30 = %b", i_dq_xdr_lpde_cfg[30]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_29 = %b", i_dq_xdr_lpde_cfg[29]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_28 = %b", i_dq_xdr_lpde_cfg[28]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_27 = %b", i_dq_xdr_lpde_cfg[27]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_26 = %b", i_dq_xdr_lpde_cfg[26]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_25 = %b", i_dq_xdr_lpde_cfg[25]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_24 = %b", i_dq_xdr_lpde_cfg[24]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_23 = %b", i_dq_xdr_lpde_cfg[23]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_22 = %b", i_dq_xdr_lpde_cfg[22]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_21 = %b", i_dq_xdr_lpde_cfg[21]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_20 = %b", i_dq_xdr_lpde_cfg[20]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_19 = %b", i_dq_xdr_lpde_cfg[19]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_18 = %b", i_dq_xdr_lpde_cfg[18]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_17 = %b", i_dq_xdr_lpde_cfg[17]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_16 = %b", i_dq_xdr_lpde_cfg[16]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_15 = %b", i_dq_xdr_lpde_cfg[15]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_14 = %b", i_dq_xdr_lpde_cfg[14]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_13 = %b", i_dq_xdr_lpde_cfg[13]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_12 = %b", i_dq_xdr_lpde_cfg[12]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_11 = %b", i_dq_xdr_lpde_cfg[11]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_10 = %b", i_dq_xdr_lpde_cfg[10]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_9 = %b", i_dq_xdr_lpde_cfg[9]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_8 = %b", i_dq_xdr_lpde_cfg[8]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_7 = %b", i_dq_xdr_lpde_cfg[7]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_6 = %b", i_dq_xdr_lpde_cfg[6]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_5 = %b", i_dq_xdr_lpde_cfg[5]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_4 = %b", i_dq_xdr_lpde_cfg[4]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_3 = %b", i_dq_xdr_lpde_cfg[3]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_2 = %b", i_dq_xdr_lpde_cfg[2]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_1 = %b", i_dq_xdr_lpde_cfg[1]);
   $fdisplay(fd, "i_dq_xdr_lpde_cfg_0 = %b", i_dq_xdr_lpde_cfg[0]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_10 = %b", i_dq_ddr_1_pipe_en[10]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_9 = %b", i_dq_ddr_1_pipe_en[9]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_8 = %b", i_dq_ddr_1_pipe_en[8]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_7 = %b", i_dq_ddr_1_pipe_en[7]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_6 = %b", i_dq_ddr_1_pipe_en[6]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_5 = %b", i_dq_ddr_1_pipe_en[5]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_4 = %b", i_dq_ddr_1_pipe_en[4]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_3 = %b", i_dq_ddr_1_pipe_en[3]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_2 = %b", i_dq_ddr_1_pipe_en[2]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_1 = %b", i_dq_ddr_1_pipe_en[1]);
   $fdisplay(fd, "i_dq_ddr_1_pipe_en_0 = %b", i_dq_ddr_1_pipe_en[0]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_20 = %b", i_dq_ddr_1_x_sel[20]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_18 = %b", i_dq_ddr_1_x_sel[18]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_16 = %b", i_dq_ddr_1_x_sel[16]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_14 = %b", i_dq_ddr_1_x_sel[14]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_12 = %b", i_dq_ddr_1_x_sel[12]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_10 = %b", i_dq_ddr_1_x_sel[10]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_8 = %b", i_dq_ddr_1_x_sel[8]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_6 = %b", i_dq_ddr_1_x_sel[6]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_4 = %b", i_dq_ddr_1_x_sel[4]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_2 = %b", i_dq_ddr_1_x_sel[2]);
   $fdisplay(fd, "i_dq_ddr_1_x_sel_0 = %b", i_dq_ddr_1_x_sel[0]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_10 = %b", i_dq_ddr_0_pipe_en[10]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_9 = %b", i_dq_ddr_0_pipe_en[9]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_8 = %b", i_dq_ddr_0_pipe_en[8]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_7 = %b", i_dq_ddr_0_pipe_en[7]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_6 = %b", i_dq_ddr_0_pipe_en[6]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_5 = %b", i_dq_ddr_0_pipe_en[5]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_4 = %b", i_dq_ddr_0_pipe_en[4]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_3 = %b", i_dq_ddr_0_pipe_en[3]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_2 = %b", i_dq_ddr_0_pipe_en[2]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_1 = %b", i_dq_ddr_0_pipe_en[1]);
   $fdisplay(fd, "i_dq_ddr_0_pipe_en_0 = %b", i_dq_ddr_0_pipe_en[0]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_20 = %b", i_dq_ddr_0_x_sel[20]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_18 = %b", i_dq_ddr_0_x_sel[18]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_16 = %b", i_dq_ddr_0_x_sel[16]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_14 = %b", i_dq_ddr_0_x_sel[14]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_12 = %b", i_dq_ddr_0_x_sel[12]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_10 = %b", i_dq_ddr_0_x_sel[10]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_8 = %b", i_dq_ddr_0_x_sel[8]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_6 = %b", i_dq_ddr_0_x_sel[6]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_4 = %b", i_dq_ddr_0_x_sel[4]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_2 = %b", i_dq_ddr_0_x_sel[2]);
   $fdisplay(fd, "i_dq_ddr_0_x_sel_0 = %b", i_dq_ddr_0_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_10 = %b", i_dq_sdr_3_pipe_en[10]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_9 = %b", i_dq_sdr_3_pipe_en[9]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_8 = %b", i_dq_sdr_3_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_7 = %b", i_dq_sdr_3_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_6 = %b", i_dq_sdr_3_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_5 = %b", i_dq_sdr_3_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_4 = %b", i_dq_sdr_3_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_3 = %b", i_dq_sdr_3_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_2 = %b", i_dq_sdr_3_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_1 = %b", i_dq_sdr_3_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_3_pipe_en_0 = %b", i_dq_sdr_3_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_31 = %b", i_dq_sdr_3_x_sel[31]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_30 = %b", i_dq_sdr_3_x_sel[30]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_28 = %b", i_dq_sdr_3_x_sel[28]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_27 = %b", i_dq_sdr_3_x_sel[27]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_25 = %b", i_dq_sdr_3_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_24 = %b", i_dq_sdr_3_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_22 = %b", i_dq_sdr_3_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_21 = %b", i_dq_sdr_3_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_19 = %b", i_dq_sdr_3_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_18 = %b", i_dq_sdr_3_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_16 = %b", i_dq_sdr_3_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_15 = %b", i_dq_sdr_3_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_13 = %b", i_dq_sdr_3_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_12 = %b", i_dq_sdr_3_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_10 = %b", i_dq_sdr_3_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_9 = %b", i_dq_sdr_3_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_7 = %b", i_dq_sdr_3_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_6 = %b", i_dq_sdr_3_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_4 = %b", i_dq_sdr_3_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_3 = %b", i_dq_sdr_3_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_1 = %b", i_dq_sdr_3_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_3_x_sel_0 = %b", i_dq_sdr_3_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_21 = %b", i_dq_sdr_3_fc_dly[21]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_20 = %b", i_dq_sdr_3_fc_dly[20]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_19 = %b", i_dq_sdr_3_fc_dly[19]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_18 = %b", i_dq_sdr_3_fc_dly[18]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_17 = %b", i_dq_sdr_3_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_16 = %b", i_dq_sdr_3_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_15 = %b", i_dq_sdr_3_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_14 = %b", i_dq_sdr_3_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_13 = %b", i_dq_sdr_3_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_12 = %b", i_dq_sdr_3_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_11 = %b", i_dq_sdr_3_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_10 = %b", i_dq_sdr_3_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_9 = %b", i_dq_sdr_3_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_8 = %b", i_dq_sdr_3_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_7 = %b", i_dq_sdr_3_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_6 = %b", i_dq_sdr_3_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_5 = %b", i_dq_sdr_3_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_4 = %b", i_dq_sdr_3_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_3 = %b", i_dq_sdr_3_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_2 = %b", i_dq_sdr_3_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_1 = %b", i_dq_sdr_3_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_3_fc_dly_0 = %b", i_dq_sdr_3_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_10 = %b", i_dq_sdr_2_pipe_en[10]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_9 = %b", i_dq_sdr_2_pipe_en[9]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_8 = %b", i_dq_sdr_2_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_7 = %b", i_dq_sdr_2_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_6 = %b", i_dq_sdr_2_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_5 = %b", i_dq_sdr_2_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_4 = %b", i_dq_sdr_2_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_3 = %b", i_dq_sdr_2_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_2 = %b", i_dq_sdr_2_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_1 = %b", i_dq_sdr_2_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_2_pipe_en_0 = %b", i_dq_sdr_2_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_31 = %b", i_dq_sdr_2_x_sel[31]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_30 = %b", i_dq_sdr_2_x_sel[30]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_28 = %b", i_dq_sdr_2_x_sel[28]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_27 = %b", i_dq_sdr_2_x_sel[27]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_25 = %b", i_dq_sdr_2_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_24 = %b", i_dq_sdr_2_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_22 = %b", i_dq_sdr_2_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_21 = %b", i_dq_sdr_2_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_19 = %b", i_dq_sdr_2_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_18 = %b", i_dq_sdr_2_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_16 = %b", i_dq_sdr_2_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_15 = %b", i_dq_sdr_2_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_13 = %b", i_dq_sdr_2_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_12 = %b", i_dq_sdr_2_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_10 = %b", i_dq_sdr_2_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_9 = %b", i_dq_sdr_2_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_7 = %b", i_dq_sdr_2_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_6 = %b", i_dq_sdr_2_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_4 = %b", i_dq_sdr_2_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_3 = %b", i_dq_sdr_2_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_1 = %b", i_dq_sdr_2_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_2_x_sel_0 = %b", i_dq_sdr_2_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_21 = %b", i_dq_sdr_2_fc_dly[21]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_20 = %b", i_dq_sdr_2_fc_dly[20]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_19 = %b", i_dq_sdr_2_fc_dly[19]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_18 = %b", i_dq_sdr_2_fc_dly[18]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_17 = %b", i_dq_sdr_2_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_16 = %b", i_dq_sdr_2_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_15 = %b", i_dq_sdr_2_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_14 = %b", i_dq_sdr_2_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_13 = %b", i_dq_sdr_2_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_12 = %b", i_dq_sdr_2_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_11 = %b", i_dq_sdr_2_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_10 = %b", i_dq_sdr_2_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_9 = %b", i_dq_sdr_2_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_8 = %b", i_dq_sdr_2_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_7 = %b", i_dq_sdr_2_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_6 = %b", i_dq_sdr_2_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_5 = %b", i_dq_sdr_2_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_4 = %b", i_dq_sdr_2_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_3 = %b", i_dq_sdr_2_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_2 = %b", i_dq_sdr_2_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_1 = %b", i_dq_sdr_2_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_2_fc_dly_0 = %b", i_dq_sdr_2_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_10 = %b", i_dq_sdr_1_pipe_en[10]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_9 = %b", i_dq_sdr_1_pipe_en[9]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_8 = %b", i_dq_sdr_1_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_7 = %b", i_dq_sdr_1_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_6 = %b", i_dq_sdr_1_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_5 = %b", i_dq_sdr_1_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_4 = %b", i_dq_sdr_1_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_3 = %b", i_dq_sdr_1_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_2 = %b", i_dq_sdr_1_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_1 = %b", i_dq_sdr_1_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_1_pipe_en_0 = %b", i_dq_sdr_1_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_31 = %b", i_dq_sdr_1_x_sel[31]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_30 = %b", i_dq_sdr_1_x_sel[30]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_28 = %b", i_dq_sdr_1_x_sel[28]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_27 = %b", i_dq_sdr_1_x_sel[27]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_25 = %b", i_dq_sdr_1_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_24 = %b", i_dq_sdr_1_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_22 = %b", i_dq_sdr_1_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_21 = %b", i_dq_sdr_1_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_19 = %b", i_dq_sdr_1_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_18 = %b", i_dq_sdr_1_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_16 = %b", i_dq_sdr_1_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_15 = %b", i_dq_sdr_1_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_13 = %b", i_dq_sdr_1_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_12 = %b", i_dq_sdr_1_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_10 = %b", i_dq_sdr_1_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_9 = %b", i_dq_sdr_1_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_7 = %b", i_dq_sdr_1_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_6 = %b", i_dq_sdr_1_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_4 = %b", i_dq_sdr_1_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_3 = %b", i_dq_sdr_1_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_1 = %b", i_dq_sdr_1_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_1_x_sel_0 = %b", i_dq_sdr_1_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_21 = %b", i_dq_sdr_1_fc_dly[21]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_20 = %b", i_dq_sdr_1_fc_dly[20]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_19 = %b", i_dq_sdr_1_fc_dly[19]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_18 = %b", i_dq_sdr_1_fc_dly[18]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_17 = %b", i_dq_sdr_1_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_16 = %b", i_dq_sdr_1_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_15 = %b", i_dq_sdr_1_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_14 = %b", i_dq_sdr_1_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_13 = %b", i_dq_sdr_1_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_12 = %b", i_dq_sdr_1_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_11 = %b", i_dq_sdr_1_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_10 = %b", i_dq_sdr_1_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_9 = %b", i_dq_sdr_1_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_8 = %b", i_dq_sdr_1_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_7 = %b", i_dq_sdr_1_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_6 = %b", i_dq_sdr_1_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_5 = %b", i_dq_sdr_1_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_4 = %b", i_dq_sdr_1_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_3 = %b", i_dq_sdr_1_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_2 = %b", i_dq_sdr_1_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_1 = %b", i_dq_sdr_1_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_1_fc_dly_0 = %b", i_dq_sdr_1_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_10 = %b", i_dq_sdr_0_pipe_en[10]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_9 = %b", i_dq_sdr_0_pipe_en[9]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_8 = %b", i_dq_sdr_0_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_7 = %b", i_dq_sdr_0_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_6 = %b", i_dq_sdr_0_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_5 = %b", i_dq_sdr_0_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_4 = %b", i_dq_sdr_0_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_3 = %b", i_dq_sdr_0_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_2 = %b", i_dq_sdr_0_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_1 = %b", i_dq_sdr_0_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_0_pipe_en_0 = %b", i_dq_sdr_0_pipe_en[0]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_31 = %b", i_dq_sdr_0_x_sel[31]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_30 = %b", i_dq_sdr_0_x_sel[30]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_28 = %b", i_dq_sdr_0_x_sel[28]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_27 = %b", i_dq_sdr_0_x_sel[27]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_25 = %b", i_dq_sdr_0_x_sel[25]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_24 = %b", i_dq_sdr_0_x_sel[24]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_22 = %b", i_dq_sdr_0_x_sel[22]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_21 = %b", i_dq_sdr_0_x_sel[21]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_19 = %b", i_dq_sdr_0_x_sel[19]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_18 = %b", i_dq_sdr_0_x_sel[18]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_16 = %b", i_dq_sdr_0_x_sel[16]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_15 = %b", i_dq_sdr_0_x_sel[15]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_13 = %b", i_dq_sdr_0_x_sel[13]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_12 = %b", i_dq_sdr_0_x_sel[12]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_10 = %b", i_dq_sdr_0_x_sel[10]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_9 = %b", i_dq_sdr_0_x_sel[9]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_7 = %b", i_dq_sdr_0_x_sel[7]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_6 = %b", i_dq_sdr_0_x_sel[6]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_4 = %b", i_dq_sdr_0_x_sel[4]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_3 = %b", i_dq_sdr_0_x_sel[3]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_1 = %b", i_dq_sdr_0_x_sel[1]);
   $fdisplay(fd, "i_dq_sdr_0_x_sel_0 = %b", i_dq_sdr_0_x_sel[0]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_21 = %b", i_dq_sdr_0_fc_dly[21]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_20 = %b", i_dq_sdr_0_fc_dly[20]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_19 = %b", i_dq_sdr_0_fc_dly[19]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_18 = %b", i_dq_sdr_0_fc_dly[18]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_17 = %b", i_dq_sdr_0_fc_dly[17]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_16 = %b", i_dq_sdr_0_fc_dly[16]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_15 = %b", i_dq_sdr_0_fc_dly[15]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_14 = %b", i_dq_sdr_0_fc_dly[14]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_13 = %b", i_dq_sdr_0_fc_dly[13]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_12 = %b", i_dq_sdr_0_fc_dly[12]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_11 = %b", i_dq_sdr_0_fc_dly[11]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_10 = %b", i_dq_sdr_0_fc_dly[10]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_9 = %b", i_dq_sdr_0_fc_dly[9]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_8 = %b", i_dq_sdr_0_fc_dly[8]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_7 = %b", i_dq_sdr_0_fc_dly[7]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_6 = %b", i_dq_sdr_0_fc_dly[6]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_5 = %b", i_dq_sdr_0_fc_dly[5]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_4 = %b", i_dq_sdr_0_fc_dly[4]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_3 = %b", i_dq_sdr_0_fc_dly[3]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_2 = %b", i_dq_sdr_0_fc_dly[2]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_1 = %b", i_dq_sdr_0_fc_dly[1]);
   $fdisplay(fd, "i_dq_sdr_0_fc_dly_0 = %b", i_dq_sdr_0_fc_dly[0]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_10 = %b", i_dq_sdr_rt_pipe_en[10]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_9 = %b", i_dq_sdr_rt_pipe_en[9]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_8 = %b", i_dq_sdr_rt_pipe_en[8]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_7 = %b", i_dq_sdr_rt_pipe_en[7]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_6 = %b", i_dq_sdr_rt_pipe_en[6]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_5 = %b", i_dq_sdr_rt_pipe_en[5]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_4 = %b", i_dq_sdr_rt_pipe_en[4]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_3 = %b", i_dq_sdr_rt_pipe_en[3]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_2 = %b", i_dq_sdr_rt_pipe_en[2]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_1 = %b", i_dq_sdr_rt_pipe_en[1]);
   $fdisplay(fd, "i_dq_sdr_rt_pipe_en_0 = %b", i_dq_sdr_rt_pipe_en[0]);
   $fdisplay(fd, "i_dq_egress_mode_dig_76 = %b", i_dq_egress_mode_dig[76]);
   $fdisplay(fd, "i_dq_egress_mode_dig_71 = %b", i_dq_egress_mode_dig[71]);
   $fdisplay(fd, "i_dq_egress_mode_dig_70 = %b", i_dq_egress_mode_dig[70]);
   $fdisplay(fd, "i_dq_egress_mode_dig_69 = %b", i_dq_egress_mode_dig[69]);
   $fdisplay(fd, "i_dq_egress_mode_dig_64 = %b", i_dq_egress_mode_dig[64]);
   $fdisplay(fd, "i_dq_egress_mode_dig_63 = %b", i_dq_egress_mode_dig[63]);
   $fdisplay(fd, "i_dq_egress_mode_dig_62 = %b", i_dq_egress_mode_dig[62]);
   $fdisplay(fd, "i_dq_egress_mode_dig_57 = %b", i_dq_egress_mode_dig[57]);
   $fdisplay(fd, "i_dq_egress_mode_dig_56 = %b", i_dq_egress_mode_dig[56]);
   $fdisplay(fd, "i_dq_egress_mode_dig_55 = %b", i_dq_egress_mode_dig[55]);
   $fdisplay(fd, "i_dq_egress_mode_dig_50 = %b", i_dq_egress_mode_dig[50]);
   $fdisplay(fd, "i_dq_egress_mode_dig_49 = %b", i_dq_egress_mode_dig[49]);
   $fdisplay(fd, "i_dq_egress_mode_dig_48 = %b", i_dq_egress_mode_dig[48]);
   $fdisplay(fd, "i_dq_egress_mode_dig_43 = %b", i_dq_egress_mode_dig[43]);
   $fdisplay(fd, "i_dq_egress_mode_dig_42 = %b", i_dq_egress_mode_dig[42]);
   $fdisplay(fd, "i_dq_egress_mode_dig_41 = %b", i_dq_egress_mode_dig[41]);
   $fdisplay(fd, "i_dq_egress_mode_dig_36 = %b", i_dq_egress_mode_dig[36]);
   $fdisplay(fd, "i_dq_egress_mode_dig_35 = %b", i_dq_egress_mode_dig[35]);
   $fdisplay(fd, "i_dq_egress_mode_dig_34 = %b", i_dq_egress_mode_dig[34]);
   $fdisplay(fd, "i_dq_egress_mode_dig_29 = %b", i_dq_egress_mode_dig[29]);
   $fdisplay(fd, "i_dq_egress_mode_dig_28 = %b", i_dq_egress_mode_dig[28]);
   $fdisplay(fd, "i_dq_egress_mode_dig_27 = %b", i_dq_egress_mode_dig[27]);
   $fdisplay(fd, "i_dq_egress_mode_dig_22 = %b", i_dq_egress_mode_dig[22]);
   $fdisplay(fd, "i_dq_egress_mode_dig_21 = %b", i_dq_egress_mode_dig[21]);
   $fdisplay(fd, "i_dq_egress_mode_dig_20 = %b", i_dq_egress_mode_dig[20]);
   $fdisplay(fd, "i_dq_egress_mode_dig_15 = %b", i_dq_egress_mode_dig[15]);
   $fdisplay(fd, "i_dq_egress_mode_dig_14 = %b", i_dq_egress_mode_dig[14]);
   $fdisplay(fd, "i_dq_egress_mode_dig_13 = %b", i_dq_egress_mode_dig[13]);
   $fdisplay(fd, "i_dq_egress_mode_dig_8 = %b", i_dq_egress_mode_dig[8]);
   $fdisplay(fd, "i_dq_egress_mode_dig_7 = %b", i_dq_egress_mode_dig[7]);
   $fdisplay(fd, "i_dq_egress_mode_dig_6 = %b", i_dq_egress_mode_dig[6]);
   $fdisplay(fd, "i_dq_egress_mode_dig_1 = %b", i_dq_egress_mode_dig[1]);
   $fdisplay(fd, "i_dq_egress_mode_dig_0 = %b", i_dq_egress_mode_dig[0]);
   $fdisplay(fd, "i_dq_egress_mode_ana_62 = %b", i_dq_egress_mode_ana[62]);
   $fdisplay(fd, "i_dq_egress_mode_ana_61 = %b", i_dq_egress_mode_ana[61]);
   $fdisplay(fd, "i_dq_egress_mode_ana_60 = %b", i_dq_egress_mode_ana[60]);
   $fdisplay(fd, "i_dq_egress_mode_ana_56 = %b", i_dq_egress_mode_ana[56]);
   $fdisplay(fd, "i_dq_egress_mode_ana_55 = %b", i_dq_egress_mode_ana[55]);
   $fdisplay(fd, "i_dq_egress_mode_ana_54 = %b", i_dq_egress_mode_ana[54]);
   $fdisplay(fd, "i_dq_egress_mode_ana_50 = %b", i_dq_egress_mode_ana[50]);
   $fdisplay(fd, "i_dq_egress_mode_ana_49 = %b", i_dq_egress_mode_ana[49]);
   $fdisplay(fd, "i_dq_egress_mode_ana_48 = %b", i_dq_egress_mode_ana[48]);
   $fdisplay(fd, "i_dq_egress_mode_ana_44 = %b", i_dq_egress_mode_ana[44]);
   $fdisplay(fd, "i_dq_egress_mode_ana_43 = %b", i_dq_egress_mode_ana[43]);
   $fdisplay(fd, "i_dq_egress_mode_ana_42 = %b", i_dq_egress_mode_ana[42]);
   $fdisplay(fd, "i_dq_egress_mode_ana_38 = %b", i_dq_egress_mode_ana[38]);
   $fdisplay(fd, "i_dq_egress_mode_ana_37 = %b", i_dq_egress_mode_ana[37]);
   $fdisplay(fd, "i_dq_egress_mode_ana_36 = %b", i_dq_egress_mode_ana[36]);
   $fdisplay(fd, "i_dq_egress_mode_ana_32 = %b", i_dq_egress_mode_ana[32]);
   $fdisplay(fd, "i_dq_egress_mode_ana_31 = %b", i_dq_egress_mode_ana[31]);
   $fdisplay(fd, "i_dq_egress_mode_ana_30 = %b", i_dq_egress_mode_ana[30]);
   $fdisplay(fd, "i_dq_egress_mode_ana_26 = %b", i_dq_egress_mode_ana[26]);
   $fdisplay(fd, "i_dq_egress_mode_ana_25 = %b", i_dq_egress_mode_ana[25]);
   $fdisplay(fd, "i_dq_egress_mode_ana_24 = %b", i_dq_egress_mode_ana[24]);
   $fdisplay(fd, "i_dq_egress_mode_ana_20 = %b", i_dq_egress_mode_ana[20]);
   $fdisplay(fd, "i_dq_egress_mode_ana_19 = %b", i_dq_egress_mode_ana[19]);
   $fdisplay(fd, "i_dq_egress_mode_ana_18 = %b", i_dq_egress_mode_ana[18]);
   $fdisplay(fd, "i_dq_egress_mode_ana_14 = %b", i_dq_egress_mode_ana[14]);
   $fdisplay(fd, "i_dq_egress_mode_ana_13 = %b", i_dq_egress_mode_ana[13]);
   $fdisplay(fd, "i_dq_egress_mode_ana_12 = %b", i_dq_egress_mode_ana[12]);
   $fdisplay(fd, "i_dq_egress_mode_ana_8 = %b", i_dq_egress_mode_ana[8]);
   $fdisplay(fd, "i_dq_egress_mode_ana_7 = %b", i_dq_egress_mode_ana[7]);
   $fdisplay(fd, "i_dq_egress_mode_ana_6 = %b", i_dq_egress_mode_ana[6]);
   $fdisplay(fd, "i_dq_egress_mode_ana_2 = %b", i_dq_egress_mode_ana[2]);
   $fdisplay(fd, "i_dq_egress_mode_ana_1 = %b", i_dq_egress_mode_ana[1]);
   $fdisplay(fd, "i_dq_egress_mode_ana_0 = %b", i_dq_egress_mode_ana[0]);
   $fdisplay(fd, "i_pll_clk_270 = %b", i_pll_clk_270);
   $fdisplay(fd, "i_pll_clk_180 = %b", i_pll_clk_180);
   $fdisplay(fd, "i_pll_clk_90 = %b", i_pll_clk_90);
   $fdisplay(fd, "i_pll_clk_0 = %b", i_pll_clk_0);
   $fdisplay(fd, "i_rst = %b", i_rst);
   $fdisplay(fd, "i_scan_mode = %b", i_scan_mode);
   $fdisplay(fd, "i_scan_clk = %b", i_scan_clk);
endtask

task oprint_ddr_ca (input integer fd);

   $fdisplay(fd, "INFO: Edge Trigger [%t] ...", $realtime);
   $fdisplay(fd, "o_dqs_pad_bscan_c_0 = %b", o_dqs_pad_bscan_c[0]);
   $fdisplay(fd, "o_dqs_pad_bscan_t_0 = %b", o_dqs_pad_bscan_t[0]);
   $fdisplay(fd, "o_dq_pad_bscan_t_10 = %b", o_dq_pad_bscan_t[10]);
   $fdisplay(fd, "o_dq_pad_bscan_t_9 = %b", o_dq_pad_bscan_t[9]);
   $fdisplay(fd, "o_dq_pad_bscan_t_8 = %b", o_dq_pad_bscan_t[8]);
   $fdisplay(fd, "o_dq_pad_bscan_t_7 = %b", o_dq_pad_bscan_t[7]);
   $fdisplay(fd, "o_dq_pad_bscan_t_6 = %b", o_dq_pad_bscan_t[6]);
   $fdisplay(fd, "o_dq_pad_bscan_t_5 = %b", o_dq_pad_bscan_t[5]);
   $fdisplay(fd, "o_dq_pad_bscan_t_4 = %b", o_dq_pad_bscan_t[4]);
   $fdisplay(fd, "o_dq_pad_bscan_t_3 = %b", o_dq_pad_bscan_t[3]);
   $fdisplay(fd, "o_dq_pad_bscan_t_2 = %b", o_dq_pad_bscan_t[2]);
   $fdisplay(fd, "o_dq_pad_bscan_t_1 = %b", o_dq_pad_bscan_t[1]);
   $fdisplay(fd, "o_dq_pad_bscan_t_0 = %b", o_dq_pad_bscan_t[0]);
   $fdisplay(fd, "o_dq_core_eg_10 = %b", o_dq_core_eg[10]);
   $fdisplay(fd, "o_dq_core_eg_9 = %b", o_dq_core_eg[9]);
   $fdisplay(fd, "o_dq_core_eg_8 = %b", o_dq_core_eg[8]);
   $fdisplay(fd, "o_dq_core_eg_7 = %b", o_dq_core_eg[7]);
   $fdisplay(fd, "o_dq_core_eg_6 = %b", o_dq_core_eg[6]);
   $fdisplay(fd, "o_dq_core_eg_5 = %b", o_dq_core_eg[5]);
   $fdisplay(fd, "o_dq_core_eg_4 = %b", o_dq_core_eg[4]);
   $fdisplay(fd, "o_dq_core_eg_3 = %b", o_dq_core_eg[3]);
   $fdisplay(fd, "o_dq_core_eg_2 = %b", o_dq_core_eg[2]);
   $fdisplay(fd, "o_dq_core_eg_1 = %b", o_dq_core_eg[1]);
   $fdisplay(fd, "o_dq_core_eg_0 = %b", o_dq_core_eg[0]);
   $fdisplay(fd, "o_dq_core_ig_10 = %b", o_dq_core_ig[10]);
   $fdisplay(fd, "o_dq_core_ig_9 = %b", o_dq_core_ig[9]);
   $fdisplay(fd, "o_dq_core_ig_8 = %b", o_dq_core_ig[8]);
   $fdisplay(fd, "o_dq_core_ig_7 = %b", o_dq_core_ig[7]);
   $fdisplay(fd, "o_dq_core_ig_6 = %b", o_dq_core_ig[6]);
   $fdisplay(fd, "o_dq_core_ig_5 = %b", o_dq_core_ig[5]);
   $fdisplay(fd, "o_dq_core_ig_4 = %b", o_dq_core_ig[4]);
   $fdisplay(fd, "o_dq_core_ig_3 = %b", o_dq_core_ig[3]);
   $fdisplay(fd, "o_dq_core_ig_2 = %b", o_dq_core_ig[2]);
   $fdisplay(fd, "o_dq_core_ig_1 = %b", o_dq_core_ig[1]);
   $fdisplay(fd, "o_dq_core_ig_0 = %b", o_dq_core_ig[0]);
   $fdisplay(fd, "o_dqs_core_eg_8 = %b", o_dqs_core_eg[8]);
   $fdisplay(fd, "o_dqs_core_eg_7 = %b", o_dqs_core_eg[7]);
   $fdisplay(fd, "o_dqs_core_eg_6 = %b", o_dqs_core_eg[6]);
   $fdisplay(fd, "o_dqs_core_eg_5 = %b", o_dqs_core_eg[5]);
   $fdisplay(fd, "o_dqs_core_eg_4 = %b", o_dqs_core_eg[4]);
   $fdisplay(fd, "o_dqs_core_eg_3 = %b", o_dqs_core_eg[3]);
   $fdisplay(fd, "o_dqs_core_eg_2 = %b", o_dqs_core_eg[2]);
   $fdisplay(fd, "o_dqs_core_eg_1 = %b", o_dqs_core_eg[1]);
   $fdisplay(fd, "o_dqs_core_eg_0 = %b", o_dqs_core_eg[0]);
   $fdisplay(fd, "o_dqs_core_ig_0 = %b", o_dqs_core_ig[0]);
   $fdisplay(fd, "o_dqs_ren_pi_phase_sta = %b", o_dqs_ren_pi_phase_sta);
   $fdisplay(fd, "o_dqs_rcs_pi_phase_sta = %b", o_dqs_rcs_pi_phase_sta);
   $fdisplay(fd, "o_dq_sdr_43 = %b", o_dq_sdr[43]);
   $fdisplay(fd, "o_dq_sdr_42 = %b", o_dq_sdr[42]);
   $fdisplay(fd, "o_dq_sdr_41 = %b", o_dq_sdr[41]);
   $fdisplay(fd, "o_dq_sdr_40 = %b", o_dq_sdr[40]);
   $fdisplay(fd, "o_dq_sdr_39 = %b", o_dq_sdr[39]);
   $fdisplay(fd, "o_dq_sdr_38 = %b", o_dq_sdr[38]);
   $fdisplay(fd, "o_dq_sdr_37 = %b", o_dq_sdr[37]);
   $fdisplay(fd, "o_dq_sdr_36 = %b", o_dq_sdr[36]);
   $fdisplay(fd, "o_dq_sdr_35 = %b", o_dq_sdr[35]);
   $fdisplay(fd, "o_dq_sdr_34 = %b", o_dq_sdr[34]);
   $fdisplay(fd, "o_dq_sdr_33 = %b", o_dq_sdr[33]);
   $fdisplay(fd, "o_dq_sdr_32 = %b", o_dq_sdr[32]);
   $fdisplay(fd, "o_dq_sdr_31 = %b", o_dq_sdr[31]);
   $fdisplay(fd, "o_dq_sdr_30 = %b", o_dq_sdr[30]);
   $fdisplay(fd, "o_dq_sdr_29 = %b", o_dq_sdr[29]);
   $fdisplay(fd, "o_dq_sdr_28 = %b", o_dq_sdr[28]);
   $fdisplay(fd, "o_dq_sdr_27 = %b", o_dq_sdr[27]);
   $fdisplay(fd, "o_dq_sdr_26 = %b", o_dq_sdr[26]);
   $fdisplay(fd, "o_dq_sdr_25 = %b", o_dq_sdr[25]);
   $fdisplay(fd, "o_dq_sdr_24 = %b", o_dq_sdr[24]);
   $fdisplay(fd, "o_dq_sdr_23 = %b", o_dq_sdr[23]);
   $fdisplay(fd, "o_dq_sdr_22 = %b", o_dq_sdr[22]);
   $fdisplay(fd, "o_dq_sdr_21 = %b", o_dq_sdr[21]);
   $fdisplay(fd, "o_dq_sdr_20 = %b", o_dq_sdr[20]);
   $fdisplay(fd, "o_dq_sdr_19 = %b", o_dq_sdr[19]);
   $fdisplay(fd, "o_dq_sdr_18 = %b", o_dq_sdr[18]);
   $fdisplay(fd, "o_dq_sdr_17 = %b", o_dq_sdr[17]);
   $fdisplay(fd, "o_dq_sdr_16 = %b", o_dq_sdr[16]);
   $fdisplay(fd, "o_dq_sdr_15 = %b", o_dq_sdr[15]);
   $fdisplay(fd, "o_dq_sdr_14 = %b", o_dq_sdr[14]);
   $fdisplay(fd, "o_dq_sdr_13 = %b", o_dq_sdr[13]);
   $fdisplay(fd, "o_dq_sdr_12 = %b", o_dq_sdr[12]);
   $fdisplay(fd, "o_dq_sdr_11 = %b", o_dq_sdr[11]);
   $fdisplay(fd, "o_dq_sdr_10 = %b", o_dq_sdr[10]);
   $fdisplay(fd, "o_dq_sdr_9 = %b", o_dq_sdr[9]);
   $fdisplay(fd, "o_dq_sdr_8 = %b", o_dq_sdr[8]);
   $fdisplay(fd, "o_dq_sdr_7 = %b", o_dq_sdr[7]);
   $fdisplay(fd, "o_dq_sdr_6 = %b", o_dq_sdr[6]);
   $fdisplay(fd, "o_dq_sdr_5 = %b", o_dq_sdr[5]);
   $fdisplay(fd, "o_dq_sdr_4 = %b", o_dq_sdr[4]);
   $fdisplay(fd, "o_dq_sdr_3 = %b", o_dq_sdr[3]);
   $fdisplay(fd, "o_dq_sdr_2 = %b", o_dq_sdr[2]);
   $fdisplay(fd, "o_dq_sdr_1 = %b", o_dq_sdr[1]);
   $fdisplay(fd, "o_dq_sdr_0 = %b", o_dq_sdr[0]);
   $fdisplay(fd, "o_dq_sa_43 = %b", o_dq_sa[43]);
   $fdisplay(fd, "o_dq_sa_42 = %b", o_dq_sa[42]);
   $fdisplay(fd, "o_dq_sa_41 = %b", o_dq_sa[41]);
   $fdisplay(fd, "o_dq_sa_40 = %b", o_dq_sa[40]);
   $fdisplay(fd, "o_dq_sa_39 = %b", o_dq_sa[39]);
   $fdisplay(fd, "o_dq_sa_38 = %b", o_dq_sa[38]);
   $fdisplay(fd, "o_dq_sa_37 = %b", o_dq_sa[37]);
   $fdisplay(fd, "o_dq_sa_36 = %b", o_dq_sa[36]);
   $fdisplay(fd, "o_dq_sa_35 = %b", o_dq_sa[35]);
   $fdisplay(fd, "o_dq_sa_34 = %b", o_dq_sa[34]);
   $fdisplay(fd, "o_dq_sa_33 = %b", o_dq_sa[33]);
   $fdisplay(fd, "o_dq_sa_32 = %b", o_dq_sa[32]);
   $fdisplay(fd, "o_dq_sa_31 = %b", o_dq_sa[31]);
   $fdisplay(fd, "o_dq_sa_30 = %b", o_dq_sa[30]);
   $fdisplay(fd, "o_dq_sa_29 = %b", o_dq_sa[29]);
   $fdisplay(fd, "o_dq_sa_28 = %b", o_dq_sa[28]);
   $fdisplay(fd, "o_dq_sa_27 = %b", o_dq_sa[27]);
   $fdisplay(fd, "o_dq_sa_26 = %b", o_dq_sa[26]);
   $fdisplay(fd, "o_dq_sa_25 = %b", o_dq_sa[25]);
   $fdisplay(fd, "o_dq_sa_24 = %b", o_dq_sa[24]);
   $fdisplay(fd, "o_dq_sa_23 = %b", o_dq_sa[23]);
   $fdisplay(fd, "o_dq_sa_22 = %b", o_dq_sa[22]);
   $fdisplay(fd, "o_dq_sa_21 = %b", o_dq_sa[21]);
   $fdisplay(fd, "o_dq_sa_20 = %b", o_dq_sa[20]);
   $fdisplay(fd, "o_dq_sa_19 = %b", o_dq_sa[19]);
   $fdisplay(fd, "o_dq_sa_18 = %b", o_dq_sa[18]);
   $fdisplay(fd, "o_dq_sa_17 = %b", o_dq_sa[17]);
   $fdisplay(fd, "o_dq_sa_16 = %b", o_dq_sa[16]);
   $fdisplay(fd, "o_dq_sa_15 = %b", o_dq_sa[15]);
   $fdisplay(fd, "o_dq_sa_14 = %b", o_dq_sa[14]);
   $fdisplay(fd, "o_dq_sa_13 = %b", o_dq_sa[13]);
   $fdisplay(fd, "o_dq_sa_12 = %b", o_dq_sa[12]);
   $fdisplay(fd, "o_dq_sa_11 = %b", o_dq_sa[11]);
   $fdisplay(fd, "o_dq_sa_10 = %b", o_dq_sa[10]);
   $fdisplay(fd, "o_dq_sa_9 = %b", o_dq_sa[9]);
   $fdisplay(fd, "o_dq_sa_8 = %b", o_dq_sa[8]);
   $fdisplay(fd, "o_dq_sa_7 = %b", o_dq_sa[7]);
   $fdisplay(fd, "o_dq_sa_6 = %b", o_dq_sa[6]);
   $fdisplay(fd, "o_dq_sa_5 = %b", o_dq_sa[5]);
   $fdisplay(fd, "o_dq_sa_4 = %b", o_dq_sa[4]);
   $fdisplay(fd, "o_dq_sa_3 = %b", o_dq_sa[3]);
   $fdisplay(fd, "o_dq_sa_2 = %b", o_dq_sa[2]);
   $fdisplay(fd, "o_dq_sa_1 = %b", o_dq_sa[1]);
   $fdisplay(fd, "o_dq_sa_0 = %b", o_dq_sa[0]);
   $fdisplay(fd, "o_rcs = %b", o_rcs);
   $fdisplay(fd, "o_dfird_clk_2 = %b", o_dfird_clk_2);
   $fdisplay(fd, "o_dfird_clk_1 = %b", o_dfird_clk_1);
   $fdisplay(fd, "o_dfiwr_clk_2 = %b", o_dfiwr_clk_2);
   $fdisplay(fd, "o_dfiwr_clk_1 = %b", o_dfiwr_clk_1);
   $fdisplay(fd, "o_rx_sdr_clk = %b", o_rx_sdr_clk);
   $fdisplay(fd, "o_phy_clk = %b", o_phy_clk);
   $fdisplay(fd, "o_tst_clk_1 = %b", o_tst_clk[1]);
   $fdisplay(fd, "o_tst_clk_0 = %b", o_tst_clk[0]);
endtask
