/*
:name: string_icompare
:description: string.icompare()  tests
:tags: 6.16.7
*/
module top();
	string a = "Test";
	string b = "TEST";
	int c = a.icompare(b);
endmodule
