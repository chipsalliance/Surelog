/*
:name: 22.12--line-illegal-3
:description: The number parameter shall be a positive integer that specifies the new line number
:should_fail: 1
:tags: 22.12
:type: preprocessing
*/
`line -12 "somefile" 3
