module top(b);
input b;

task DoSomething(input [7:0] A);
endtask
endmodule
