localparam              AWIDTH                       = 16 ;

localparam [AWIDTH:0] MAP      ={
  AWIDTH                                     
                                              };

module top();

  parameter D =MAP;

endmodule