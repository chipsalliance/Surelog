/*********************************************************************************
Copyright (c) 2021 Wavious LLC

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.

*********************************************************************************/

`ifdef SYNTHESIS
`else 
// AMS netlist generated by the AMS Unified netlister
// IC subversion:  ICADVM20.1-64b.14 
// Xcelium version: 20.09-s003
// Copyright(C) 2005-2009, Cadence Design Systems, Inc
// User: shadzibabic Pid: 26886
// Design library name: wphy_gf12lp_ips_sim_lib
// Design cell name: wphy_clkmux_3to1_diff_tb
// Design view name: config_vlog
// Solver: Spectre



// Library - wphy_gf12lp_ips_lib, Cell - wphy_clkmux_3to1_diff, View -
//schematic
// LAST TIME SAVED: Jan 21 14:06:49 2021
// NETLIST TIME: Jan 29 16:30:00 2021
`timescale 1ps / 1ps 




 

`endif //SYNTHESIS 
module wphy_clkmux_3to1_diff (out_c, out_t,   in01_c, in01_t, 
    in10_c, in10_t, in11_c, in11_t, s
`ifdef WLOGIC_NO_PG 
`else  
 ,vdda  
 ,vss 
`endif //WLOGIC_NO_PG 
);

`ifdef WLOGIC_NO_PG
wire vdda;
assign vdda=1'b1;
wire vss;
assign vss=1'b0;
`else
inout vdda;
inout vss;
`endif


output  out_c, out_t;



input  in01_c, in01_t, in10_c, in10_t, in11_c, in11_t;

input [1:0]  s;

// Buses in the design 
`ifdef SYNTHESIS 
`else

wire  [1:0]  sb;

wire  [1:0]  s_buf;


wphy_clkmux_3to1_diff_NAND2_D1_GL16_RVT NAND3 ( .y(s00b), .b(sb[0]), .a(sb[1]), .tielo(vss), 
    .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_NAND2_D1_GL16_RVT NAND2 ( .y(s10b), .b(sb[0]), .a(s_buf[1]), 
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_NAND2_D1_GL16_RVT NAND1 ( .y(s11b), .b(s_buf[0]), .a(s_buf[1]), 
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_NAND2_D1_GL16_RVT NAND0 ( .y(s01b), .b(s_buf[0]), .a(sb[1]), 
    .tielo(vss), .vdd(vdda), .vss(vss), .tiehi(vdda));

wphy_clkmux_3to1_diff_PU_D2_GL16_RVT PU0 ( .vdd(vdda), .en(s00b), .y(yb_t));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT03_1 ( .out(mux_slw_cb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT03_0 ( .out(mux_slw_cb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT4_3 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT4_2 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT4_1 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT4_0 ( .out(yb_t), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_cb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT3_1 ( .out(mux_slw_tb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT3_0 ( .out(mux_slw_tb), .en(s11), .enb(s11b), 
    .vss(vss), .in(in11_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT1_3 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT1_2 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT1_1 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT1_0 ( .out(yb_c), .en(s01), .enb(s01b), .vss(vss), 
    .in(in01_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT02_1 ( .out(mux_slw_cb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT02_0 ( .out(mux_slw_cb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT5_3 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT5_2 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT5_1 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT5_0 ( .out(yb_c), .en(s_buf[1]), .enb(sb[1]), 
    .vss(vss), .in(mux_slw_tb), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT2_1 ( .out(mux_slw_tb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT2_0 ( .out(mux_slw_tb), .en(s10), .enb(s10b), 
    .vss(vss), .in(in10_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT01_3 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT01_2 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT01_1 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT INVT01_0 ( .out(yb_t), .en(s01), .enb(s01b), 
    .vss(vss), .in(in01_t), .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV7 ( .in(s00b), .vss(vss), .out(s00), .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV5_1 ( .in(s[1]), .vss(vss), .out(sb[1]), 
    .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV5_0 ( .in(s[0]), .vss(vss), .out(sb[0]), 
    .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV6_1 ( .in(sb[1]), .vss(vss), .out(s_buf[1]), 
    .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV6_0 ( .in(sb[0]), .vss(vss), .out(s_buf[0]), 
    .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV4 ( .in(s01b), .vss(vss), .out(s01), .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV3 ( .in(s10b), .vss(vss), .out(s10), .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D2_GL16_RVT INV2 ( .in(s11b), .vss(vss), .out(s11), .vdd(vdda));

wphy_clkmux_3to1_diff_PUDUM_D2_GL16_RVT PUDUM ( .vdd(vdda), .tiehi(vdda));

wphy_clkmux_3to1_diff_INV_D16_GL16_RVT INV9 ( .in(yb_c), .vss(vss), .out(out_c), .vdd(vdda));

wphy_clkmux_3to1_diff_INV_D16_GL16_RVT INV8 ( .in(yb_t), .vss(vss), .out(out_t), .vdd(vdda));

wphy_clkmux_3to1_diff_PD_D2_GL16_RVT PD0 ( .vss(vss), .enb(s00), .y(yb_c));

wphy_clkmux_3to1_diff_PDDUM_D2_GL16_RVT PDDUM ( .vss(vss), .tielo(vss));

`ifdef WPHY_ANA_TIMING

specify

  if (s==='b01) (in01_t => out_t) = 32;
  if (s==='b10) (in10_t => out_t) = 47;
  if (s==='b11) (in11_t => out_t) = 47;

endspecify

`endif

`endif //SYNTHESIS 
endmodule
`ifdef SYNTHESIS
`else
// Library - wphy_gf12lp_ips_sim_lib, Cell - wphy_clkmux_3to1_diff_tb,
//View - schematic
// LAST TIME SAVED: Jan 29 16:17:51 2021
// NETLIST TIME: Jan 29 16:30:00 2021
`timescale 1ps / 1ps 




 




 // END AMS-UNL Netlist

//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_PDDUM_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_PDDUM_D2_GL16_RVT (  tielo
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input tielo;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_PD_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_PD_D2_GL16_RVT ( enb, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss
`endif //WLOGIC_MODEL_NO_PG
); 

  input y;
  input enb;

`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss ;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign y =  enb ? 1'b0 : 1'bz;

endmodule
//systemVerilog HDL for "wavshared_ln08lpu_dig_lib", "wphy_clkmux_3to1_diff_INV_D16_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_INV_D16_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_PUDUM_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_PUDUM_D2_GL16_RVT ( tiehi
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input tiehi;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_INV_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_INV_D2_GL16_RVT ( in, out
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

   assign out = ~in;

endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_INVT_D2_GL16_RVT( in, out, en, enb
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd, vss
`endif //WLOGIC_MODEL_NO_PG
);

  input in;
  input en, enb;
  output out;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

  wire out;

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign out = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

  assign out= (en) ? ~in:1'bz;


endmodule
//systemVerilog HDL for "wavshared_tsmc12ffc_lib", "wphy_clkmux_3to1_diff_PU_D2_GL16_RVT" "systemVerilog"


module wphy_clkmux_3to1_diff_PU_D2_GL16_RVT ( en, y
`ifdef WLOGIC_MODEL_NO_PG
`else
, vdd 
`endif //WLOGIC_MODEL_NO_PG
);

  input y;
  input en;
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG

 assign y = en ? 1'bz : 1'b1;

endmodule



module wphy_clkmux_3to1_diff_NAND2_D1_GL16_RVT ( y, a, b
`ifdef WLOGIC_MODEL_NO_TIE
`else
,tielo, tiehi
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
, vss, vdd 
`endif //WLOGIC_MODEL_NO_PG
); 

  input b;
  input a;
  output y;
`ifdef WLOGIC_MODEL_NO_TIE
`else
  input tiehi;
  input tielo;
`endif //WLOGIC_MODEL_NO_TIE
`ifdef WLOGIC_MODEL_NO_PG
`else
  inout vdd;
  inout vss;
`endif //WLOGIC_MODEL_NO_PG

`ifdef WLOGIC_MODEL_NO_TIE
`else

`ifdef WLOGIC_MODEL_TIE_CHECK
  wire   signals_ok;
  assign signals_ok = tiehi & ~tielo;
  
  assign y = (signals_ok) ? 1'bz : 1'bx;
`endif // WLOGIC_MODEL_TIE_CHECK

`endif //WLOGIC_MODEL_NO_TIE

`ifdef WLOGIC_MODEL_NO_PG
`else

`ifdef WLOGIC_MODEL_PWR_CHECK
  wire   power_ok;
  assign power_ok = ~vss & vdd;
  
  assign y = (power_ok) ? 1'bz : 1'bx;

`endif //WLOGIC_MODEL_PWR_CHECK

`endif //WLOGIC_MODEL_NO_PG


 assign y = ~(a&b);

endmodule
`endif //SYNTHESIS
