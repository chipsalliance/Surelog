// Copyright (C) 2019-2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC


/*
:name: basic-unpacked
:description: Test unpacked arrays support
:tags: 7.4.2 7.4
*/
module top ();

bit _bit [7:0];
logic _logic [7:0];
reg _reg [7:0];

endmodule
