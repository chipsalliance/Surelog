module dut();

assign mido_bytes_in[1][2][3] = 1'b0;
assign state_d[2][3][4][5:6] = 8'b10101010;
assign state_d1[10:11] = 8'b10101010;
endmodule
