/*
:name: class_member_test_28
:description: Test
:should_fail: 0
:tags: 8.3
*/
class myclass;
function void shifter;
  for ( ; shft_idx < n_bits;
       shft_idx++) begin
  end
endfunction
endclass