/*
:name: typedef_test_2
:description: Test
:should_fail: 0
:tags: 6.18
*/
typedef reg quartet[3:0];