module top;
initial
   if (0) $error("ASDF");
endmodule
