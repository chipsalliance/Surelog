module top(output logic o);
   function automatic logic theta();
      for (int x = 0 ; x < 5 ; x++) begin
	      int a;
      end
   endfunction : theta
endmodule : top
